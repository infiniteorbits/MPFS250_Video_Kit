--=================================================================================================
-- File Name                           : RGBtoYCbCr.vhd
-- Description                                             : Supporting both Native mode and AXI4 Stream mode

-- Targeted device                     : Microsemi-SoC
-- Author                              : India Solutions Team
--
-- COPYRIGHT 2021 BY MICROSEMI
-- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS FROM MICROSEMI
-- CORP. IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM MICROSEMI FOR USE OF THIS
-- FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND NO BACK-UP OF THE FILE SHOULD BE MADE.
--
--=================================================================================================
--=================================================================================================
-- Libraries
--=================================================================================================
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
--=================================================================================================
-- RGBtoYCbCr entity declaration
--=================================================================================================                                                          
entity RGBtoYCbCr is
  generic(
-- Generic List
    -- Specifies the data width
    G_RGB_DATA_BIT_WIDTH : integer := 8;

    G_YCbCr_DATA_BIT_WIDTH : integer := 8;

    G_YCbCr_FORMAT : integer := 2;      --  3= YCbCr444 and 2 = YCbCr422

    G_FORMAT : integer := 0;            --  0= Native and 1 = AXI4 Streaming

    TGIGEN_DISPLAY_SYMBOL : integer := 1
    );
  port (
-- Port List
    -- System reset     
    RESET_N_I : in std_logic;

    -- System clock
    CLOCK_I : in std_logic;

    -- Specifies the input data is valid or not
    DATA_VALID_I : in std_logic;

    -- Data input to SLAVE
    TDATA_I : in std_logic_vector(3*G_RGB_DATA_BIT_WIDTH-1 downto 0);

    -- Specifies the valid control signal to SLAVE
    TVALID_I : in std_logic;

    TUSER_I : in std_logic_vector(3 downto 0);

    TREADY_O : out std_logic;

    -- Red data input     
    RED_I : in std_logic_vector ((G_RGB_DATA_BIT_WIDTH - 1) downto 0);

    -- Green data input 
    GREEN_I : in std_logic_vector ((G_RGB_DATA_BIT_WIDTH - 1) downto 0);

    -- Blue input  
    BLUE_I : in std_logic_vector ((G_RGB_DATA_BIT_WIDTH - 1) downto 0);

    -- Specifies the valid output data
    DATA_VALID_O : out std_logic;

    -- Converted data output Luminance                                                                                                             
    Y_OUT_O : out std_logic_vector ((G_YCbCr_DATA_BIT_WIDTH - 1) downto 0);

    -- Converted data output 3Chroma  
    Cb_OUT_O : out std_logic_vector ((G_YCbCr_DATA_BIT_WIDTH - 1) downto 0);

    -- Converted data output Chroma  
    Cr_OUT_O : out std_logic_vector ((G_YCbCr_DATA_BIT_WIDTH - 1) downto 0);

    -- YCbCr422 Y Component
    Y_OUT : out std_logic_vector ((G_YCbCr_DATA_BIT_WIDTH - 1) downto 0);

    -- YCbCr422 C Component
    C_OUT : out std_logic_vector ((G_YCbCr_DATA_BIT_WIDTH - 1) downto 0);

    -- Data output from MASTER
    TDATA_O : out std_logic_vector(G_YCbCr_FORMAT*G_YCbCr_DATA_BIT_WIDTH-1 downto 0);

    TUSER_O : out std_logic_vector(3 downto 0);

    TSTRB_O : out std_logic_vector(G_YCbCr_DATA_BIT_WIDTH/8 -1 downto 0);

    TKEEP_O : out std_logic_vector(G_YCbCr_DATA_BIT_WIDTH/8 -1 downto 0);

    TLAST_O  : out std_logic;
    -- Specifies the valid control signal from MASTER
    TVALID_O : out std_logic

    );
end RGBtoYCbCr;

`protect begin_protected
`protect version=1
`protect author="author-a", author_info="author-a-details"
`protect encrypt_agent="encryptP1735.pl", encrypt_agent_info="Synplify encryption scripts"

`protect key_keyowner="Synplicity", key_keyname="SYNP05_001", key_method="rsa"
`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_block
uSv1JqkTm1EmiMxs4INN4atlU58ollS5Pm5GzNPjYV6y6gWTshK7I4EyS//CjQ6XNGqk1ktr11N0
aURO6TQQkhXtGaviEgDSwkLkSYOTpwj5khYibQKSIYjCmwcWj8dztko978qxtNUPXVx3JxbbPj8b
cVhrLLSLCX2pzlgr6qH3Fl7XqTR0Q5P/VEN5RWGWYu1HqysbhY1UsyjIP91rJYyZG0srIr+5xNGg
mwe+3++ycJZR1aJ2FvOYHnWCs6S5YKgnUDMr7NNve/m/1qTNjBsjRevv16v0od517f+E74LkGwwS
RUJwyEIvOU6ZIXxM9HZhstL50oKi7hlD4W6r4Q==

`protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`protect encoding=(enctype="base64", line_length=76, bytes=128)
`protect key_block
W2awRCTmUqGIUJBpONO1zvaGqX6f9UpZFSte+BTy9uKGgv0FpvXw3KGzYg+FtQQRhUUty9N0bTVW
3RGCwnVVcTl99L8llU++PDadqrD9jDaKV9Mvjh5mEj9owKbmLwW135SJdROyFu9xgsVLKj+ZagOu
hBwMw1G0aYJkiZR7d1k=

`protect key_keyowner="Microsemi Corporation", key_keyname="MSC-IP-KEY-RSA", key_method="rsa"
`protect encoding=(enctype="base64", line_length=76, bytes=960)
`protect key_block
qU4SVu2u538DeBOvGDQlRA66ytPRSdraDztPe5UxDlnnQDPpv99XXBVAwUQNg1CeqqIkT0aLcoLT
wmfQw0YmsgTdEezJwZT26yFVg21VzqeqPX2XXS5xAHKAAXAhwaH2+JLc20ZBwtC8IAxTWBG4svbT
ffzfkavG7F9UJK4dqifdoakTFkxsVPqnQ05K+cYrD2G2fKVoXSKf7tTLiKiX7ao8l57t9RSuMqHJ
V04OI5dmkurS+3k7T51LuZ/7gI3e4xp4PJ3MwJ709/H2s+MEyFveLHiMzZll+Q2B5GEiCMDr6iZX
0hUNI+jxDMaDcGHmKOYQEvVqCvVIfW2Kh/tl9MtT7oEVwLpHf0Jn1HwSUSUa6GDcVSw43MYYQqq8
UvZ9Yu4yFz4+47CEWVWT1pT3DRHX2HuEndqKV+onFRSHdY3XZfPB56dr+6n+DtnUgBxGIgh2qO6/
AVKk9hW7NDiyvVt8hZiSgtoYflzIVlHraBV411iByNqwThmBiJQPo+a3u9RwQrNrzDmwObiaHoYW
1JMi3j1vtJ66H1aQ5oHdU4BgDvkA9yuYkhehof+09rfpwfCGLUOhGtYWVfFYJFxH7nC6+5dOG058
mzONlCTfbf+intmnVj8swij8E0RSxBu3THmrMXqBcSnCBgZ9nFtBVW9XHqCIYPW+IzuSjO9h7Iq4
+VRjwFPNI4gmoqxtPKFdLdLWBsPz+46/D2h97JsjsNiTyWPcd43XH9D1EMU04OAlr2LvxAEo4FIS
7wXTZg9XOEeWB++uWO3dHrofugb4am5jtuLtG4CTUghl/dQu1lSIHYWi4jmqnJVUBAV6fn2hAPSe
EWzF0myOdisVX8anVMJQkY5A/5MbEaW+PpWOgH0vBE9hZN/67PjI+iVWjhVAzL0rvzt2by+nrzfO
m/c3n3B7FlLSR1CVIdiIj+iI6WvT4kVivusUxMmVDELBAYOWqcNVpxZiYIf7LhICPR7QTHQthYlv
6axGgoQk/H8Us+09ll7HWh3Ka+cJfKcFJ6urHrBgGfmzaiy9ogEU13ADF+28bS3ESbP6Tc2HyhTS
4ryaIVuom0AW6hncK0srze17i8hEUWa+C8Y1zt9PL99mrCRhHL/7wpXd+cO1RPxZZfwRX5njFvYk
8h2lh4wyrcYD70fQpcwp+GAhhk8xBlRzOlos/cGlXelNEDBhe+sDXagrUaqqV6ODQHTG9/bfFuoJ
GHKUU7uTQSPD1U+VDCL8/H6SjkrolgDSXSRuKVxxnniiZlvWITcaMEthw5Y0Rani

`protect data_keyowner="ip-vendor-a", data_keyname="fpga-ip", data_method="aes128-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=39760)
`protect data_block
aGBun/jiuxi3KsznCcY8KQm5BYlcAoie5/N95mvNEgiXgV/YBWGq8TojIhvXwiL7qQodPrC9k+oY
buDGJ2FUcwrsrG7IDkzek0wW0SUeGpnRznenTVnC8+XpQTzNZe1FdK1B4zYDvrz/++vTfcaFNGxD
xYLpbu78QLQok1oZh0imRzgLOWSfrOgCvEztrViqpPz/Tcg/9L4EdlVx0H+/fkRDD+t4zNiNyH4O
ao9i9hgW2dJlyj/cYncJQ0z5QNA3z2kipHtAL5qnJSrU1pzxzkelnY3RyCD0gRbmqPLDDf90x80S
hVdnOesnn9bw7HyoVMg4lqx4OKIAouCCkVjz6cbZ1k9KaAM0r74d7LO9hGHw1GMuTtlNFzlsEFHD
Ru86C4RzllCKNFIEYtNDHw6R2yZyvA6Qbx10FEThgu9wjZHWlrKSHLz2H1v/8pWoTeHp89oJFYrE
QBjdcL9ngO5mlnLGD0zKYwWjazr1Fk8wx0vuv2lLuXxQRTO9m1Zpwn3R2e4ZXn+tsVll//1jILbp
yqBnwoXrXPIQsUYGOm5bx3X+41TzxaT3linGWthIqXNvVfRiB+/6CLxs0vijn5/IVDGIqD2gvR1z
ON6KQFTWY7k9mxZh9ZKnbJxNlrPmIOO3wdr2i+JOjCu5sRc2vMwJGsOvnWflAzwGrkeZhTI81anh
k0sBamb9gWhrV/48ilmWw09R1nX14SMq0jMNAjuLJOto/XxdB5eJaJCq9osVc2MOZiLM0ojk8frN
r4L/2RJrjgITpZ0SMUtnrejFF3Zrqqr0uJXn2bseIQk0XdfVTrjt2JJDdWEPA82tKvizI1e4qRxT
AUbKJYMubFgz8STYxl+Qs7B8BW4DKz/P4nXzf+wzqTY1OBpGAbr+a6Ak+zTROayjtmG4rbCANW6/
fbB3BwQjsr7kocTr0N3HT+ot0zzS8lgTGtyNvJz06NNOPq7vBE95KBequV4WGWHLns5eZgdo6H6H
60V9u0mSiJZpQEHypHzT9avs7/v10QqxTv36TJJZWBM4idGELGDSHkSiPQJVlzpfR78Ydo7X5dhj
ypbs4gKh66u1A+9xFmicAonTcW45GcEGzCq7WdxuqK9JxO396+IbO07C3Cyp3XnTU718vuxaVV9o
rwUbrsokNfR1GnKtkkgb4S6iVvZ5P/SNQ4AyrN2XoZJt55PSuJ1CAerg/h747Rbot2/Rn0gye0OE
LCEs2H6hetKFA08YkUbmIW9UDZAQcMt6ZrWfPty4otDPOuTtzkNfXJSyl5EAzNIWP2S6xzzz6i2v
8T/WDH8lU9u0+KS6kb5RBTNjyhLKaXgydmphXA3d0GogDzAPy0biwQ/j+HYOFjfmDLBgd5QwoW2+
ZTuzWJA3as6duC/vt7P2pzqYcYDCExydXCBFd8YWMXkdE/Ut4A8/5g3I87QeK3WRwqn+c0NN//H2
o+VfBCIzhenVMvejQ+for1MzWRE+XAw8X1LKi+iTiZOd1cTwT4fOSzn4q67FYCAhz1PGJO05O1I5
rzQ08o4kNqrfQhrljh3bdHg6ER2XlefjLunhI33kZsqwYmvg14GGduhU3YfMN4MciDdfwC7qms2+
UlhqNphLUrN073N9ryZfBjjRKTB5gaoNgrVDgc/v2g+YYkfAHJQ29MN9TddNrPOFNOKcyY6V6JLH
Sw9+2fNtehVnfZ9gN+6HxYX6wmNidplcfrCuMPCrpxzRHFpe0lNCUHGjW3qu4Rm7/sDEq1wB2TK2
nvrRpiLkPby62c4ChLePvdzjJ6pxc48cb9hua4aWqmXeWNqkDe36Eq1Dp+jFJRJ+d7oEh27EesOp
/eagsvBAfkglU6jsMf9iRIkihLT+KaiBemjJdDG0b4hOq/DCVRmg4WuS3v1EtDLZsZ3R7g1nz9Q2
otJxe7keE1XSQXv4TlOiZafyLQ5+/5J7Hf4KyzzoEcpkVJgz6c4TQPEjhnWH0nE77hh/+GQzxIm+
XrUSgLA5qxN4FlRIe5FmTX7V31dbnig7jvEErwX9j/t1/7TevKsw4TX/yumhvy/HoXF2IIMYbOrF
ekGYaBihWLIdEuSgNCB53zPsDqsyYDUK385xqjVk0xy9qPxWmtW8GsY2Jhf61xlvtDnn1Vufuaa6
WuDWWQFD/Xh+4L9g+USQb/J2uBb7i8UUvnAqcydN31KfMklPUyvTRCP2CuIluP75HUb76OMqmcjD
WW+QSjOFCnD4LKyD6Es3e1tPU9fNUZTsdOshFmnE/ISW7pfaYz28GSqoD/Vu0FmC5p3f1vOH1yWL
Ms/ifyTn02JF7GduxMJFyJ7S99BYXy13+LV6D9Pfd7VhZSltagWjlsPThiGj+IAuxrmjzmm9qnNq
tqA82m5IZ/xnI8YOaPoL3UXlQq+KfRhNMKcPNSWOOtizqNDzrnCYTQmkRytmlAAU/Og8kMEd2drI
YjGvy739xp1L06x12Zwcs7PjgccofLK8XRd0WaxKJYxiM7aW+lhnKEh7aP4cJ+p7BQk9/s7zsttq
aTcBDuqF7LNt19uhx40YjRk/Wrlz8QTCSbdydN8TbDRKcZ7/I2cif4SUGsWfOCoi01m+rnFX0+WZ
UEdXegAyLVZSUDXAVpH7pfAHF1vCtN4e3IEHVBvKp1zxCZxellnvSe5D7tGOtxGYfwdHZrDUrQ7Z
5c1Fm/Kj7aUKufSup5jCsdAf39K/K1Ni1lhlwjCy95C4EXJj/3gWF4JHZBKHEoJdMWKbQY4oPTs/
IW0jhjOIxQIcWdUVt9MJ0ImzQ4+kojfnlSv6ejC5NCqbd4HapAdDWX+WW/AnxVCeVw1g2mpj4lQB
BSog+tstVSRMrf4wVnAkd8qXUJUjud/rUxlVMZ6jyqQJg/RLdJBxFcfWa+QaAwm2o9V21dJJinVM
vvpZ5hPt9pfIYfaoupVJlXmuIisTFLU2X7LQHc6itKuMWcCcJRpuB+SdNFaO0CEOGPF5QTLF5Fns
G4iiP3T0jDT5PNLsxe4XGMB2uIBstqexJc5jvbQueOl8GcUrP9SjMdMnFtBhROetqRqX5/dHqE5B
23Jt5YixqGM8Ou37ygN5OgybkvHGYfLIyYID5Mp5XfyVl7p2LSSL3pUyLfRPT5ErCUMfizLIsYCA
8L/bEjxKv8UCe6skr2ttKvXb7o51l6IIC7Ji5y2A7eJxbNqvEVX7RbY50XDJOVKXENENacnjs3Na
wUcMCy/HLlyD9rYeQk4bbPB0ahXY5BuDrYcbL6Qh3bA7IK01YH6USjJb5AMdCq4NxOZKZBWBnYbC
7cfCZxglMdaUx9oJj1VtBvoaFi4UNQ4AfagZPwoXl2sbIr1ZT0+NUZYT7jcbrkyrRqg25tx/vSJm
JLs0qvUbAo+sOVzhq6fY8gvXcQ5cY/IpKGBlJPktrbymXYJ4g+R7ebLwXQkNtmF8OewVHJvC3S3r
+URukeaNa2Nn4SV2hwkkNEVTc0nJ9r69pyzhl6LZP17EanahHD3HYfX2K8x2z51+xViUzeKtPKkW
IZ9evo0QxaNnoeb+6OFBR3fY51g1/ZNnhNBGmmXF6K5npdn3sJEFsr3TADnk185UbXA78z0Cs/QW
5XBj+b8r6W/TrlbXf6F+6EBgerKd7sdjLNOFAUL2SgPwOTeYRh0taSoa0U/gmPRCFveFUAkTRNbL
VVGx+bnpdDK+43OyF0Hsab9rcoavCU/mpgiYqO5mHNYyKdYuRj3VK8phIodA7RdOD6onCb8dRn20
agXRMYHdKndMSIifwDbqC4bk46jNek8+odZz8eAAOJok6jfU08NiA2iOM1jFf9fjLQ80ZfEjfBdm
4P5CPVvIbYlxuR3bNjUD+jtz0svQMjw25HSM/unz4r5XFOULnmUvu7QwcGU1EIxqly+Nzvhta1sr
SbJ30tNY2/fIfo/aDTV4R8LKYwaF4iiXt9hzvTEpOHIdg6QxnSXT4bneLz/vc6EiSLOpUmvwHMam
PxWf5ReITaJW0KMuYQl4pPZVWcRRbVHk1BdFbkSTGYmTbUSUgYjSPyhKw3IYJD7RNAR2LSYyCal/
MAtAGWnamaZP47SCDg5a1dzMaa8at4/6KU1eotrA9adJ2uVIp2yt3umlELgJ7TAenbzyutaRnDo5
TGVQD2xIQ5xEQ8QjJZuwEHyxKegRL3eb9CQp6MiCAE07oc7GqWUkvqSgkQivyyDmBAVGxsWxfeSk
sndgPFbk+zzbu/5MGOTsmJ5uoJUKnIf1ecJ6BMoXn7xxT8D3i2ehmQitw1JK6AomF36bcCPDqwtn
hGm887toUP7Y/f/ox3zrPs06j+lNMdUCqcEKO+7eo1mKJeTpQPw17iAPT8EAl7gLIj2Zyw1G6d3b
pfjVSDcADdmKN1LZogJKZRRA6ixm6GyARNToFYdww3Ge/GpjIsd+pwJxSBcxXsuQcPNtNtuacvLC
8RNk15blJszn5Y1xOJRojTxFyt3eWXOsD1HCJSUa0VxRltXAsqzrfeyIwhA/SSL5gYAiHzTojmF7
2uS6J2gCm4QB1+KI9rFB0cFA3EUzKiWZ2GG6Gy7Qke9BcsBa5CGwCbdfRr1u1WLgx2NGJQZToqQ5
0ByFzxsCm1RrVmRexJc+HvK7fig9Jqe5t1c7bspXyN915HnmZXHb3BN7v1buZkxOxXEAgvIrBIbL
UmvpU/ybCxs5GnUjdZGJxkK39JNs1sC1cocwfopThdUVbSv4TGppyxfxH9u3oJjyGKjjPUL3sc+Z
6fjNs+OFFZ7ewfw8k/pH9BZGP0jdSq7DbDDhnaG3MlWIGDN5gYWklGmRmvxDGCAAu6V9ULWkk6dW
TzGB/78Swx/CT00pMYNVR79Pgoypt+8w8MPSAyiC1vZrKTTBBMFC8vISxFJlzrdnaBM0jAjOENlJ
S7BAiwZT5v4g+iL1zIC5KqQ4Vxv5hrYssdBX1Yu7+rCQywfQj8mVH8zlp1t+UxWoncDoQtOujfAY
RAh0y8PAX3txQmMyPvj1uB6McE4iQU4N1YdmEO5ONGKX/r6a5V63KFg3vD0+YjUPwPwYtr7zJrc7
Jk+bkiKNKKFFSCjQr9wCXbTiDsCPsPqp9S3URPRiFy49oEF6wVHNsGUzdqjapDLbTB+buHajgWBI
yjIAgA9O8saH7Jr51wnFvgZflRPTQcMC9qPNtzPOEbTPIqHwWnG/qmb+s1HNv4OfZ46eVlbIYPOo
fjNx6NcAjtkxl/hfO5O3LaePL+5oTWGnlFZQEWDgdBJeSmlId1poB4E2FMqJujVaWmT7nqX7ucSN
ZWxlZ4OpcqH8HgOyaztGlsZzFBZ7mo8lLhDXMgNQErStjW6KYgwxZ0UnvbXdjRYrQ8rUecR/vlTO
GKkO9OX5OHAZWxLCg48oO7xMGc2fn7HDmXDkRCklU66uEGfkJk5Bz7MMAMdk8Lf1rAkmVmZjTENX
mE3pTBmhtk0ljG3LWCYdFg+KgdzxAFMFaYUznHHfuWHWipx7mZRp1dBrTzXiTob2SQuJpNXVMvwW
eRqhO68MDNuYMpMFhPh18s1hm7yCXOZHxwIDy7pd9aEpf1Pep1oi4wEDWG8YFpq/dLlhIiVJXZSk
IvrhDmgG01K6gavxy3jxDyP1A0Ylfruxyy+eZjAtuZSLfPlp63m49QIj+qFGPCdvUk/FwJWlAGat
+KwB6SAz3xKDC3tiIWS9C3g3AdqBspBBOEFjSKwZMCPWtxe9kpd2nNq3BiURc2RCNjqLPXgcq76m
wKWAONsGlSJIJekdpbGYdxRtChZArBV5hhVdv25Px+hqybLNjM9EwDr7PFDF7Po/nkoEgDMBuD2S
v+XDxDpbdy50mpS5lAmIxXvM7QTjLu0XQYhjiWmtRSRM7Az9mpuhBo4NgIBlXvDPCL0dXrGEvj8k
IDCElNP5v3ddXfCtkYU4U5qKRphlF7agMwYNQCMvF2JE4Kz5tnZvsKyfhKtrAd+4rjZpZ1zutpAf
x59H06DqYi7A9MC1ajMiLaHpLCs6lPGia3+KCkyL9Fymi7D+oNm1+oD+7og/zRSon7BaDFjB0Wf8
FpMDMKy2eUu5MLjigskcnVDTt0XyF7TCxxBtdZ9hHKqjDvaHY/RC/pXuVcTm5dfWArzR2Z8yEsLV
IREw1fzcHZ7Syr2Nryysu79GNXFn+uegrE3BYztpXa6rLWYGTqYyksL2zHiUZdpgEqrspsR576nG
o94/gLCR0fXrOyFOB68/0kI0oIs9okyVF/Ev9cxm847ArHnG3Iq8VSTFWOgsJ/XKrC1F6UfpJGZ6
OrOTY54BVM0t1FHMC5cieuZFbdcqMBdZXEwHdJp5OF8tebeGP4lboSyKv2psDUgvwUq1rsMfVKcC
3SymmylOrjFNKx7n9mjSoCEFa+0rJeYxlxScrCUyNxBjy13dFLjFQj9hR+XvAj+VI7V2ITE/Az4v
JZGW2UmzLB6DrclyXG7e0G/s9XQnJ4G8lqiAfHnx/yuHCmQPVBJ7yyOTYHkQsYBC05E51+und2w9
3QNsrwRmBAOYccXCNb0RyMlmyQAQQxxiRB5qoR8UWgmSgrkC0JJ6YdQ/k9J5tHGOkwgfEd/AL7bL
SlG22xprTw/5YhnikQYKavj6UjJixwMdDZTdtT8pVUaDwX1PcNqBtpgUoKDhNORl7Fj5fS+uBOxx
zxNLhxgvWVl+Tc33aNOEzmSGWQKVtWfYBeFjf2dP0xB6nMxPl6UBvmm+XcoqAQliNUtjlCQV12F/
WRuwD4DW/CnR9j1gZQJk0MqdbLjt6OtQfGmhWwbqSOYc5sq+a9/ZVuRtUcWK3y2C/TYLSbRK8ENk
uw7RWMEzOYTGfW1xu/a+vNeuL/5H9lzkIJj0cVtqtSDOQ5VuSeHCgpySxsYGzpBpH8C7D6SNmkr0
Agc0YwtGgnf+hua0tM/++A9PZowMTkVoLUAbUa8vNjw09T0riTwkQPW9/Lo7/98kOKDNrmcwzO4V
wmAjYGYX+WLYccn7LnDHru0cqsiykbGrnPQQRDCmt7Lb88uhZTMRCDWEj3nvGBKpLXv/V3T8iJWs
ty9V+jljdKRxug0ii9pOZp7Uk5sFx4wGaIKAxp0vMtS6+c8HzhNWBQqb4+tRBSpreH7bxjzzCjgZ
oE6XmB6e6RxxE9/UNNqMMaxVzZzikeaM2rO4I639t//hSAVPsqf32Z/ZHVBsGywOjuJX1msrphsb
/juxMTqEf61+rvBlLmiy/VFKMq3k1XObPKhC98doaP06W3MgXlVailvhjCxw2+Ln6I+5T0q1k86N
4PmSCQsZ8x1w0XCPqKVXeZ7034z2GjW4wtiMrvtq0UVa5YV/7IVewPaLnItrGdMgXlII+ci6kpH8
hRSOnWAzw9TiYcDB0GXYboZKNDP2KLmRMPQyFEVdzcuKzgE4liu6Exn0B+DPWsJ2P9MRt2nLCRAx
xY7iCe8coxab6SG+mg18KRDbLEOvBrf0DqFfAjhzDak1+9TVnpg07ZeHKaTIZh8Oq0cGQ7wIAyQe
/foZ/0BYY3T2xrmrsQeGVMQtJHN7zKo1O7GuETlQ69XnR+AymST+PlwA0IULw6BfbZ87qpU24Uz7
jxF+BIrvmxtr6t7PQtwJgmNuC2Uqm2vCm3p8AEGpuP2Pc9c8cAX9h50b3B7czrVeKRuv+6DlB7af
Ch+2hjJLWqjtOuRmWL/XCsieXeUlm0qjtM8gOZ1U0DKOzwP9nNcT5D1/q1h82fevKsAjpnzqEfVj
FfldbV7qAfpVojUSBiNlFS7yHbx3mjyrwQ562MaHgcEcB84CL1SoH7IBj65kq/dT2czywTJgkoNr
w5XPhk+2mwfViWkxVIzHWIrPXH5P2ZMHdlzkUmJglA3bT8hr0+JlzD5IGmWzl300duB2o84IVtYu
kfQNfasAK4W67yqJOV8Bu00lfHHrT12nNWsbVKwQxNDvnxSU1NlDJ63NaBSnSox4afwY0YxkHGqT
N1DRGRdPqhhnnqDGnSaXqDe5TBRVTgr8qhxDa176DyfK0qll9RJ8NWN9DO578Jz5a0XHT843Coqw
cIAaO2aGrcpbdhrIMiNSGUBXIomsX3rqldJ2q+YAkTVuHBwfxzlFfI2YCpQtCspRjYFC4AwIst4l
IT8zQkYHcmYpb85spWqjdO8kIX+b9hWEt84VtnykbdM/vSzi3qTfCopMQnyjJM/bF6dbAYA3wRnz
Vqvpp45zij02goakkq93S2fSh/uyU9Ax/8T/LR5XUzu0GbRZyFFfiEWDI82Kcv2Ism/MtQNK4U/0
EHbWgiOTmU1XRXw5ne8eIkxz9+2aTMBDE1p/sm8jWf8Fn0fxgUQCMGaWvdd2KCeJtBO0FNtl8fFv
eM+ZY7cL/FJivovmwHDWv6HpwIYbjhj4rfOM49Y7c1YWtQ8RG2BjhSCi6499kKHrAec8KlQGf79c
qNcl9HPn+5Yi+uG46OLEdXORGzFa+zBbSfH2E8JkV+EjbUDFnbexS/PY6zS6AVFAt5lDLRmco4Wz
swZhpFQmmXuYzlSkNrxeoV02B9X6y4Xlf3+k2PQcJrz72VS2F1hZ5Wu4YeKnf2AYeGzy/kYNYyg/
SP8lnSAwO7SURKtFAFkXcdy8t2ZZac2rBGofOub3iQmg1c8y0XdtFfObpEW7cPB8WBqWIIZf/ezG
P950HpfNSi8zYhqy5RCX/JqDZkEveEV2AgmuFPwrZnbGFMSj6vS6ZqdVeswdSc5L/Igm0P4ry/VL
D6HDARwpQE7otHmQmnhPpaKRZlAF6xfU7weOJgeiXBnBgPQWxlIq/K7D3ferg4j137onYLN8W1QY
9FmjhEqDDZtEEgBskyH3+t3I1j/OoVlJ9XjHVDZLxw3DyFeIlgxGHow9kkmeX4uFqn0UKyEiZfE9
gPH8mSfkwzvRquBk+jIZbfHa3SicZH7+oHj8APb7mJFbwXoZjhNW5Dd6KgwROVWbCcJUaV18/LzQ
YVOTbJHP3b5TKKESPLjCljutsTixiE8il71t6V2gPg4wlRUIAp7N4hcTAGOdnC31YuzjMj1u4JUg
fDhAldeKcRXhM45by7MRj/XccJpkLNvE9C/nVI2N4lm3ot/wwM/NW+Z4y7k4kEJhHyxLlY5EZygn
MXcaI/BFzU9rOfZSTDhCpSDmFQ3G9f9c7SVSvnVM3AEYoid06F5/Gz5vWSrZe/+3LEn6K28gkTS1
SuX1Pz4wR8wcg4y1Mn8fcuM4S4NnKqpAlQQKxNq04ix/FGlqWK34OHFuNXQFBFaTyReIhFvAV6G4
fuXbu8og+5yTR4O0lciXdLdbtxv66r+coxetWa1j3pcYfi5+h8Hll7zxwyZSYi7t1Y7zVkmmuqWY
P9dz/tte+yDch4Iu1iwfpvxd8LcBrpg2NUxxLF4tZkfeiYyp1M+WG+x4JgciPqSrcnPK/XTu9ol/
pQIpjJTjp/pSQ1i87sk1bzavMpkFawRBQ69GbPRggscCrNgs05tlM4lF03u3K5/UPgA9mRvzzPA1
ZwXfBLVZPpkVwg8VNv69m7Z6lFXahTJCXo8U406PEZEdRD1uYWBUkdlmpqpZWOVOm4VdtfABR2I8
/r3BMfVeb469VXYlbBy4g1Ygu91Oi2IfnQlS9zmh9jR0pnqtu7HCXZi8LSVm0e+AjOKhFL/VDwgh
2G3zyUUaQH4IOGPiCyQZgqVvTcJsN+atj02QLXZVEFk1zoggxPLyfW78aqymZ+8QfzIXSsQKXqD6
g7l9+pyOVaJgh0XRAX8A/HuNT/omqo4Bwwg2mtuA7BWgP7iYOPr6E01rsKWjGX508NE+aLRrDp0c
8e3kURe1OR6EvfOuei03+c/xSAAtiY5fPR/mxcgVSkx2Q543scXwOwM5i2zvJnrtTvJp6jJnBzYa
3Kl1JYZ2eRUuD6cDhMpzWIbyvmXC+6jeWi2REfBZCUmSaVCYKUXNVFBSHbdS3TBPR2JhPrp/6wjH
gHt1ZxARRybtGKVoNKy5lMUWW55KlSDk7AFyJhRdDGVVpbyn13zL421kMY5pQX7c1spFdrdiNkrS
L9HklW3yL2zL+Qg60lMa0Ke5uSzAx1CHlwusoluVmlD0IX2wDVS41wHicTUa9mBy3yBLsOnew19R
aw5Sqx/KnzdeDlpNvYAgK6+wmMMr9vyjyaZIIAz7WbY2+YXSDxF39HCWL02cYiIflEqyPj70fxVD
eqbReJDs7SHV89jviQZppWUmemHqwzQ39DU/wbGhyQWGyUZi9Tbar3gghrZgYWbiWTSv48cQVtqe
TC8c1/J1yZwCd/SNjnAcLo/qUY5XSw/sexF4CS+idJqILuEyW+XkP1zdKYk8XFO/dPslleazCAQA
gMxa46NxLM9DO97c/LjAV+8ze2qMBzJR7EdfQCCoZ/TxHB6oNjX13YmyWesrCbDFW4Cst3AIyBm9
TGmS5CHNTi5VzuWjnbl11MmQqxbIsuUWfvx+GW+TRcghaDV56757vDDIAldxU+RrNFzzM0syY/7G
70T9z99bDMqCHvhU6VlCyh0Ipt59/31P1+IrOgsJib+7dGmzmdg4vsuZ3smdIFP5eV1q9dN4a4H2
nyEi+gPnMyqQS8IhrTJSbmSZUS7oyNeH6ClpUv7AZaSp/3lUijw3kWNYY7/IzUYepAw9kSezRpwq
l9LNp0KAfC8AmP487WWwtPQAofA47Ld/fAfFv0yK+wDC7clxog43MNcIcsWOWbg/gA3dto/hSq5e
aRy7AujnjOkZJa+/iccvVM4J37c1pYq2ejgyUGDhLlb+cHvGlu5hXG6USjv3u33p4CaktmXM217O
ViDBhk3SfAf0WJKT64ie66uIWZNQKFRpR8YrMoK0EQi+4l7wjNZzwL/vlw92KPEhjdjZuPlFEm2t
ag5H+e/hH041IMdsGR4lCtTHgyPJwZrAzYSsTqvFh9q9LQJWnwja1H7g+u8dcnhhuVAsUUJ+Bjcy
zGMQ+vgA9/dmSVyNXefBUTi5a7vXcsM8VGpDrICn0giNGo0WXHWT5Cukmiht9UuXRGbWaiPdArxg
JQo3cWutDfzgZmOmt+JxlgDgUgFhjlaa1/N9p1fNC+M52vuJxweG7OD6pfsxvtuzqV3zx9YHe0FF
jJdPpBz3LGNtaehyPBN51V68y9yAmirRDavzk4vXih9UkrYMFReMYG4sCbipX2+myrMccUJ3GYjm
gMQBIRrJs1z4rx6Hr6IBTgqdGhJGJrIzaJ6XMBCi/MSYr0e/9iF3LsoApVKZVsmuiOZTA9BiSIDO
HbWyuoExlQhnJQhKrKGPBSVl85YKmAi4gpVOa3+EjIIsmzqKj334guA4a+JB3rv6iN5DVX0A9VxK
owHBMALA9wFx2QbZTjPB/AJOLqZim9bNL2vLRFq857EXhQ1Ftm2QoP1gGNdZg1l4iA4nvN6WVEcS
EFTFYcj+zu1E5tyI8r9pGt7Nkk6p+t1ZtCRgJC1IzM//0qlR4hT+2a5xiQdWdkfuTgiXkuMIhG25
wHg8sq/YtQeVQGqurrr8BjmYtRxTL7+W1uXuS3+SaGaB7Du/2BgdV6rb8nykBVKarrBIoIEI3ZC4
sJoYjBWLW+2bIb6bTRSjYuDwx/npEwSgdK3pHzfG/wM6/AIZOc9YYs78adnbNC19m7j4KUNZXUvm
4+ZH5zLEP/ift+g1FWPIPh5Jnp9dhXrRFsVicKGkhMmdf6K+X6G5sSNtnrC4hzM95Q0Z21XnHuq1
whZm1x/JxdCvrBH0/BURjIAKPvH4E1fqmDhKqiGU3acQgCukyXbAiXMhiPVDBYaMnAb3uzcJChDn
6QNo87AKHqHFCV8XIxeTIY/OX2udZGyOW1++JNMIVXCdup1nF//org0V/XS3aQilgoGjVckzcSOW
NyFuKVafISL4Z0Lm7imQ/LvopMLCe74e4zQ734GEoiUuvGLI7EIJbMH6AeRIxV4Grvf/jfPtdB6P
LZsyLjzhXt701NDNZ3LnWxnA7S4XfioDr4P2QHgcpye+Nc90YnZwMSQ7AHfxKp15J/OMynBusees
ZWTSfgQrSbevnBZXCuDFfcHJcvwlZ5tpXlg/ngoiLyD9kNtgtk6uAS5V15L3+d0lw/y+VuEYuKuR
hnIU07NuyjCQEulDc38Q0W/9WUgvI5l/HfurWTelZRcJkjSlM6+/x3VTJXaHmlqdVfaoAoA2Rbr2
J+gtBQ8t7tmspfciv3EkXfIqFWdEd/soc4ZAgkc4rk7GfxIMCllKdYoo+4+YX1CbZCJwMP3FJKsJ
j3nWrzdmNQkt+KngV88tF9py/H9d7mKwulM/kaDN7mnKJzTf1ygm50yg/dQTTOe0aBrNtaZ+b4P3
Lh70v0D8FOfMuDNuION6HQ599CFmAd0ty9WpfCNa6DiGzBbiPFN8aQpAIv/DS7SG5NJflMgOsNRd
2/vKO9kgus+01MIdzReHKYczMmQ2hneRUe4NRyWhai/JfSKewvSPPk62HYtWZm78fTR15vYYDWC/
RKjJx1vVhekb0dyca7RrUAiObNhYzYIiaeogmTgOCRPkLQlmYdF5R1cIQsLLYdd3S8M0N2TdsOn5
BCgRUdhMO+Of4NetW1XLH+bXbicL3ufI9jotJTva0luUgkAO5RSFmqLCR9ZuMV0IkSXgDeP1HFxl
Za/VCcM1BadibyHhUyFyiLyyY0RfNCwl6bG9UnHKPmPabBoUp7uoRGbn5iYLqhBMPhqaUlHFzftC
GhUbxT4YomQqmx1LKo3SnA74lxi0p0f4OAgziyWMaV1/Vmx5pyh9Uh1be6qocFludzbQHIopSb4x
OwnEcCCDKZf4tHDzfElhykLncLWzuYq7F2owGVUmyVmfUF6xyC3IlrrvEWXQ69aQ0fw2M0MPEjgW
nZdwgNpLlrGDa7cxXkzwLSEBW4Gz7GbqdBakVvgE07NsX4sWmsH+dgmVV57VLhYO47VcMbqh2lsI
0RVkaVfEVPzhX/7cJUbF1rbCfO45QoyIxd03oFlfz22SD8LRfbrbP4I6q7BcIlHBoevvIdfj34BZ
un7Xojoh0ESxNQN8bRZvT7xVUAMQftkkAfBJOiIlFi/T5MxWkXVWgvIh8HfunXl41qYDar4qA1qH
p20mH5FjoVVJPt0W43jYIgEzc2oGuJzxpZOw+wLEyphc38ry/uQjzhiwzxrt5T9VAFHe0U401Cj8
4PAJAhkUFNnP7D2XsJcLqnQhdKSY8bNu1h8NuyWqpjurAekVV4LbpstPfRPd0JIVZhReYX9MDWeH
tt3Mq7PCjjzFWsdfTq0DK/ByR2q1V6neUNQ5X3kgP129NW4BjClsqaF0bW8qVwXHBeFmaGA2i58q
uS6+qAj7WYT2YuXlo63OX1k9C59qs7oHwlzSPn5/baa+B20PCibqIoEr1ApzWyu3Oo0e90EkdyL2
GHwBxxzTsB7YYeejIU9A++AUFxkMjJkeT1B6RAkIsjVsw8pqL9884YiUzUcojj45C+jBm9C1n5di
l4ZLamzluh4JOBM+fKRoSGHgTTRA8NtfIICHarOIUzo2dkwjREArSnc573JTXCzywOJV3tzCKRcW
+CXmd+nYr4rR5VsHy2LNphM/ckW3/Fj/oGlbM7soe1dbGnI+I+ZaJG3EHXvE0ceKx8jlPGCzo0jI
5AA2QT5l8qVD0qPeasDyxUuKCev4IuHc3jcfj8LO+U4cxUTFGuzL4nKA+kXAWdC67EU81oCMM8mb
Q+SwyDTEXAEb5Ka1CDoxgcPuA8oVfMjANFnp9up2jTdUncORxeomOSn9H5I4HyGPaK2/nhdJPGVy
ygCm+n2tuWDcBCVB1SzvT8bP5Yjqz+A/eUYQdxEzcWcFF7ZlUTbR+1wrcZesfisPY6T5Fd5MyfKU
YilFi9AMPx9GOd4knTJqC/qJNd1m5bCpZoTRlEtc3Hv7zhyoYogOhkGD4R/1Q7bNnUkiNhygvkzX
Q/s4eIFfjNrbYSJNDJ8OtS8GwcS9zSO+m3OEq6QsZdEDui1JWxgD6kUo0fVpsWVKJPgovQ2dIaOp
j0FKT1m+OZzPlVPq+Dpjzr4Oe9/umxugv2fU4YBRHvBlgjXQWa4IQ3YwHl96+CFPPhX2CeXXKla+
IBMdpVWYT+yceNIdaKrXlB3NHMJ0zzKp+X2gSeXNTjKLSbwQZ236iPcTfVIw+TUWZJm0R//uv8Y0
pqKd/z7mryJ5izrQAy/Xwn8DKPF7bHSpS8ZX7zFhL+A2rPqO06uN2G7Unx6+LUOnYQ9KeAh6ukdr
5N1n0bTzoata5EXACC9i4pUneRhvOQCYxqYEyadp3ih4AI/8Sfirvd2VvOXg2b5Ae4DziJcM0dmu
ReT7tFqJo31DcsVc66MnxQp7MsAPzcFWYwAp8LfoHntzhfJyJwMXK4m2Xo+U4N75fHX2y4wmowkE
laAPEtl/jtzDrHInamCpwNnpZTGYLvb39Nm6XgYj/FueDA5LxbpbNAilHnP40/78qBtEcfwmzSRE
RDtf3hlH2JI8PsLoef9VXhIYz2SZhYqqnN9Y5X2fPVEObUURtlTeFBoZ9D5BecwFWcehiFEohcaU
dT43CcAXEhH3o2aoipVzbG8ZCoc1qBXL8N5OHKLHSBjlRquG8PHZgYPJ2NhkokjFOBH1BayJzBm7
tTQjUViDqmSKToCWnXaRSEiJf8zzZP0U+LoVyv0AGeb0xgBhamRMN1lcq9jmNqjkmGi88TJIYMMu
bpMU3n9feAPp37tI0FYUL2Jj+BQhNo+Ho86Le71qxlGwNfM24ykRYFicQ4yiU7obQFTSsc8JtzfJ
34m549wcSgDaBtiJbayxJFFkDWWpu0rObBpDmMyY7mLBTR+ZP3pHQ0vqAS4Ez8+IS9pYPSRwrkN3
5jY/YCtmw3W1Qc3J5Z0zihfpDZSVu00fNfHLFGTvSFYr+1hW/eSg9tV6sieMApXnBz36xPk2aGco
Jgn0j7T9roCivV5P+5YbNlVwHcyytJrA/HBh7Ki2G5v2lSaLaHhT3yHbvnBREYh7bHShVacG7//+
7lb515m0z3Gh2OmMftMkRFo8oV0mUb+pvcSDxaHQOA73Nrl2h6RxwHJkyBm/fbA6L+Z2GsqE2B2N
x9zlSfQsqh/+evmAAxOkMIgRX5jxAWUJnjZVgbIuZgX22b99yz3bg1gNSciA3jShrC/ETBhcS3d7
RpdVunebNp1cIzfOkDs78NH6PH/bXa5i/FnQfDxQrWaxCeSmJ9BkfNAiddZFZ/QlQRCbqib2W2GV
Oa0gz91dPTHssxku8FoYtWBv2HiABmmwoxvG96KM3h4wY6TKbl9rTtaNVB2UgYZbeu442lMLNKk3
Y7QUub/bPY3foUqdb31TL8PJoz7AJFLaSSg06IJa1YX+TN0FVxOAuLYCXJ2iJXiBxoidRscnx4jN
DeF4trz15xhDJkMcWxVT56Enw+O5hs3/oduqI/AqbJ2OvO6TXqtQIMgqdGLcYPq+rKIhUwVIjfZC
KOo82mf0jeFj89aHXlcuNLkrnbGhy88GyuumJWHs/HBhvw70oGRJxwsmCXOwSUiBE8TXBAZIxvbY
tYJXWJgJ4KQ/BtvlI4XqC6IPM8slcsVhrtMEZs9cmBsc/oHoUbhWcC0xYnOGGOJnLIXe3UBY+NDJ
fbn4k5FiHFO/GLQdoC6u7tBslXoK7f5AFmLjWMV0c//s28X0CrhgUt2rZl81g5UXIpjWoF4ABWtz
aUltW8NL8+zz02mTtWjVyBOEQEO3mThHRwk+Lh57I7aeZbm1lJRfvA236zeajeT0QEGLq9Sh7Qby
HilCsGBYLCmNIz61K0yFR6iqLLM7pxHK2ShXq9Zq01TXbjQpy5EvKPvFrSVgplldXTsAlEd09758
/JpkR5qLTiOugHfgukI4kscjpRQH054VfL+Iyzpwbd2mir3kZxAOSWsy6klFpZR0cECC1OfLFwlN
8YQEKtHZu9sUT2Hc3CDH9KNa1Fi0yx4FMdxuIz+KdXMsdbxRMxQO4JIybnOU+YlUj22lO92etzLS
rR7PlJ9CDd9tw7N8LUOTDxlyzElWD9SwfbCHrWSggGoNjUWDsY3rv+hoR9fDVmT/LoQ3ou9APmh7
+0OxZLfTuas41ybzgiHfgHivMNy2W/lS1otoRqanFQhXNOccdn+CrztyfUGdChctRdeuSRgCbydv
ObNzZFWw0A2tDKjJ45LCHJWTizW4O1HztEgoQjzyt1GdHmRpJ537kQj7rbW/vAWdC0ZtHCGgf07P
GgBeD1TL4K6AnzaRg0xQSZOU9zVfwTDTFnFsA9HzPuCp6L+ZBHrepL7lc99yD+MYNjdlm+hV4Tw7
bjFr9cTBCLQbltbbtnXgJ1eoNkIlz3EZjtmHykI08BcAKBcA230/CH6JW19eFi/CUqCTzalABfSs
LNuc/AMoqODjaUFJQX8ooXkj6DZ4WAhNsJ+lOJ6FSI4hse2t3F5ReeRzPkaNaEUZMgRMleN5VU+2
tQmAmaXSzDtEt/3Pu7U6bneg+grMDo5OqHuhIWsNHgo2GkcnaVEgxDkEWU9tuAF5MxNKh1zjDuyl
deQBUotWGzdkvaPkFpJAfI6xtLZhqmCdJu5sfQzgiv0uS3v5iLSN2yVJzmXiGLDUymdfOZ6C7Czb
Lu+iYIY9LEVzovOI/bMNvO3VBMwdwvGY1sfbtz6GWM5xyYULgYG9zvOJH5gicOmGPkY4/JY5TAvF
/hnn3E3SuWhjEVlKhlCKjIOivqZs6HnVNQO3AWhL4IPptsyoiXtbfVGnMaRgjMaDvFFzwl/jmA5+
qnQB03JGHCLQ6Bxpfq7vb1mjAj/pj31XZpQ5Os4ehFppeUTFi5PlF7aL5ZOkK+ZfpaQneqMJoxJJ
A+FvvgitYYoqVraGtFKSyOTK9LbLzy/dNs/96HaVSfkgctvjYAsoF6yc6F/I6qV2wmfdZ/7NLhcm
5lQGob5iBDJVrHBSVRj31PXQF1osLWkGWD1kp9NlQgUyQPEsqAvdh9Q7BR6eHQLpMCMrOgQ0Za5h
AFX6I8RFWkC5btWraBykNaHGdpq3BhuYvEPVEnfwVfHIVx+su+ySrpNmTlxFwb9PoNsj6+wLFqX5
O4tVTTtBXZHyQgTq1Jtzuzs1UmjjmByfZHMhVz0vYD2pIqiaU6moAu8Ts9OG2ikL/ohoVBKr1qMt
/FGwTOEkES08gcYmcFbOLd6VcgOswF2iIbzhKRd1Bev3MmYQ/unhhzY4aAPIz6YhKh/1I0NbOCXI
NrEi4sD/wIIcrv9/7DvF0B7NW4kuro61EvoSBW/K9NdC6oRaLCRhibe4frgEQ6HQjPCAFGW8PHKR
Hb6C+Xxm9hJ2hHI/LyWu+ja/yN5JeQoHhy5hC8cVic4VynvGTHQ2yk0XXtmoKWWgyZhK7440Rwor
+5LfMEeJAh1H787IdVz7l6qjhF88zoD+8ETNFgZreBQjsuTTWoUnhp6TMnzNU57Ofeo7txstTI8k
8TBcxf/ru2xEAO25otUt7E3IkXjOzRJ5/yGnW2L+QHbZ8vCJTWhl6N7f1s63oJtlaXgELcYhpbgx
5/LJsTolS5QfDRLvWiCLpW5NP8Dx8HY2ye8noOd2SUOMJC98SudrUkimytUiQ9uH6h5bamgjuJPB
IBLbvSp2JHXVGmecF6uvw9MVlcT0QpjKpwrn4DCvIiHVMpw6iOGZ72M9tvB4+Coyb5nwDGJhS9bn
73Mcd/8R8Q1kTmeF8hKFGo2e8kzcd4iY3mpR269h/fxENyv5ejpRaY3CACWNp9BXsraVqB7lws3W
ln4pE8k/cJ51MgyxwLrzwldMGbc3FsgrllrEwLyjOPumDQYaQ/b+RxjFSAVHc8mHzmw50uSp2xk4
9v4YrfIZuCpnKI9PBHZhzUTxS6/D2ELqu/krRG9p02LFn+UODcwjpSIZ0znUkZ3JdsVupzZdI/h8
/PdSJfw5pH4FAvTBSDoah45VI6DYvpPKsIiL2WMGebXRe07dFlVnqr2p2vE6JNtXOKq1d2GLzp4Z
awlEeVf9R4Hr1Ac3D0SnrtZ+Nl3gptvJvRYnEhENXHiM2ooU3PWKnjP0cbg/zzllbCw+0CaqMdwg
3rwoqytqVu7CODKcvSJFyGdkT5v8OkYr3Mm9vboHKfkTLscI3u1KWLIiaa0ThBgmrrajaP/gK6xv
kIqv79tPDOevMZushi7O2B4TCrVNdTpWm2pHcvkEA8Yl6e3e/klNqDq++sUrrHWWX4/bHAg4sqRj
zirPLnl1zwGAaCwJEmXSdhws4qBmWC5OrszbXwVjaTSazFAj7n48ciSySEaWmOtfwg7SSgKLOZMi
LjwYjH0YkPGC+BZ/TOgcf3kZANK+yBmyXtO8XfdeJej/UhUUQPIOyxkxB7smxxZjOD3Je+hM8cVe
nilUjo8EEoPJWnN7YJK95QSIcQfHGjQwNsiMXdOa7Q8qegZkh1pJmYDY6ATRMt8gVG2xWeE2pWet
z2vgBCyDHb3GF9gEh9aJs3msj/UJTZ4WQa+cHB4UJbA90Xix7RTF4nxva8TYIPDn/m6qjZHQ7DXL
Avwhjj2hKYDi0n+ZwcAugjnsjjexYhXeqj3gI5TEAEA9K/OVxr3vfsY4VvoIczbakNGIeW/GHHVb
7FFp5pWiQ57myMKQTw6sWRjO/Fgc19Ft8b9Xr4lAEWuDi7DOapEsHME0uPq6XC1r02K+fa5oxBQE
+EyocGlYn1CI8NK7y4NmjormA+z48obnQWDSrXCI8ZJXvD4x520QiRVmiXJQh3iiU7iSLZV0Ei6A
69k+4h3EgWUAN0zTJEPYcWhbcFYKOpCcHkvcu5621CnckvTcreKFXJRqsRPz37TTRRrHzFV+uk6k
iCHs5XBhIZcoCFvl6shEZlRof6L2BHsXPwh6MnxGfxWLgjTWtRdvW7U4fBKD9IVhIn3woRBlgFCs
pDqQej0eAhG3MMov7Em9HMFaJCIiCfUvapj7zItiMQhKLycgxXHT3tZ7UcpYjsrBD3vReqQhjPVH
/TpD4nx/wUn9nNBzEBu52s0I2ItOyPjxFgk26clvVaoPzt3wZlICY+b2Jw8OKoe05RR2D+IibqL3
WPxTEVZWZ3zAKvRvNnFJpMSEtTrEEIgya1vFPmHsD4+Jp7wYel6/Bzagahl8hNlmAjomTwmnNQUb
ikvoV0iilSVKgxtFVxoA2J0xIexqSaPlG39qMpFFiy65Cj7MqY6JxZnt2Ssp67lGyUmMuXgVLLdu
STBNL9fy/1kYZj5TPdYliFGUCAZp99y9fqlQiBD8WCPSxrhabU1V32E39VpIqO6q+qVhDKhSLUwM
EGU2dBHmQXLiBVHcwxmONdwTNGRNAbTzbkX/BF92IYkloRNwg1/PUejWXvFudWiE9gG3sN/1GKbe
ZQU3lDRebsygMLnRonOYywXbLGgZO7ntYa/oclolm3YayzfRdg/IeHu43xiB2viRawfaWs8lbP+q
j++VQnBTlVprKSNq+44dDPbtWzjCNqmtyrodLGZu8KAsqdztGnLrQ4qD315yI5rsIcUdbMyI0wxB
xdwqEr6XiJlU0X7Q3HHGrfSOesCK2f9m+FStEYw/M2zP9Tn8KiF2KUTUPlZ9ljFmz1msE5dSPvgP
FL/gEPs3mioSAtPdvHLya8LAqX91SNU9317tzQiH+xO05r9vVZ2aNOjqJ4SXpWtvTSRwEzmRlm+X
V4S5tVx4UUhVvhibRl/j2npRQjIlq2rtD8AxEYFcTTwLY7nkbVyTi7GzBZCx4QOuae1w1C65yGr3
+MzLZnNqcX3xsrdBlAvUL03NyAriSDgbw1eXshn4JbfPcxN7eqWscEoTTmYkpWmsrzB36e9d8psu
WvJx4gym92TRJ8T43QjuKLr3dk3esa6dwiXloF5kSvH2yorx3JxEUwY6DZdiSeo3x00k0Hngswn1
P1z66m/YeWjI/VsuLE6uN1O/9RMOx29oeYMPuiupCWHQPFTlEimAEmCITwCxCAxNuEDEp1RbTYA2
71PH5E/zHlRxYqrLJD3csT2ggQjr5yn71s4usuxZ8o9LrwsJbdZXMqpo3KoVGrnzpt7rkg6nkT8n
LvFP62R9Akhlw9nN/SlD6hhgXm5Jam73HWlTeWpicCDBMqFGg92/seU7dyH2/3q7YwoATHaeF+Ye
YonDQwLtkC/msojaWmyUEaWbrodCA9ZUGpkTivxTFQObj4U8Sdmuyij5Xa/Z3f1zNQ5iLWXkSDPk
5d32WvbKHNIgkNUYSu5goLcYkYYR4kKAGQjyD8qnq6YVsaFu3xXlCWMDyoT0Pc+MVAoWMMHHFeep
HuRCKUP0Hr9Egg/8psqDXQF5u7gpI9OUaj//Rc0HYBFy9GDH6yUqJgqkDYurAHVzA1wLZvvmvv2h
x+vfHAbvRM4aQnf2Akbp5Et23k+9sYEZYM+RW8gFOAULAgBQ+6OFpP9Cj++vvTqWKspR7VQW4HsH
yyaFC4A3+fW+5Avi0KoMhnhgDhRsNGPy0tjrtcaDgAXwo3maaR3nS3myB5tdJv8/asowxDbJ11ec
qelkvjkW00HWTOxVk8tpDFSRuXO4q1fX1Nz1TW6G0gqV1NNur4mUsmDdFVqW9zBWPuZet2ywPJ8M
ck93b3/OmjvDudOs3GFnd2m9+7zjMWy8g3dbo0Zo3IiIomtvwjytHFvj9JF8lQ2f6Qs+MU24Xa1D
yphWB/i1BS01TmZaNbkkgw7LgfbhE6QvU1Ri2oUgpfYdlyBVBgYXRn2gOyLp6FbTAXZ9mb/5Lb2p
x9UcXrhz8s6jZoplUOInHzRlxkegwhrDbbcPclakbMNB8poCBupmMcXBZpu5c4i2ToxfSjGJT8lP
6esrJSQKjudQpEGMJwioBkE0RVMsVkpsaAnDioJ9XtXZQitzUYMUXmTj+oAttdNSsNlN/tNM+bKi
KBXzwDObqmjCIaBRWiM5K+8dhb6VQ05b7yvBdXGKaJ0PCMnj1Al31/I5GKzvQTnJ5sgT1+9XmqM7
Kf1V8f/IrsIDBuyqQJ1BzTAlIX9XSVjGJsbTnL9NDZaOL4kYEMUFpV3DLePEDO7q/m2fV2Y7OLJ2
NAZXuNpxtEQ3HcD3WQvGe3rA0zTXNJf78++Rk6jNrYDtdBR2I4R3PpVIl1KQ5C/NHXkBr3Fgh7el
qkXdeFiGAphy0NCfksXr46xBKLZVENX+fq5dgYHDYFGV883xPgGoB4hJ0GAGKEPQ8K2NyKBw5w2b
jSAQRQZwKd5wuS1Lk6XTgpirj2LEizHFZp03EVNyZWsNkRUlYRJQXhaRUzAG+slaJhKKUEt8db0d
OL/OyCJvEhsAL8+AzoZLf5CcE60z9kHh11o58sRv646WMG3P/V4Gj6qI5jsJk15MOdFX4ZywZl6H
qjbx4fZ0wwG+rShLOpK2w5Sod+nr5mC1lk+Q1SI/c57bZxvUPcsZWrZTrr7+RApUhTWgJjt/V6YZ
g8jT2plQGR9MUZfQt1JSm+P9snXXfhSdeD7APlzoeqU62fBfHh0HNS2Gx+9v+n9ludfIcUdejOvf
D41UVPzxzqBeKtxgVljz4gne7ZQlIEZBQ+yELYjjogFMNMefegw54o0+QkpODAuURJaAGAZ1tmK6
SkSbZW1JwxY6RdVY8o0xlvkEiHX+/jkSCPABD4ugiqzIbFhbJ4k/5eMp7pvJJwqqv5Sjs2pi8M1U
GdRYO1UPmeeBut2D/RLk0ld3XMkn4fm8n7WiA7bVL6HlyoKjOj0oIvY/KFQsOD6kEs/ULuaXWzbW
GqQixEagVDW/s0OeeFYGbU/rJZdL5qiQJDOqFdfv75bmzLsXHWEzmrDXP6cwqOZFJr/8pq4oWeRl
oATWHzlQ25FB2VC2sZNhYyUJksCA14kjNy8quoaaUhqhmLfLLM/x6MX2UDD4qc1qSdr/fb1t6K7J
6sdo3VygROFLM6Wgy4HVHZ7gJW5xDyf54R/HPBXgJU0gr1Ze88OdRcajT3wJIok2YEYi1udeccMF
r6OBFJxWR+Atzh9YtcxHEklaO7JOrrVJT4GuOoLeECln+QpD9QiUAcCMmYLNSpbSW7A1OC+xPRYn
Sm8u3ehx0xwEvmy9EeezQyjlLCAOLXDCcUSCrdbLZ0QbcpmXMByo7x6GqsblnnpG9yYlpoQRXjWR
WSqWVTNEXEKHo7HD2mi2G2a/6Hf5rdWuEdj16q7RIX2zMStaNWzRrRJqU7XxhKB6eJEDKUX+GkDM
S5/Yf6i27+c+FrZBG3/ViWJxPIlE5CP+zgbN2BGsH9Wzz9Cl87BqP9LgxOFePRkFPpWZiAGJE99g
xupUOF/kVFiupKLyxMOvz9G5tcBeIMQZ38VyYCKVwcPGhBltwGhgaoqI3lGfv+wDPLoLpsSOEiHg
kXOpppjknK4kmC5Zf8dOLBaKqXeiZij0Le8uTK9ej9Ihgt59Y8Nmv5bsVMfHLIcj0MS1j8XKmrGz
wxB1C4gAapdIdczlmNnv1MxF1++Pg9C7QXcX+JsfEUjNY39JXdNj0KP8+oONWlXLfMW1hcVeHAFz
aaybiKpsXSJpvl7kQ+9Tl7XT/8aswnuOvsJbicFM56nrkVr6McSyqRjefjah1TT2K9i4vpFTM4UQ
EpCsKJpVCaSoNUJuGeA1S2ElZRZ/HbbFtJ0a89XaPbzsdmzAuGiRn/xW6Khl+0MkrklCA60Qv46f
acReGj8C0T3Ml0RFRhVgaFbYt9/PrU2x/kd242Bi+FmhKFGW+KuJQ3s+dXBh5JTrxNtiSCVj7eY4
d047um8wi8lV5A13y8DbEZO7Q8upbRyIxRNAw9HsG9udI98f4KUMcNqZEz+yhDquewdWxifhv1ig
zeUCaK9WmpIGKzijbF2r6jRJYbYinWFPrqhX2qkyl4o8KfQTRxM1C2emWx2d+e4dDdHocGprSR1/
wUvfLFvb266KlDrUyp3hcr3OzhKNuY/ZhBYXlNmQnNTG6pxLaIAG0M6fk2cqMEihMYFXAg2ScDih
nYm8e0m9ph41rdeSwaHLlejl5bvcJHQan+Aad7NLeWC46HYLwzQYkJzATiQKzU/Io/fBYt9xQxDK
S943/orvP5dmG3nXbeuGc076br1oN7o7YDdw+ezqvtfeCNJi+xg6W0vjd8kCsSxKWAgnF1WGbTn/
DZvZr980UR3ko6v+Eyjn96TUYcBKKxC+YlTgrSzIxVChPQgV7t3jiQ71LzFl1cyvTOt8dbWv54Bc
ixuGK0we0VWMqYUNpMvJE1Eit4UsW9KH9V7kvmu67D/qEBZgxRSlgy/8wl1QAh5E9+NRs/4lAX4C
NOIDtgj5T0miaWaI0ajGlWnUB2UafFArQCN+1u+mlE+1jzwNp9/ECDW4nPgxSBV5jaofmbqroNnw
12zrC8p63W8TwCwdWBd4lIDy3aRU0Zua5oxwm7vvZFVeu0RbIZcemtxa2eddRv8RlPUX9obAgA0/
0Eo/KXe7G3zX9KtGlsNUtrvKwWD+wUpGTS8Wbosz911EQgEJ1tdFAumhWEjbLDc4fcpBaqhs/aIq
aiVOeUnTnSBqjwhNRu60YpieoeScceVH18oh6UB9XUShNgQwWkG6rzqyDcRlEQCtmhVNi089/YOL
WX601pGN01LLQWwdT9nurvkhtNQFDU6oh5zrpRSOjdRNpAElKy2yBTyOF41gB/LKm/e4Id99wREb
meKRkeJUI2jzjBRSyb58/6UuV2P3DTrgxbWqR1P2IvRbG51kJfyBXv25RMzbcmKDDPa2Gxf2UZlH
PUHEO7wnS2R3qi0bfPI31AYsCaKRpzgzGZO7R+FIo+hLXi7M5FcSUjn3JpB0faYosF6rONDjFeIG
mAOmYkV2Gqnnkffv4e7/KObmxSkvWZ1mhpAa/Sguc5qgltWBc1xDnQBhHz/SgeH4Iawu5J1aEHqe
Xcklnzky2eq/knAQWpx3tQMJ4zyEBwnnMO4krqiQayk4MCMikilCKDttC4yX7+a0RjjpRo0LeR7p
yOCD3AGFL/eZCXAX83oWEjJmCXQg53a2PC8iYHI3Z+tcQlliuLwc4mMcx/LIuAm5dxCQHDty1nTn
mK6pYO7KLj8tMTmUVKNKCpWumokIhpyeXWLPDqC3F+CnAwFZeIvvbSDvLvPnq6L9ZYawiJY3qygT
AH4UDPdPXpGJTEVY/GSNQQO0Vm1R/5Ru2gHOzgSm7h+2qpVwRZFEtjoB5MLpFeRrnVs1Z7yrIbAo
DhUQft3/Hm/ruNzyvLk4j1AGMHmVVsjzE5lmDuaj0YABxThIedq8RvCwdxnV/r/RvKQZhaEvd/Hx
DkV7iAv0h8H6NBkZM2jUxbgACDFqhyO1r7XiGxZa3Mgq4I5s1lNDPUFTtvn44hOYfx7K5ebX2d4c
mjvsx9gjdPom7EWoMwiRj7nvJwVa291sFHrkCuG0GCuTb8zzcAUUpUux9NQwavukccAXX8L+WTHw
D6DTeUJfuf5Ix6PGy+9SVgw3BYjlRX1+WmIkjP3Qh13WC4RCJkXFZH/HgLgLmqnJ8ujj8KGopfit
e8FCIeh74vbQC3z5wtetiAuEGm0A9v3lgDWZL1cSKtbqKDk1u/WQPHTY8Z7cIbuCEkdhUBswaJlw
A/jUVkgrxaAP6dfM7qZ4mlN8m4sq8MN00oaDJngxXX074curTDOeY/ejLNzGbN0U4Q0FfO1vv+NQ
9Pvvcy5FYC24hodrfQZQvyPRltun97NCzg8OIUavIJ00665gC+uS8oZ3/8Ah4dtdyOfmx2A3I8S/
hA0doOae3iJ7im7ZI7xoUPzGSW/jr95/v0AwcLeSJvAbjpQnw5BA4uHY4Xg/9XjqopL3xU1SNiOo
rse5RObUo62+rv9t+haxB9sPqf5dEeRGl4lJcDw3ei4dqpwni2/hb+Pe4oNnZqFqfQCWm0DYIQYN
aTyefQc8f58TxfXulYGkUmiE5hiWqyhJyOriFXOPaFiiWHmUsFYqThorhEYgpbAi+dln5psfH/aj
XQMeleKL7ETGPXyWGcfb+aGOCLfO/sOXCwaToYDaP19bMjJtPOdJu6DkRb7r/YJw3ekO25GeGwIr
X3ChJtkRcWbmezPxSdV3Mo12ErgMUTyttPQdeoVvQQ3MlfSGkY6/EG/n/KUGIcC14POAnAWV13Nc
sn9ZhWUOK3LYcP2gLFWhCFi1BfCvGjmUy6+y0+6J890GPV04qE4dd3mbEZyB5hiXVK3UlgS5u0eE
CeD/JWaiBq0kMrVd1l9WxFgwH3U4+TekDHGeIIQeDxzauZpFFAdyewtCAam0N3eY01owzjTycIXE
2icF0WQ/ohwgq82hb++sQG7iegqdrjuWWm4WndvAM0/5c1Ib8/dhcFA2sxUER9oBS37JwupnImNT
BLjnmy9cj/DaBpiOWBHb0tAIx74XQlR/6t0VyFWB9Nqk5bsTaAMGQ8x8kw6R9+phiHlDnaH2qxEM
bjZHQma1SkAKqfCc/VZ0+bMavHJmNBDJU+q8gUw3MV1n855CNRKYTBhGHxiAe8MIYNn9ILpYmXfm
yvi54SNq4uzuhqtNyYWUfMy5bS5/RUbBpnSDUh6BP2DtBXuSa9LXxSQowdRP8u2xQURU0nwwXIyP
7Y5HzlCDHnKiyaB5ogxWYTmH7mK//zswr6waoGtbDxH4UXEG/y41OEaeRvZkwF2vZLCj80TQC0wH
d/MJclDBoFsfIVfNwiAqa20hYYSMYNv+EWznf1jKXreUw8uPwifmDINT1F2Ii9vPnZQ2WekGVmR5
1ZLb6QbV9mrA6TXLzN5CLJttwUbr3nTjep66cIi+CqqMRxrKEJtF3LNe9ldp2TuMb7Odg6GRkY6p
WMoTGzDYXGLJC088RYmmhts662awgUnZbSvHEb8UvTjAhCRhN6QuO3NTkaaQeMXTjIvxtccl4kHg
PMFaN0Ia7kM1YnXhy/cG2bA/362FgKVNJbKXH5oN0EZ2UgdJNfq8nwdDc7pCPoNiQSbGzTCNhjs2
UW/037lwsEKsjRo9+0yJC8YEfRVDL64p4I1TSB/gM6fqDGVzgOLOMxjydQLaTPbBWCNdHF/76BnT
Lz53xKuceg6m0B/SoutB67WSbdiDByIxc3xuhnQIX3gf4PJ16i4SoaSK1/MSmdRDKsgW/AVIf5dD
6JRav732dy7ELh+XBgthWHUn0RGIdNylQRw9Bw5UsPCdyF56qeDRdx6tAacADa1WNUakjzUNXnwf
mmpDRl21Ty6tXDxsf2FzfbUB2rOgJI/OpZ7xfYpiP2FLBgZkK9C+wf94G0WT8m6mBuOkMrQgWDiB
4R25zPZGsujCqKLXQwe7siEVr6qqbZ+dRr0/O29sPMEOBhYl6/N6Om9nqn/C964lT8mCZa0Y9Ek5
EMLVEQ6yi+4tY1PT9T3GBZ2cGUwLjRgqi09ltQaylaBGpLMecmVyCRz62AAaDbJ4qLudx4wQTuE+
oquLghkd0ipOHYYOLXnU29sA1HNj0+4ZfgBa+hawaJ1d74ATmCqFd2sPVL1VKegmii7yH10Yxtum
EpUxhDX8ovbWGHcXE89RuSf7tSOB9a3ArmJ1vS8aqPc3TSXC2WNRg8gWV4DaGU4N3FifCttyo/0e
Ye7yLO52UxeOq7V1pQqx1cvldEaOnykrmB8ZXrcXxQ9rPLJ9Q6cVDhlaPFaqkpNii44WuT1xXDvo
qMvVuoGH/neqozejuagQVXA6pt4J9VDIkFH0OErieKTUN3i3kwMuR8ju5uJ7kdXm2zt9tRUrdsJG
/BKBW/yC5X/PLc5nHHKrhFu7wvgq0AaoIzStdiq5Bhn6qsiKxwNBnwWYQ7aZH3vc7nZJ1fH+XgH6
AKtrGeW3x7Dqdi3TpHULkyGVX1fw+0mCBJJoMUhGRldTCpDpzNl9nm6QuJEAsbhTfPAfbkWtveR7
u+vBlhFFp6harrTHkYJJN9mZTNqJAqgPhAwGUo3xx50ThsIACMOdz6y2ePG75lGdIQESiAe+EdkA
Bh9eSNb97Xtu9C/tFpOQwp98DQU3UupkdKxVwq1yWe8i4tI7gMJw93ro57aSitxZ4lL8hKmdsFXj
bv6JdJ5+0PRmkn1IQ92XJ/XSe9C4JSnt0DP2Z6sWSiZnI3KdSADqtvDrZJ3xSDs3J1e+JiAjSALt
YmNmvGtf/kMlIjY4/iITaN7EL4AlNk2XhbyUZwjChq3yV7ToN1oqldQUEeCVhRI8X+sIfcjvvWlq
o6cuxyuUPcfjULchYeF86dMqPT74b7I9nunb3ODbJfmQXxbql40Entj7QOT5SmWJtCmPicu2C64+
3fjGTzLOLaEJ1jS9fEDXZQv5NaMSyIfHBBmY2YhVBt0immbVkDDZgr6OvrpGtxOrIXDcTIEJywjl
LtGuqmRXZcLokhIW3bXHzfbIaGMWMBdSZEAqa9ze2H0G5EbqNS9HQkvlfSp+fBUdKXDAnN7bTNGl
J6uTDovirPXzvhM5h4StkYBkdsl6Bg4wyCr4FcStElIUoGzjplUBsQZmG9O2gjoFidOhACSIQGaT
pQ32YnsP3F5TwJmq7ng6+J9F7p6QZp9F3+oTeTg466YXybqn4Yyh4mbkVrCv4swi2RKpUzkL8W2z
b/WhsS+WOG9PN6uFw34Gn0Eksi33Fv+DWkEqp/cDg9yLY8urM0zJJCTkCYY2BlDrVfsEvLulX44H
KW9HgcnRdH8YVv7leJfkVHy1uGLQcfh4vH7dbnAuMegHuxBaNHTVySTsO1SU3l2RCzmLfYvjuZaC
YLs0tiXcXcmYRfRuyjQnoikqEKP2isYh9AowO+VScDb+RvwyXDRM0iUWspV8KuFYnlUrw6YAp0xF
g3KojYSEoNTaNAPxDqsUwLiXyNfgK6GCPlVpqJBpGyWz8HoOeUWx1ts5FbRGUupKKpRV9ggAi8rZ
XG3rH4zCeV1Qkp0tlcUpXUo1ARjFa80Qs5UWjx4yW70sCPYUdLT0rhy86XJYsLZj/GmwE8MW5Swt
qO611raV/DSwq7/CdpXEze/lRbJHpDTE/trGRhaLcCUGKb6XFKDdVq0qImAb+GFYd1TAY6mcVh8o
/D/BT2Mb37b+/pBYKNZc5zPoypdpSHESWrDklU9SFJzkh1517J44Xa4c9QCRUsF4iKgipe/lf7c8
tQ2Q0i158HlmJ7y8sJpRKaUcTyz9Pygk2XB9FcW+sRKK4zb92jld6WXJZc0kq2n0FxaQ6UKmBwvJ
n7TRLtLHZOZ6uBCKwigaok1MU4JFX95ihrAiZtEjztjYP6pGPYWBRkKT7C/6q+rDp5UsJJwdFsqC
9sF1aDAJhtVQJDUBl1YIYBDzVB2Yo3uzf/ABF8V3NV6U/47ZCsJ9W4xSUtHr/5qpPUiaFW/u2vFt
LFyVXHRmeQ3HpWhcKG7TpKzzQygF7mYey7bDcC4RdXLcfEuJ2PDy9BUEkBF981BZ1GZVMAplFMgx
Z7DQTOFCvt4PT8mIKk4oaAlP9Dcae0Dco3s33qLYV1KdKvjrOqaLRGq6vWvuUIa+XgqjUAbl+yqA
PRGhKfrL5lXArm29o1eq//gGuFfvPkVNf8XooVxK8HIDyEDWgcC0IKEo8xe3q3WSGJ7CvkTl5SEQ
S7eN+dUhbe3l8tUlYmUAxO6kmDRNwEDHN4etsUgB8pKmmw9cfktiZ4573YjglGYGn0Z5FkYfcVeW
bh6KvUir6IOQbgf7ZdnZXVgrYU3tagK0VjrwlCecQNfyqifSFYsF07aLLaPN+xtTWwC/1yWHTwgi
y9YGuLzj1Hdvh55+F/e6cJ1stDjlfrG7jxGzXcP1psYHym2hUvd1onmsadfOeadac9wxKfMSdWjg
ediPhEX37KrgupOOY7khlDIXrQVsvmICxKL9/yoOR7p6DpLajqM8Za+/PSRCsIZOMtM3dZuBqO78
rIcPBQ5Nh9rRdJUeITGmDXZjUv5MJauzeeXnvAq5rbpfTV2p9d3AlTVaY57Gt7IBG5TQDP3EaWlV
m+es8HS2qMSQ7QeBftXXZBEasWStus7UDFnhpMUNWOPk/IxYFk8MreeJtjlJa7revXI/pnI1/w/Q
VuGkVyrpQpVcofIJUm4A4PbFL+Ft2OHAzcz3viKiASun1wcufXwQ1Gz08ruonXktSO1FVOppRvYB
FDPHOAQY4cKkgBMR8LTUYBKbZOsPlPJJVJDkCvZ9hzAar159aQsxgtEkoteS1PyWHOzjbtiMRVFx
mBkg1LjlmkBVnWofgFUkE5pYhrju2YdVemt3hHG1+AbyQcaaCet1DriEfNfzTSOa0tmWckxQOauJ
P0hvwSb3jFgWMXoEF4sWRbBKpRyrMUACzYp0kUMGn8+KClHehgdvhk+Y0pZRGETqDA2Ti99VXuAj
UbuoM+htdY+X7kVES0cJHnt0q+diLeOA6UbC1r2VSwsBsXeKSGkAP4wG7rVUh0Yb23ZVAw3mENKv
HThNKpBTLJyJq0esUe97Npq3pXvUPmsHDI/TCfZXybnrV/eG/pZMWUttOQbEaPS5reRrevRSRivD
WZetkYDQTq1494Tw3XED+ZHK96c4y/u3yuWNJvAVUEH9v+2zABisSxmEuRPD5p0b58WJfvw9bxwM
PnKGUcR4mb4XG0nfLBQ/Zw05AltG+hNNK9jRdAtWDTV0uWAEYAST0evT2lwK0reFOqEIvkepiBo7
qquMcZoo/PReXRuMNW4WVPVYnZSIA/Er7j7JhvFNgvpUDbY1R1uGbGSE3Z6NUsMmNoe2UqDWCvry
1UtdnSUM/MB8Gv64XhPaqdOAV4luaYDqD+RQGTRKSbYX4Hc6pCm/7S437mm1KU+ejNYKikQxiIYG
jj8XGgEHEo9tHCNwJix1RYjOklizdq3jCEngC5avCb3tSK1S62UBg297fDK79CZyNYLSSvh1d5bN
XInp0pjX2OHwvmqJNw/HAT5DgNP/6PEhdgjVhfxtGHkzpbrnQIbSI0PIttapXCAtO1Qj8X93vvit
ptmQ/OO+8rrgopAGKG75XRDVVNGXOEbQ3Qd9O2QBsI8neSnWo3yjlhjuDOZ3DI74V5kOVq1cskiC
xCwrM45KSdLm+M0MSzHbWEG2AmXCp3GJF3njsmh15j+WI5y+8/v7smpQyagxvKlB4dduYgrVWOR9
alZr37jnG4RavxbOJHLIgK3kh6ucozKVqSLkDAb9+QIRVlKvEVcWyrlefhPulml2ufg/ZeNgoI0B
SzeNTjKbC52qXWke9oP4H7J3h59EtFh+ApFLwLhXH2pJoJen2K9P6SH1U7HEIX08BSvCh4Kgh7Qm
+NRWCVEYxqegFiaM9ZOc7/wDGOjv0DNvDBsWJztfGgIz3466EeYpBQ2/1PptGNcUcbHewDAeoeE3
07poU+B9tAB0AUHmLR2to9pQ8mcYKlxbZJiWcqLY2ozRcKDMQ/uYegJvfvr78NMbmosnSaCk51im
AmVLeRLrrKZErkLd9GEjD+HTVyiEr87GGxpZNiFUoSVhxaeRTzX06JcicK8guwd8WgrZoui2MARW
XmLb99PdMBPliV8+MGcfyN7dBKUm/BHI+hHdhrEi7sDZ4Fp7DLQDtJqqaSQixHaE4eeWQWpaRWwu
eAndzXvYnIT697zssXbCBRIVT26vTj7Jm00XkyRmluKzCCcJ1Att6x0FudEndKalMCEJ7rAgIiyl
rfwkBKOG+VopXNpgtrrW4EV+k6RwdTH/LeH6Fm1ixgwlnYZ9AkhPfeZ7BZ3atu7zka0Yn6WVHjor
jo8govWwguz541VxdnYioANtbzW9/okStXjALC8Sf++XByD1M4H2FNW7miA7L6LNhnzmqzP748km
NlCSs/I7UkDoI/e/LmDvvi8mO363NxZNTvSpWlEcvzX+BnBAws07qPi9tgIHo6ZMCJ8ixS5wpYRo
IzPTDveeoWuZox1UvmKPe52+qeHuygVNBXmXeme/bRZVxJ0PQ3UYyoB6Dui0O5fh5ubzZ2qso9lo
U5btPemKmFAi+zhp0hO2bBcYXVAgkvL6l6newa4OBj7IbW6rbcKWzUrAIzddr7Ma4SYU617JYGrp
vkpG/6Hg6p0GfBsB97pRl1vsgl+rOOm/EW80pKIri6nYIuGyqdlT2z0mlQhEepZsoLAsWSS1xVaz
0GX+lhRwZPmxHoVrYOmZ1IRNWeoSGnuaT6FornTpDnpRS7qY/CzJfnwPE2R7zRBWKJnJTmz2ZRtL
wEYxvQW2ffLzkxcF/GtMWjr1+gjfnK/WiU8S5H27z1NeKddSGSAV88voc2f8osUmUBweGFbmJqPZ
nSSmVQaUsXUbSrVeSX34RHSfVwF7y7jiIYsuIIpY0R8J1d94bC48xYJhQHtXTRoPX2qf9O5W/gD6
1UpM5zhnntxQxzAY5+Wqt/JdtAK/yRgmfm6hSXKRXatR8foxc3Fdp+l34p8i5os2AT73pRETzfDk
BKc39D+uFTXX+kn5YgKQmHGulFGK0Dh91yCrv7PeTIugxB6Sf7Eezl82bZbJom9yx+kV4y6/8TjT
tS3aE2mMdcTKCj+13XzRKM42F6SQqf8Ae8zBSR0IcW3LJIem81Bim1JQT01UwYGGHo7EvDLNS442
XkTwSFB0HsmaUeSq9HZKxdiFuTxjYBc3qxElnA7p2OdnCJorWy+3x6ryMIrEKIOHXVEzNMVRNfqv
4bW79L5JzLxLoDMcK8bL1zy0TCW89CayQR/fEctjJ0blHe3R97wgnqrZoT6Q37CvYm1jMp1fQc+W
3JEPuuUIngBLDxMF+FhZDlG8V7OQXCBPDH0tz8a94H+K/VdLXvZvWSDwHT4VJDaK/f1KLUbdVIxL
t5LX+2YPBU3cLJT3UgZSM9dHhdI6ZRed7e9Aby7n0RrnISId/Ekm3oTAHRZqIYKQnw3AzxwcKBZC
GqHMzhvHxrkkwxLFqXiMt4LV0f9QEQCDsjol1rd/szUvKN9y8Itg+Dx6hYmD8ppz8RT4YkuKQZ1q
W8EBk38ONr6hoPFRtWXRpVyDDyP0oMYI+itNRJzMzwJsmWcc7j/PuAr9GDdWAzpg+XUyp9jzLe3u
yy6ngegJs16BSewVw/i4YbLXSIoG42HCJRg2Py4zgrU2XMn3UE+D77Kvt/mJZVC3vf0g5GYnidM9
7D8naPfTz+91LSSa3gY9rJfVViq3+xQOsWXwU4GlJbAOdxf10itA9b/8vMSLOU7ErM/Q1aQyDjzT
i/+k36DPLp3rPvzmLe8zMPpgswercQQ6x1+2TvUrqzY0XydqfubkTDk0a5VqWGWQl5sEhXSSLg5p
+kbSAQazs3cx5fCD52eSfFKXgZvrFrCpxrDgh/6PBAQjpE/EktXmvlVJ9El/6mIrVNxFVUILSt0K
WY3i4nusPtR61FWBjb3f5dnPtLODuYX9NDC/2XEtZxKEj3rV11SNaR6pVfSHscSq0yX9p5mLD7EJ
uJYn2cUt6qXcOTK5jdJKGgznOrgNiwgiJTARgGGNqLao+plMvjzccQzyWiid6IGFqsoQl2nuX84q
Yta33iBoFlpzftvYAX9OCGGH274AFaTajI84kGJGRb/ozWbSYi1hgETluyogNggSGvSX+1uOuoDo
wlyjAX0oZ4xhahuhXaMQ/+V+9sHFTrKPhe6SY+m8Ug3iyvMl15HpDHrC8GfB4QCI4ucLB+Rmgvat
yt3AdUuGnNKGZF1GwBRX8ovaTxEyCl20D+iXnGM/5BGvPk9JkJft8xYCRXqvpLupkTgD1B+2d8fZ
T3ozwpzQpE5CLD1A4QgtwlbLO8mkClzG8cSmWzNcfGIHEwvsCY/dmaQuSqWslx6jsEYJiIqQhfJf
PEJqoBzbz53kYAaNmrVhdmDOJgC0zz6Nononz6ydL1Qg9cyLY64QXAJde6yPnBE+8RMhv05Inn0z
P5CFo53vAIcI0383yRlay4cOK6pmABheMK2QV/auZQq41EXkONdhcpug8OFTX7KYQxt48Yqb9M2L
lAKz7zJ+O8pWg2Sv2MgBTeTsZm2lDNEX3lQlqLhC0vYyzOZkP+WkRX4exwbZmuHwtHjuHAdmBoHF
IVzpBom35kCjVJHcRUwmUlaZFaLDcRuB9uxML+G4qwfCpuQJePsDMAHqsawvU3RNAQscnkFy+V0W
jmkVtcHco2GDoQH1srbB7ADNSEQzIHuFNKzv1AXqkdsMlzqGdQpQ+QclOUkPoUns13S+YtqxxJBp
7mzHwkdCoA+GbBHWpwUzrT1TNuIMI8dTw8588cyy3kmsFXTpKoD6LZFxbZYaaUsTKMh1qreu74iD
9I9nMfVZ8IQGcYFDAr5AxqXK9tpBwTpkD+5jmnbGuS0DpQfVlhG08z8lxZ51Fapy/FteYnkPbYEb
eOQn1iDcuPS4HptpT0suGQ76gAcZkV03RyI5Hx4ocs+9AHjUBsl3n4eUSBM87WBsfIDe167Bcyra
gua7lJyeqyIwydtDIUY7eX51oV7v6lTRMF+PlZBpd4ZkHg2BH51jd3A+Bz39OEyQLIsfjmGmvedu
5mGd/RQsWxDZ0ut65nQFQLJ7ER1pOzZ1/1GgKbKe1JK942nziReuZ4JrHpNAZ4tx4OGWzinyd7Xz
wlH9F70oDsxJdsBDUvcKmBhSZDfkKKSbCF28pMEpTh5XOWWxzJ5UWlLXIHWEHsxVY1ewXcVViEYi
IO35i0pfVMq6+8+pWJv3+rP/e+c2qD3tEwrmFhRV9zvBtTpMwBX09q8sOIn441IlMwpwUqHsLXZU
XE+dEqe0bCYZVR05KG3MyR12GC5aK+sbSl8BVlT36j8s/2utkTHCeTrvmXVM+tWYalTK/qGGJtLZ
exYYvigB675s8HoYDHIaoLlpXqIhFWLI9HuB7CteutuP+KT4bUOMoWHhh7BMrcvFydrZCL2lMUo2
s5I/sF4fkGU1/03eLVhDp6uBT15ko1zNKe2qUGxKi+f+a0A9uw4yJIXdBGiQb3Pv8tSOoE4nfxgo
TR2EtXyCf4hV2IcPdYx2y1+GVo6CTMGwlhk8rD6cL9A4RLt/YhLf7zGGfKXe+3Sup07NzlFmHIfJ
x7hmK1uBbGvUU1abnVKDHt3l+cuoJ74j8nYS5VU2dQd3RdklMvtv3BLAy/5qV63nvngoV94cdZwX
5HyKi8b6gTrrCEFCVuIea3xP1Lo1UCz6TiRrA5ugf7lsWU/WXY2rd7ox3eTOYapFXx1p60MJ+Xnh
KIn47Leh7vbWZ9YTMbksXRGZD50QsdagD1gr6+jU5gQWAAdquqxqgS9CNR1tWgoeQFx42o09GG7X
/mupZvWynTRq0C+YrI8R4dym3Tj8PoHiWX3GFte03icnsNG83uLeNXDQ1g5an+e0b0GnNrsleyXA
hzLZ0YFiRx7tEjit/e4Qfbj9W22b3Mn5/6az1jY+2UwuIDfz5slqbV6RDYmpAwTXVxQWNBiaM5ux
ejZtP7PyDRxboeyyvGRQfUYx/SKS3HYGDs+03e9j1gDS19PWWWE2quQN8cpXk3YgzW2OP4wJpzgB
nq7+qH8NeaSNAI5M29F9/cT3g/MBvLAMNKZf8Ev1ediw5iDRcyF3MZ4bXePfUKfp0pM/X+TOEZEq
dHascZENY3rpnLOYqUUF73pEk9Tw+sZRiQKkuC82+air4mnD7lgtwtkL9maMEnwOUk/09Lr5/VD3
JBVpA0dKnIjaYQl23lRx1QNZrxbzIhCsZos1oSfxwcTd7WQU2KAJB1FONYo8ulDsKFgZKnywJFby
xbpi5kk4FGA/E/ngOongJGFOkgWFCd7SoxBqyQw4ze6z3vxqWXptOMj9PEje013drIx7IZmTxuCQ
fTSwSr0VNS12qY6YUTKH2GnN/mrdu8wPNdPNJ5DbT5D3396sYqfNX7sKqkC9a9BhbH7PvPgJn078
vjuDfv235zrG74aHMh+HPJce2r9u1F2fXsR3ynDSkwEzbV6dDopa0jLdtZS0hwdrb0MkUmGafxaD
ebL1rcRTYUqYc9P3OYYldzgCGsTcJ81b8Ug31B0KatsBtOQRsXfGWOrnayYlBHBTi7Q9vzUYri3C
X7xxrtmy8aWbdRKkv92T8RMYPE0jIneDKgYJ21TIU5r0JEk8yiqXz2gmRC3SHh2bWKCPRa/B+KCo
yZbHvf+Y9WDVdJN7RcpwO1h1BKPul9WbM9jEPLwV5/qR49NyTKsGSwIAVpx0tr7DMnSZDPzVimxN
BhUFrC4uDhBftS2HLp2o26mNokp5uybEiYrdWvLAkEt/o4EXny58H4FcH6v6rzsej1BOqi13ohFn
NShCQounB6nEuKWbBev2BxZY1k2SZcZN2e1KFmpCP8VXk5fggZ5DB2Csc+iJ33OVzjZ1aZTNtkD7
4owOlMXO0Ue42WrE3aSHsoCAn5e5wyggmp3TXGJ9caujE5EvB+c95rgI3nZESOXztOfrv9R/Gdpg
0p9xRuT+zE39s+VYqVtZw/oajUBjHnJ3DgVTkGMQvq8daDr1wISA1F7JaDf6cOTt2K3s5m6iVWnO
OR3bBxdxfr6R/XoCZPcoAHY1xT93rQu0fWGUZnYFYXHYIXfzWrPHmAXdE7C3KdcUXrqMKtMtXEPH
ncgd8GkwNho62GrLp8uH+8PuqDWIb/So1PaYt6+E1u38vWzxDgEFJswOwLBImpFR3p7QEcy05fID
x7T7BysR4M8EqTS4WCVfhFJ1j1KSCXm0VTycsDMSCfev5Gu6vQrZJhb8L8Tzd5ztHtLqYRolXc6S
AiBvd3Ut8D2hYkGPMtQMuFU7MImVekTyvZkPQDdHmzgmzs+lSJ2Gw74HGQT758OZXKkM1oXKuLFK
PNS++XA37wMU1iSM5eqzbIa7Arm6wDjR/op0Jv7bto7CKg4PmYRTy9tBkDL5RhaldmtdjVabTBkP
aM5BRRYuJ2WQJomZ0NeWu664qNBFc0KH2GEo7DOi2aqBqFmi+8KBoHr6UNzIRZxnjCBDiy/i1Yi9
dkPv3k1NBAXOMUHFJGjXwLohVth3tkRQEsFNB6zy9RgbA69DLA4ohAK1x6jF1La5j6+vS6XrIVY2
hxS8ympwwsrB1EAY+247CcODt9sJscGsFdgQ8rPeU1zSjJXs49+eVZO4RM3lIqfOG2XgHH9Umpcn
dkcOc6SsLQZdrQizkCdMiuJweIWzT68Dp2a8ibK2HYwR0yXAmv8UO3jfuZkoBIPyXSllXw2u6p5p
lPS1rtaGlw/sqkmw3eprlABliL9pO4CBT9RLxTzzb9DcnkQN+40YurdP0e/ShhqBRInk22NZ4IhU
Q77oL1L8N/6TriFFRl/mAWjex5fBDaFnpUBbF3n1CZPYwHA2m+j6zVLysK9YuoAoxSlxWChBZgTP
UcVUuHelIMlwClT6kIkB7d3qPWOqJdQ3Bfd/cHhLonDhZZM4jpG/Q8FfcM7PxOdZKoqHoWOX+FCm
pjrmKiChcODPGTe2imqkezacs8jAjcupavUCHhJXvvoYSPQkvc2KukezzEn4RbTiueTIMpEIXRcP
PnrntQBYkhb+E6PRkT/YqxPHAK3lDsNn4WtZ29OxNMTAaOYlHYQsC21Re66F9zz2ZSyMYomiNm14
08GPafgG4vUT1oABQm9C4Xfm2JeAqVtWzksom900EbZr7NVZepfhA+1QibHO8fFsxBb/B+X7n9K+
9l2B/ePaw0V+76lQOIWdcXM2VIHoRzhwUAkDnb11HLtwCv9gjzSmgngJ1IMZlzRR7hguc/qtNxq4
/3FTsfbhc2jWAPbhNDHOuSelwRzSXX1SAi7Ega7UF+xofzwU/vZlv1SZ/XdJ9F/MoEjhflHLkfQf
a13erYW7cpdZJB+cng1ZgHI+bjzQ38qokoCUMCETkyhTbOIsfa2GEXQgccSgg0yIuG//+Qe/UIgV
b2ihqLYC60EPaC+IezdCcYLFtQ3/S/s2YK3dpQvuj3Y6TXFpftdu8bb+8nbftROYlgprLebZx+LZ
rY+jqYry4s6ChnDJARD1AoivOwF4cwPpjCAFdT08BH66g1ZxKL+KcnBfngAbhtYBBZM8JIjBWCn5
EDuR+e1asSiNezxC+n8pmkZuFyAYHjczA0cOyjsk8riLFSA2jTTemqw4V9Fy/9gVh9qFpd3BfgpG
bvYljLIMvj5R224DcWfrgFQhu4UlBSsFtYsKExpKJswzP1kz63LbhyYvPhNgfQ8oq0B/nyf9zngH
67JVNmmqvQ0Daw3Zfh4vtY29trAWEmP35WPkoa7A94EQGan2T5dhDtIT2YMqn6NQ9dS0fej1rzi7
eawzB457km2fH0AcxHkby1QZxLW7oADzAkhTBOAJ84lKhcQx4VIvTUqXCpe2RtbkLXvDpTHaElAL
Bq8tvKSyBsSIpZHJ7/U+GUAz/200QZ8cVMtXO+J3Yx2zVBlAyAllCI9uC95tBemGCwlqrECUWoHq
WxV7kFjRWRjHPP6KPl0zSvLuXo9+a+LXZHhQdudOlhiC9LbU+BZPZ9918bfYPOJfornbzLBNdcf0
hlydz/f5T6QLuS+mQdNN3YiSixzzeYdQH6HNArnFqXzzkXWQpRs2Eph4c8G3FqA0Dsc5VJopHiCJ
WMGQ4Uyb6HCRFogbB6G93OMMPaMv9OlBrALpGlcur3LGlGcwmsc9JxWwl+fhYGBQvbFzlgh8GwRV
fiUVCLWkdZMjh3un0q+uS7TZ4HWNBol/743c/1axSlUhqUONUyiiM5A+zikhXwS6Ohqe7EpgOHP6
DkbRWA4638SMZ7O7f+J8/C7i0YhfsuheuGWcN1je8CrJORDpYMy8NBHjv8xa1RiGGhTrDP7SFfOM
RGcqN0m4R+wZ3T2CE4tNh5lr96rlDcavUB3UN2m/5XsCv4U9SZbSxorA7cb7TqbBKmBBWLXpFPQN
OF/8G1t516ly6WMGDCYPUwjSa2Lud48B3qE1zyhZKzYbuQFr5j1L4C4x/598GERwDGeI0zOLscfj
3GhKlVFwDPkcjr1ahHLsyiNwj9pVguku7rhqGhRAPDNCGNKWdN8gIT0QP2UTIS60mmgqoSySGoC+
LpMQKazyRFmz4lE9EjwQjs6bWMeXCal/RqxO5vIFieGVcYtjUw9FkEPpu+fD1YHmKOLulruxfccn
GtOMl+2wKVi2CRMPwhx5zjEIXU+vxHKBLM+Kpl+PL0ZD+8J5cwkx0+10ofmAPFBeBW7qh98zHVP8
7ghmBKRGaiVYO9LgCUl6pbHQ2kCgV8IGJ2msJxar8TjbrnrI0GShrw3Wtrg+cskzbG+/uOSbXbSY
xTvdmf7cZ/9zkMf+NZmt20vGStKJg83iFmsjWo4NlX2xwBx0graLdxwskjKlBMh9pZ+1d0+uIAeN
0gSS66Y8ltdy2/MfVRSxY9IrjuotPlDeC/t1uv6IZkEBWmm+o6qoFSU8s2L7cot3r9dip9KmiPzG
hqZaisCKUE7TJi892zMQt2eIhwzHoQEU2/9hXb6LwF8pC5NRS6VooxCkh7YqA3zX1dsk2dDxxMTR
lAOSPnQDkUW21j16kdovaKLkxTcXP4QTSaSY8pm/6hN1386abPFW95eYkuwfG00LUpSQO0gt7llL
0cZWqzvkgkLiyprnb+bqt8Ids8J/uZArDH5/yw8IkwoyerSMfwc8LUFYi+A2KYek07jrXGBPJMgQ
17Snu6joGpSvCgg0u0lL6wTjdqFzy3voIPrQZl+G1XkaaMSqZis5JzAk3cGiTqk9lmnIldMAorv9
WI+HPfIlPOP6fA8V8JajyXH3FtL9iNwnVOKy/sieEglgc6aT6M5Qq8IWsN6q5Q03JSZsLgAZyxd7
aVaNJJwNz06dB9M1OlRpFwpRQiKWCwVq3oGVE9Aok0G2yV7sPsGz+GnMMKUUKHHdUzwWPieqNJkg
s/1v+PEoLosZr3H5y8gBDnf4dNzG/Gg2R/7KdydkF4OaBW4jdJJevsmMCLhJIRsRWMqflJiVecyP
i/+8oxjGtVhRH0BSD3tQ4JU79zw5HqxTz+eiSffYG0JU52oDzs5UbxbX6kxOCC3vnYpD7ImDbuhJ
C95nJR0i/+M4A0UMqmrdLuWinopZYc8xbBbJ/WkknsnlyQ1RxJvFW0xBkVw0robL+gcYSXrgWP8j
tihhH7tEggsVjn/LrzfDYK0VJIGD0IrRmLsCFFcUvpQhnc5r942JkxPfxee7ONBlqPMM140aeV1q
4PXD5v2qE2aQ2ahxpLkqahmdzey1/OB5lWvBejzUo9yjMhciSwIrwt8O2WeLRjFnPsvESQSf/OQ+
eITrZWq5aqIZ5mmNVTx4ihWQXtBm0R0l4Q5zXqQQDjqdWUE/I2oL3DlJ0gwBVRDMhoOg5duRmvPi
nehN+gNlpoC3pJ5YEGkntxbePlETAgOgYEy0zxERjToblQjOftLQuaUn0+zSTyFN9qqzBAQv9N+K
gkzlpZCZMldzRX+r7ARmX/IIGXrdoMqyQ92zE6xmpQ+pEBM8yevbYCUUzG3YsRAA+LyMcLNHEpzi
IDFdb6Z9AlpaZBiO3JlxjEoIScXd6VHmu1rUqpcMAYJIw3CHiTwtF1KU8HviH08uKFg6XWJ0Dpij
W61xTr2APL9S6wW1ZiFD7OiftCVGkfUG4mzUnUQEigbXdLAmLPk1oGnhNeqmWFoVZtLEwWhd87pg
QGB2oObkwVdDAqZwKJcqS9EY9AZfz4OV6K2K/4sfpPdvr7kgGj54eMm8nHULF46S4UEHJx8jQFHD
8O2iutU/fZqprMR4rSO028j0xFrJUxdHeqi1FxVRp/7flShU7idp+7qEijpyoA6xt+1yvUCPRBpR
ug7YNoLOgog/8mM+ez1yuwpvJI0wF5lSr1oFniQRrPGwB23ciMjfW8a1Lo0rG+eOxI48koHLHwQv
xNK4OWOi2tyir5KJziKNMgcpJjEJ0w5nAjvS3lRl6IN5y/On8wS+IQP34/l36KnnTQ3GsGZrh0Gk
DZ8h2uzXPsjvyMFCB/Bu3DegJLSLhTd4BN1lx+t84ynb+WR0cIf+lFcGhJpyMeCfPQIhd6IbgG0F
bAisJ/rgAmHiRP59zd1AzaoIc8LI6H2BNPruV0KqLPiMjOPQ+oP45k0cLiY+RpBk53GumyoiHp2x
50QCDaedHoN6/ftzkmt/DyafA+cfpafxxw1XBriJGHG9WaF2wB6iVOPK5TYOgpUAkSNsAbhFN+GG
nb3c+Wvm2MKew3PEsdC9HkixouOgCBLArV1aoJBXjt4V7bc+InYCO6eUXRwdoz6Rqwzcgz4WVTYl
+W9JADKoS7oihbak4fdKuQxqPmtlUFId6yYH/CFXXSUTZVKaNzF/8MIGhExn7g416ApdJB4DqUiy
+j88YpaIF+DXmPpTTYjIA8JVyQtRJUb5io3+wRXik5k1hiE/uZuNfm2fEwFij46J8jnBmDXqAF+X
ufa8IQFu8PEEgCsyW822qQdMxtUUC2+5ECONu8rAof4xNHmIQroAUGeoHnGPeAXAWE7D5fhEKjOz
mXADO4ig+ZeoTr0ZTJyvLYrbvleZRcG94qSeshc7XAHOGIoOs75opo2t1YRCxXOAa6Xcwt1IsljK
MFWR4UXoZx0mW/c+X+TslJH3mCN26TKIgAu/ulDd9avWvdKI4q7q/oYJKDD25CXWBLRwe78r5UrF
99hKVmNbBwsAM1hUCSD4XkYaRKC062Fu6hrYE9zU4kwWVsmYB50pnlKYFy4/VXSj/gXpmRNinKo6
fJjvdGHAKmBAYMygIb3kmXWPuJPKt5IZxGmoGxVzRM34EAyUp/nyFA8PPLeuxpjGgalCd9jVoSTo
caU2hvQRLO3QQ74cl4NwfVFZ5GYaIU/zSvyHiSnrIyBrDAhyd3GZQfCuwOMIJmgxEAl1tHbdZF+d
Y4nwhhRBPfcEw5+SbwelPKGtLcE+00WsOz+f+klQpmLB+8r9PBTKBfix8CnLFkxlRJMfjcSglSH7
GLHBIBeng02crwk3P6oVAQF/dnSRtStiOGwfXy4oibIxZzhH2ehPvuhI2hB76fIhcST+RbymF1EH
kFIwzi99Bs5B3RLWVAceA9uDHxn7+xqTNNLpjvuvaybaGxuHZXg9dalsthtEXf9PJYibydFu41Ou
dUYSTJ9mNeHjhQ7TF6ab9kKFvxLttMwGWXMGOb/A7eZU9qHGjZnXX68Uj/jh7SJSgqlj+l/ntQ7g
zVcf8tk/GPjcEyoN990FQl7VIpfIroJvWJjEyqBh+8aEt1XAkTAz07awK4iqq6AXGASeWxcGTzIz
ljNndK8XUYuTUh61Qt3xyR1tzOaBu3XnS55e9ZbfU7lnnLWMpqIKK8w48UDvNnqbM9kAh0t/Zp2H
nAAJv+zsLjFv/eL4+f+t6c+Z/Bwlxnf3usWVk1S+lJXqe3OkI3WIzKrnkC7UhTzSBlLqKIOuFagW
Fi/T3mYKKi0NKB0PokGVSR04d+eTJY7jxHVsrSa5teLQQvIS7T9hY4TVnVjNYaVi2grnKG5yHLUk
XKRxYM3+wVVnoo6F8LAKzL3caPy6/eifkuwEEO++mLW1vAvib2YzKfoemxgRae1r6Rl1n4O03o6Q
g13WKYLSzsk9FvbUsZk95iHR8WoYbVB5pDikUUXe9vASE2ndmEDK9kjLe7L9Ybr72LHSOtExifWW
v/cmMLzfhMFgaCKngHW7En5AFAvFj6KzpGkoVBlp1Jbd2v1/Ihf2sVhh+i+3Ba8liL6ithuoTxNr
NGrqk0RAFdv6a0viTWMLK4kPQY/i5u0UHqgpPC7yylOOW7pMhYU9zR83NAB1UoQ0vjeNBKQhjzvB
LC8yJanuXP55N5VIFTmh0DizjdcQoN+LfsaP85Cvmhf9majg6G/tB6eXBn64oqlUtEVAAHd8Zu+r
WnlRpUIYt9ZJOUHVzVtP5XjcQQXldIF7WgTwp69sFFT5XdMgDu2D9l7xqCz5bdo1rffL8BjmZ/nL
8x4M7mRwBfZyEW+KMM1XHhu1tPho/N81160+qcgDjpRvnp6D2OTi+RWXNJ8wSbwOQYGSM1molu0L
J7RH9zN+WwKQCxflUXEPq0OSNCgRfCXPxEIYgJk9cnaoKUwAHfIAWdWndgz2l4swD00p47WRk62M
sq+1zfnRFtHAioJpM5wXaHJNb53IbgxEuPasw18/DfdgW+395G14Nn2TZ128mf0NPLIBXO4S2f5g
ymdALM+p/kOkaCdHDq7UOOLaxG49AHFPT7VZcHjmXLgflS1mobD1wepkbtG0xtTuKdyuPYEuuLxl
/iTx1vQRYVcPzqDComAm3VCEobepyaZ0a0GiIEEyx5cZP8f3N6KGPAq9cF6sI+nj0pWriRE8VPRX
8a1rc9SZcVR7AZJ8xJjddAukXn6pSmvULJl+TnETo92s/EBCn01oXImaa3exl88gFRa2IYuhYTN/
TsIwnZmHAe4p0H0WMYI7qoaIsJ5vJhYWIILptb3LGQ3RaDZtvTvWvvEumYPFe9x7KUCLW0QRsNbk
ga8ocTr1YH/lE797uVMvYkmKEwE4+2ZksRjv6l2lLGgC7OulTtC+4Qhvt/ZmQm1sKZJCmAqzbo+r
e2hjEKkp3Bt3dSRuPtfvt6OxCaXU2VmozwkddCA+yU9xa3Q9wqkDVXV9AVM47PaECy7Sm8nwu8bG
hEbAzwfcZsR/vIFIbvm4UiGSLkibp8KSCQkUjY9XjkyAb//BB2KdddyYTeYm9aOD5a0MfVgwdnOX
yMZXessz0XdquR6F2VStrskxvzm7OuuHWXyi5UwhiAipfIeVfrf0veh2gw45G8XWMn7GN4YduFZF
EMZW347viJDzKM6Gwu82Okcq1JGdaff94eSh/3rkGKYTU6HF3zkeuuzBjRpG0BZQP88ygrirVSzu
kXQyEMDrxI98Dq95ovWkygpUVuBMA6qLpNsSx/msoGrE7phIzlZz0xFa5g9hk9MupR87V99MfQ21
u4ejZw7VUms1rupWYENIxxSNpscD6MyF8ncXTieq/3XaI8LUCdc+4l7bzK+QQ9TbsPbPCSWNpyvh
IYnadsfzZidHQMzD7fCodLuwbtCW0EgHteOXgTyt9UWUhb+HwZp9eAj6obLJn4H/dwjPemA++DGz
jX2RAeEd99SiBUzK6OIzo078i7/49RBMPuYZVkVmJGSML9OfYyTcJ8d+H3irUdrVjrG7I/pItx8s
eL6FWPr8RRygkfRVfOD8FqjoXipJR3U4D3ezolFSPRXwkJi9hVhjbg5jpGmWOhqlM3jIbi2iYcSd
AhP2Mkv0Za905HNu39vZ2++qgPxGhnewCb3ZisACTEYRI3k0opAgUlpl1Uqp6KBRuUtfRq7Q+4F5
8BxngF+QhnxLbqfLsiKl8ZQ2Xuag9IIArHORtghOIARH1FJd4HsniK4FArqoC1z0M3Ye+EdtPFHE
Va62D8bVGnbERlWzoQrtwD4ZGUbk6iSdRpDM6OMAcHg3cHlewICH/ZbJbR7W9IQEmwRsMI0c9UaH
AM4H+DrrF3iqsesRPJosLgzTsi7o02lf50WTKx+dcdRLnAgjGmICTc74jiUVZ4515I1bkuiKKDtD
ypEhMpRtyJxdBHjdXZBCk4P0a+FFdgKf4E5nBH5DU4JoBu0Hp6uSJckraJJo+GD3bKvdkUr5bGbB
P1hyxPtQDb3vY/l2BkRbRgGoEtEEpX0QXR9cO24H8xgC2e5AclmbEeT1zyoxtn2rQ77IW5iun/gf
HcDQTAwPi136B1G2547Dy66x5y6K0Vhiu9wb4VFptmBk0k8NOYVdO5Iv6uwRMu7b+Ot0BcjVfHn0
Mg5bFJJCzr2SiqhqClGYSYPyzJv3D03qH6QfhPUnadw/DbwXSqYXZucPCIhYYlgnTzZkUV4hxgDg
auuEpZskq/++p3tWvmvSIXiXt+HpNdt0x5Pr22OWJPWMnxM1Dah3spdFcJIdoE4f1aQnmZYavx3+
7jkrU8l3qB7z27NlGz+wricTjil+K+7BJMnkPKo2AgWqGBsu4Q9/AzXBA98YkodAZFrDVHC3rey9
yjGjBGOPN6GxZqxjuAOvWbtucWL/V+UgHxrHG6mBhwWpPJSzC2i4lUWADSW0kkTJ6dTZV4PaOhoR
GqT3xv/dmhwd3T8GOBBDdD2gr/IodJHwTdZ0cmtVVIUMJRwvFEMDU4GtHSwUpQmBTpmF2vtzwpKd
gBdKBPB4KAWeVdckfJh4x1YBrh2LY/KvB8jo/UtmET+bKdea57F2ffUmphzKlH0yq7zuCUFq9eFY
yMohkEnGK3WkWo8T9BchYnoKFCGENf2gaPKRFuE38VyjYw7hHsTDmw9NNuwkpklhQNCoxZxR9PHc
GRHTymM0nACuCAJPNmT2PVqE9F1p1F8n9fsxq+MbwAR8AZglvv/30f76cIn/YsrhpOT3X7cPyQe0
sMGXjymKMmNwm4xlHSx8gndhlVYGzhhvv3TcBDxouhDst7ajZG0P4u+gUXkULWJ6GsMpNQi7BY7Z
12kN4OnScbPO21NVIGRiyR+Dscfbxq8jbD1NFOy1j4YUPi5HIGKOQ/ZfYbHAj4sZgry8hp/jp5w4
TZ489brfkvLa7Dii9puWGww3IAl6KjH+q1/4mo7Hyb7EzloLwRxfmrTQHK/EKabIg4TFLayIeReR
W5LX9OBw4K0gl04EogbEUoZCgIhc+EIZEmQuFFVG4+oJyXsnQkLCt9oB4B6LluOBssOdFP7MsWLQ
2gg2lwgQzIGw96eQabrvsCsyiGdNyN66bvqK/m6EYqMf+hMY8QX2p7JKNw/C+aJnYZFVeNIx0Phq
FM8rky0kFH6Xp7W0OPrgvpM1Id1GcNMJjoQEdzGjnzM9PQUtAuWgEP6+vobaEHKrlI6MznBE17Hj
yOa+X1SnhjS/xUpyM76cpVu6EqKiI07u+YzULG+n/9c0COj/XjWi9p9VFu49MHDPHcWJbKoRDPlZ
k9WZJEGezFUx/6sfSok5sdLkkUed5bYKFVfTildLXTIA5fglhyZAvtigAq7WQxVXg4eO27SDo8nn
I80/h4pOwc5vRvs1xXllP39Rn61Y6IJf7BRNnyDBN8YIU8Nx5KK1eYPVXEvwQuvS7lBkSnBmFZUT
bLsVWK3g2cIrb9SbqAuCWCJGYScLEVJLZEtnNLkTi8yOx49p2FdmHn25BmISDYVW2e1gYLGoF9T5
rf7o/cPgKA/D/2QxhpMf4qwng4+QOh67WrQEe9LPwfxQUkK6F7QxhcOpjnFPM8FCVmADOp3v9/Bj
Mx80KtS3lKGZffWGbZHPtdcD6swCol8D6JOhyNCA1Fml1bo//+ipQ+irOvUEzNBGquGqdYCrqgC9
Hg7atp/YZdHZFiaqQDQvT42XvXj1nj0wWJE+rR3E+kLwEcJRcFgJhuaSKbIdslxxMNRdNEglqs5b
YqEDRDNdz/JNmJQNHVLTJZsbKcCdBmcs0AJr3PonWuc2nqklY8cW7cT61LTENQvz7W2d6GkQCdYv
WIcpucPBGytMtpZ4TYHz+KpLSZ0t2v2ZJyqnEU8vxngQ5/zbQBIIuaKXUbW68ZvdcPX4mKFJssan
pRrKLFb/TTgz7IgjDmBvM45Nth+e93pMJdaob1HEWYkaxLLHaAAbrs3cSS4fdsB39N6mMv1CdSQe
RqHXXGVPiJHDZLxleYeCRzj54Sk54iXMmUM2l0iOnrbK5PBaUgfJsZXIbdNNBSPekR+x4oX61l3C
KOWwP0h2vnJWVNQQFUuaVORtkLhRtSwA8FwaG3DBjEML56dppg0W/KnVTGj8FhZ86Kv/ZCZH1aAq
Lr01OBFxE0NnsINMQT3l9uMmHBaeW0AhQ6o/+H6YZsLTMOIzzX7Gjl7KP/HsjcbL59PDzqOXajq5
jQlcoMvQe1EgXLUgcDdXQ6HDdWlpUl5GQwpDXwzdUQ2TK9AY2PlnDyLHdWI1JpZdFP/qLv+jsz1X
orIMYs5ZEwZlCrbdPvNBmBLnIluLcLvRiC1juYbixXHYtxr0K5tNufjfXaeb2SkfCepndGKs2DqY
USgIyGSW/sukKsE38q9ZpT0aTl3TJmmoNO10OvIOk5y1RY+c8dcIQBB9TPdAk4CPEOwdHkYiZm6k
78NnhElpBmA20rB+fKjDT3tPqk54pWDN+VrcdZP8fco7k5TVdjtdxQNmzxTNSogzL297fjC0NIpZ
nn1falFW2wDBI/sDQw7rcwqFIwaqHwZ/kt3Rau6zMkGbulUdgt/GLGq2nd0OGll4H1NXxPVP0/Tf
Hsk/zJZJ3vVjlC7pEiw8HoSO/eL6Wr7jN+w/rh6R6tkCDO7cSyd60fHnODkv0wZwFBcfE2L1MVDg
wCx2otGkTYlGLC4sMrHcnPcPcU+5rurAp0eB4uy0b73bluTyjQIl5BRm8/IG5lAb9KyY7lioRmna
APfGyufbrJu4TejTIc9u+exYnbjHOZUN22quVdb0GXSipqb8uhCCan+DFusunrBxVr0Lb9YivlL9
A5CLYREGkTA2z5QQUwrBOuvdR5Ea3J8RXP32YZMOvMeKmgfRBSfsMMotykddrxgpkBTeJQJSSI2J
3Hdn0Werg3tthKUlVWoiyH6umEdsbq8jI8oz3Ita3JWhtbBUQA6UC2gvH+yl43JRFz805OaupBh6
6WojWJHcYR+Vmii/QsgUoKVVWkAdGCJQssoBrRDdx8MyFn/A6KucDZJcNrE/Cehvd97o4fa5ryvr
k41DOh5TnvhlA2729dihiq9wefNC59qB54WV4zP5dsFbHcoUNrbYplPBMo3hJPcE8bS/4TUvQAJl
gdaUVzWSFiNhVpC5rQDJX015kwhPpOuQjtfwUVYmw70cNA5GJomF9AyY+EsA/pGKnXfyvrYFYpEH
3N0Go24uPTrmnZgjsXZRhkH8bTd6tfLqwaiqL39LloL5RhL2S0m5KTfqS/gzxhOUzvd2SdQxXBN1
Cm36xLks7Dd0urdiNEOdye9eNLV4BHaf1LGanD4MopoV03nwsaVaA2diWNS3WtgTU+QHfSWLQ45i
046kofMYjdKprXVuLZnIjuzvccQkzExGfVU3vMFYmbP2AHoFk56J0z+3/WSQ/MqrMvtVB91u+tXU
GZvXBVOezPyk+Glm8SFe9dzYFWT/uSsIkhNcyXUn2TUkkylkPTFxEjtfTmDDOnVpT63KOGE7TX10
SzLWqjyj8m3QPLJmyQHcMVY924DJ4w9BRevH2BMbwG4Wevd/OxnS8EdKW+qA6ok9TFY4CVlYbVzt
hrM6e2OgfrARkT17MGavxVcfePYVp71XV7pV2OcZfvhSoabBQhpHO7l9x3tOzYh0LOVzhsv3C+Vr
RfmOoBuCptrt6U54LCiziWd4kV4oIDXGbtPvTZ/Nbb8LGQAIuvlCn5IUzUjeOh3nTMpz6eMxwovO
TlsFOqqyWxDn6hNNDu9JQIe/OhhKTFk/1Nd83YU+fC82+bnaJBqvGBYROjCDdQ38AadVlThLjtnC
xRV1rqn2coBi2ES+8Cs8SRkJvxdDdMCEOMufOcEk+sLxB9KU8+YX436y7mnIg47G1JeQPqOWuJ2/
kEdQUw2ji7VpoDLj/2PujgcWgn9zfcP7VOUtsbBunXOErsFGujPxqmaBslCXsZ+MZ/O3j1vKBWYI
VRe8AvedV8wbLbb/YjyX24QagH8SnaUa5Va74fKNi508JxmffGiCku/fRm7saeen/B1C0nufDUP8
LilMV0mJyi7T8HBIoE9HBEGFXANWB8gjdEDxIlpTOjC0LSKaZ77CAQlvoN8pLMimrYY0suybV3Pg
fEQMkCS4opNDgOeJPBghPMVP0t9GhYeN9WV8ZCjre+7TXcpN5aOObcOrK0Lzb/5MpH4e/SK76Ggy
cRDh+WXV9HcpxzL3Om3k022SXSyjwMO+nbctYtNRtPomHcnBfgqFDa52gqWuD02S8z4ogW70RslD
S4umRr1yF0QewFdOl9D9ye2fCS/ttlgMlI9hbwyDH5wa6//sDhP/hZGqAEEo8xEMKmdxHuCE7a2S
w4g+pwd8VLz8CfOgAtSsGMPU7Ou+WwYCjGY72I6EgJ+DrkAK+n7zrBNhNvPL+i3ZiqYT6L77DxYK
ULFzgG/OtQVwwlDnTPP072WX6n7HbLAI0iiN0VgcA69E/aAVmKCwyLP3xaolLRS7zlpT8z7TdyvE
F8bkNdJ3+coDCHh5NTO2r3afHK+XsW8hxISqcIBcvZYgNae9RLEAtprE5rpycc0catZDpLYfTDj+
KTZJGEY69qGE2lYhin/JgYYX3vm9OcQsZFaEcWcvDJBo2U75DISs/iBGUj0jX145iGoJhdf1YHIo
eih0PsXxdcT+E3UKDwfyr95mzEdxoEki01MSslYktZdm4SaUzjpewlNd4kMwKgfLv17yox1YwRPz
rW3NhWnQSZO6n0BhERo+yN76hdK5uBJnk1wsvw5xnucQ6efPykhLlqBoxgcB6Y3VUbrCLvJDnG83
eXNz+1c8UxVO+r35xrV6rm5quzBJ/C+G+8Lizjn8AVX8yDzTM5Npuy4P38eqqUyE0KFfWgkbqtiE
xHBZjhF1L9s0B4H/zbYPFOKoxyvKXsXbz5IrdmYixMbjHMImbwfV8QwaUYWff7XJ2jpTv9gX0kSV
fQW0usjTZFL5Ik49C2NNVgEptP4BzC/+Ke+vzonANGzr7aTLtndyPVH0NXrWxJlZQ5ZLaTPOP/Ct
Z12R5cIa5jesZ5V47qX4pXsKOL9Q71jHYPBpOO3KV4FkkvwsVLkovCyDYEMYAN70/cwkrFu5GXq/
WPCXSXF6ujnFNHy9T0UfICHrRWrq98RHe/X+tofM2H1hJu99yxiAuw4umOI/WbfIU4fDQlPqMwkR
Hs3rzDEgV0FgWaYa50wNAodT6RZ7NDPSTMwqJmXyz7Dz5pnomB7lZMULOFzVobJKPUqtYFvbTSoT
GEaVAv8UY6v7g+JzA+dcLIJUokT2L6HNK4aCxwhB478TSmFRSaehBznSjz07QNTLUKKn1ajhgYEq
djeAPht2fpnUsBwhvcwL09ldsehQuHrUQ8HTHTTKGDQsVc7XEn9b/b6sZXMnYnjmmHusUHMbOawh
zkh5JgKGFqZ/8EqtFwM248pqBsjB4KIVn+RkqrXpFkJzZFnVrpax2blGBzxvmumTNumWiHVMG0hI
DpOJaDpGanExx5yKMvFdR4q+9P/mQq/ekl9BLnk/5scgvNqxSZwxv+1LRZoMymcfpWdX4h0LQAsU
lH8fV/LoHIGepfyMotWlKm0RTqAAX61Wwk3+oOHJlaRbt/HQgykTe01FeI7cpN+r+vhaEK4WYlo6
779mC3St4KMpqcXgc+vReefB0tC/JHIz/u1rQNZZXSvsCr9ZUFwqGlOeCKvsbq0DqDV5jnKmHGIP
UCczvl8Rp7TjohNJTvgcwzi43WMaWwo07vDhyc1VvSEju3InsU6FSZEAeOSXgYK2csWaig90g0cw
+h9IUANvlHdlFgC+3sq9etWC8aQ2X5y5+HIfDykTINAoM1CWRu0SJ/z2gylAAXEWDoP3HTTLXKrH
YZIZk4K+eQWY+5dlaOIOqHFMlMHGLPxmW+alP22lPUI7asagmwpZxQ8sSUMctTZjGKCW+sHoIO+Q
DofflhK+hRrOCSkRZgPMB5aBMDDs3cDsPsfPIx5IrKvRjt9BDqwDJEkE8B6NHmD/HT+1uJafnMir
c3pDOvnZO4bAGDV9bIujU9BvEj9C4sTitVIdS5XRtqGx75ssNFkcKhr3QB5gvUDOA3nmjhlgkujp
AXi0BzUqseRHZNyuxIlBcfEQQi5+OhUQOPvesaKAKtrgt3qcNj/FjKW/QTTw4EdRrYv3bcryYCvq
R0f/Q5Or84o/WKNLx47zpH33nxmw4VzliHDRZK4bIsK0YADLlkCZgCxQiagnNIaKWxblavg+er77
mdL5CnSWsXSqEvtoGJ+A7Tvw7BVTKkDKvOqRrFdeBmCZ992CO13Qcd9Q95wzCChFZL5h9gWSPLXn
hEUgwlgGpTSCKvH4Uc2WEu3sR/WM6KkYg2DvyMXObEjvklHpxU4D/Q5QkK5mg+NmMuW/HtKO4Eve
taSn42XE2wC9xeenEwJetWEn+gaIkagynulSfRVrqfeG8Dl1HBEG4VpHio2vo3aIhYv7IOcPtRdd
qmxRzSOVDIXLL/Z4zLqwqPKLy6YzvvuMd/ab/gJ5NPKfVYWUpD5jKb6f7pJEwhr4xeXMdPJXKTjf
8D0UeuOmhslhrlKbRuzMtiq2BadmM6alqKBVvb3w9sUq2noC0uT5GZ3A4eNRGOPQCQ8veZtbWUbi
EtozjOONymfsebzQ3znZ42XZ5yoI5dVMoaQdYP3IJA79TB8/orVdZOJn2PtjTiKO+XU7XqbWfKz+
JQAr1oV31KhI0hPnTqadOqRwcIOsk7S78gXpzIPXcSi12XqW1DbgRcspQkJvWg5hHRDoUlVxvZVp
k+49fL7yctFLsEaNhuZmkSwt62pEPDSpSMx40bPMSBxulSf5gjyAm9qlz2I3c73E9Hw9S5OxGZJN
IBmkURwqw1vqUwBnlZ3MI0yzB2R30xvhklrFBteH4t5epPevhqO56Um1MwVYny3/w/PNTKvnFgGH
5FLd18OCmLBL7KIA6kEnTl97BWAddCTvwphCoi634F+DE7QRby2YPGVIezJUZZX2Wd+KMNREKF2G
xqh6doxEitsnUyGYCY+Ef3DlPGbmRt1c1vXaoR5wimev7iSWn1fx+vtsHrz5QXMbg/pGMoZ2ljDF
UVd0HslV/Sz1Fc5ZDDcoQQThZt/IAcXa5T3I/Gr9PZFq7sZH7I3+wr/mJTc+A+xHEpSzOhVpo57r
1z6RBQIyn8F/qxZFMzwnivfnorzQ7THXuv+HX5wvh1OWTYpTgZM73xQwHVPUqT0T66fTCbqicPeZ
wG+fcQ0wulXNQgLZpRfxzJXXBOV5rPtVINpVLkLrejxfcBgKzzEIZVxDQKcHdiI02EjZ8OF9udxu
p0JdiwPdqKo3IwGZS2c1VUisPCDtymIvRueYPtf5dnfBsB8Znn+3qLBck5jsJm/EBh8vqbRawGqD
hRZZpaW0iRSX1eqKWCYEJ7XpxyJeq9/11Op5W9K/WZtulJnl8YnyFNs9AM0GEyWe9qahpKXc0vN2
5bSEf0heF9APQV2cIB07HsTX2pD9SisqwagOaH0KrdD/IPU7eKbU4em9M1K8MLHZyopRIokdqLhI
59e84cPbS+kAHWHMAFYzdd0QHCs4TbpGZFxppI/AeSk1w5Swj8TCkFREzkeqgOORtl4Pi/b/M6Br
+XlynaknIqDFh6a19bdH0YtmjczHnXj6w2J5TWndJ5IflzTKOxnl6ybXt/jz9JbUQJud0q188YMs
fMvvLnO22x8LTjhR6krmLYZzA0YmDlbGyi6RqnCs8Y8ko1Hmog7baJPGgMYbxjxjRe1GVGxsXk4u
KTecEzueSQLa+QR9U8Rjv85nZyHFRBjhOfMyLkSEcdeQAFWauNwCjB7alN+URIOMKwTPV0Cim5BA
zHUJki2isPzFpZEiSa36S7xbx/FOAZNrl7etrLu/0uOV+R7PSrNeXmkhrBXIHtsbBuxsGLfHznxz
r/w4SqlEtZ7kZyJVms1ozr/Tgm6UPzWxrnrHhuYmHcxjemvo/+Mh9Vk6x8ncFfifoxoedS7/wTa3
ayNIUh+1MgliG0GRDzSl4GSTiOBmQQ7I0Mb4vu4d6v3ISl+8wVEPIwZ+Zo9TnXTqdyZiuZtzKCqS
1YmtkNAINjo7JBxfBuuOu/2Dx0X56A+MpIPCSUbneLB3UFZiJT1T+xHErb+ESXClDKpd14vby9kj
Hn2sG4dJPPw6J9DzwX/aslD+PStN7e8CnioKkj9KNdo4ON5FAvIbBpkXoVUOqProNw241YPXviup
aNCvNbbjJvZfSG6nPHpf13eBCbrBaXO6zBbby35IRqnb7oOcqVnToViLTZTmVvIe4FJ/VEqcBvtK
fqIVUhO+1A1wjuJQBa91e6lI1blEnbSRQ8ln/5FwElVdtL96aMEg+o6uBbfDMQNQE5i86dlVF4xB
tw8OJ+dbPpiM26Oo+uHnAaUukdL0+qSAWeAQo5xOIg+LsvS5xugus4tG5YCCDAFHDo3514g6OqDW
J7QwnOmhY07FkEIpWbCLScsQDnfncrNFrIXsQrts0dAEnQ+Ns/tdlwo2Uie3EqRRVX6gZLsl1EqI
8ImfXAa+OThdU1x/fGs5h4oZ5WjQDOY/D94/Bc7aKIg2vkPrZjHkqKoVKdyDzzMHj+sgdSUeZWM8
gBw3im9Ot5Z/TPSQcSHEX5x6zOuOurlrjoyBHdhU76LJ2eyR1wvEB015qDJOdajh1PWlTzS8ZvrN
tgaRfZFHZAIqlB7AzQC2b5uP/6lOGX+9z/iS0qm8sg7F/RZz0LcLP6Kyw7F0n66JTFz+NQrDUSgp
cIgPqrhRmQ7XdzNuivyaEBFH2sijGcIdLnrqYUhZNiD2Vh/gP1NS7EyzQR9QUzD/NYSNn5N77l7n
SsCXFLOVeyxTr1MU4gPGLeYdIOd0/i8lyS38RbOFrV0lHAFDhQgZ3g/yCLKoi+z9eLoCq3N2R0vQ
uGhMI7Mz8ov2ORA6AwGAB/b7b4keP0Phs/x7ojo22C8YD60pQGQw8ki/qSJJgH+7Oqi2UrKCjF2n
VPhlSMuvmzvQ1jqOniNSbSYu33+kFqhjTdXc3sDhMduTfEH8dzL9p1WcSqusb1BsHSj248pxdPmf
dGOcIKUPL7UxS/6G9j8Ly2e7sRn7GX0Xa5VbptfryOT8fqlpBzlM9YIB83rTKXp0ln5KjloeURr3
IVmRYFXSaS5WwWAXQfviVxiaMdFfG+0mipEVFeCYonna0xCKqm37XdDvPb4UZHx4+9tpvYlLkEP+
+46uxbFVLIF9gphScQWDgwGunnBCqVXI4UJFbYxhH/LwtjQBTMz4Coi8o6CJCoHVnsHrtmPW9rv9
kA+dC6qg6xRjclG84ly1QqTMzStzTdAQThkJF1H9YMIKADZvN4rsCyC7eLGRwr9cHMi3iB1gCFNX
97oQiJF/XwynJwI3J9wBVrrpUY8frAsUA0wMERv/KyPD+zoPUf7c1ayDQtdo7N8DSJj7pTdDDZtE
qFeneUO5/cZmQhgJxBQvq6H0TPe7mJd3eSxkLGnDmToCAsLLwscigSwcBPsazYPIWktDv3THBr2X
SPTAStCMiZ2XMjqoXgIIaTzw+xHy8tqTSOLsvW/ksCyreSBGITj+p8XnL0bAtIbVYUNC3tDaz+gK
658l6hnsIFLhk2isHt/115QBdN3WE56DP7WvwHsEEwjiLMshdbk0O7enL3LZkmuZASJo2kzAl8BW
3C/h86vm865H+cOkog41qf4c7WBgslyS0+KBCBJloKuKCTHGUJAqV5knkLmYjnx9IG4ztTVO2nYq
5ALm3J8Eu+zVtgY07LkFR+/7/lx6yOhjvSkdR17QZQ==

`protect end_protected

