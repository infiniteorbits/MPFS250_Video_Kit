/*************************************************************************************************************************************
--
-- File Name    : h264_I_Encoder.v 
-- Description  : The IP compresses the video as per H.264 standard by using only I frames. 
				  The IP expects the input in YUV422 format and implements compression in YUV420 format.

-- COPYRIGHT 2021 BY MICROSEMI 
-- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS 
-- FROM MICROSEMI CORP.  IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM 
-- MICROSEMI FOR USE OF THIS FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND 
-- NO BACK-UP OF THE FILE SHOULD BE MADE. 
--
--*************************************************************************************************************************************/
`timescale 1ns/1ps
module H264_Iframe_Encoder#(
   parameter G_DW 	  = 8,
   parameter G_C_TYPE = 1,  // 0 - 400, 1 - 420
   parameter G_16x16_INTRA_PRED = 1
   )
 (
   input              PIX_CLK,
   input              RESET_N,
   input  [15:0]      VRES_I,
   input  [15:0]      HRES_I,
   input  [5:0]       QP_I,
   input              FRAME_START_I,     // must be before frame start
   input              FRAME_END_I,       //must come after all bytes from frame
   input              DATA_VALID_I,
   input  [G_DW-1:0]  DATA_Y_I,
   input  [G_DW-1:0]  DATA_C_I,
   output             DATA_VALID_O,
   output [15:0]      DATA_O
 );

`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="author-a", author_info="author-a-details"
`pragma protect encrypt_agent="encryptP1735.pl", encrypt_agent_info="Synplify encryption scripts"

`pragma protect key_keyowner="Synplicity", key_keyname="SYNP05_001", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_block
d5m8C70CaEK+QUi5epv8NDm37mCI9r7ZKiUl74wRL1JtxUlqeBFabwUl01+1dq9uAadSuxr/UfLy
rJkZQ4vMKsDFwiOAmzz9FYX9TErX7mbO7WlBkwxv56V+SNaglFDdc5kCsFZoucQ2EwKm2bwfKY/i
lAC1YsyfLYJAu7ZrRYz/NA0NL2yBr1udfED95S5ObH0K/6xsEcdO+zh4TKBjd5HvDPMApb+09QId
bd3doMcR/wHoa9vGvRLDACtE8gymHLGxg7uN9bFPZ7hNT/fH0OKRrXqucJqxbm0Bic5GhUFO7jeG
90vkhCUxpyQd6wX1m+jlQrrpGPkk8LmkzAUxfg==

`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_block
joRxwvbrKI6AeHEAv5+LXWj3rted6ecnGhKImDQudP68dJCPNtFCNq+Hy1B+9hkZTdOQqNe1AOIX
vEeb0YktV6Mm6ToO/1RhNohz1Dq570uFkof70xblnTOY1AJseaos3anGmSpWNkO3icMAFp7dx3YI
Te60wDYnLfDmSfVL8+c=

`pragma protect key_keyowner="Microsemi Corporation", key_keyname="MSC-IP-KEY-RSA", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=960)
`pragma protect key_block
T6gQcvYiCYEso8WrnxC/em9fGkpS/AkjZ7IagvzxP/mGPwWaLizFSb6Utqcsh4xeSbGqyBbe3ZCY
OI4ZWklbZruYBqwLbzySIP8lf0xRtw80c+cj3Oog/DFt34ZB+Ju4evNya2B0Ih/Mf3+EBzzJquEb
j5wbmhhgvkeKwjyGxhCSwRrQ1nQvvAxzBA/Tq5ulqYJh09dso0YXq1Jj+ydfupnLWraLEEJYqyMt
BHi604LIX1MOAvEasjWGBX9xv0jN6YgChUqsC2WIecMGh25f7Rn0Gu05K54Svd9HETI0tiTFC0fS
grf+Y4ke57ycavcqV6e9BAOP7aMDb+RMHonZj7I9BRx/qq9SqBz4SIPnxYBzgWH7/H1slTof0t16
Fq6zCWUl9kOwD6vc4dKr56AdofIQBJBlJgkqOSMeHQltVT/Nz9nURaw2FScfGIS7DTNKwWd77Fze
k7JiQd3naDmHF3gjTuC2JoV0KQNNjZyME+Ku0/fOL7cdYTAUbiT6OoExeSLaL/llGL34vBWl7K1l
2N+V249XtpTZ01Ta0fxR2RUmRkSfYPdO4YL3p6M6LEKqsNFY+Sipaj6w2wi4s/9YZOnkN+DwEFg5
yA++PWnWT0vrFEQstVzzTjf+42YTHkxNAEkNbx7geKf8jQIFse08YFSCp9kwM/b1qKEMqD29rxhJ
rI8N61G+OB3mPsedvj2NgqQpjO1VIGFqI1m6siRmz6G4opv/sW/fXWCMXA7ftmmo4FB/b9zQse/d
CcAJf0Hrsh8Rf+SPdiidVeVZOgzY9lklLzhNLj30TYFXzo3kAv+AnYusWQ+cBT++gp7M3s3nTt36
rz+dFPabEVtvc+MthF+fIND+AT8LXGJ/dAh8HYnGYQliS1zo+A3RUc6y1/o2qWkxRBJocPZypBdU
1zC+Z9Em+sp/FwWs6SpoFNUz/vVcoxxjpHpl/3x09KsW3AtEuUWMle35KoWt+H4yKKuZL7EHJeSo
PPReL+DnmoKZihCuEnJo7cGqZIGNKcld/mrj/PovN74wW/wzN1VFir+MVKpSgqtw9gViU4Jdrh0t
I72XqRbMqmeXLQOTC61Jrnyd1VRV40uk5WeWOiefDcbzydKIMueUEmamRSPhf5H3mWI8oh+Zwy4p
op6HXVa5FZTXUFoz8SNJzqp6txu3QndGMQMI1hEKSrT4EQ3ZGS1sP2twldCP6WHsacASirjv1/wG
26Y/DmLoV9NeDJavnZvT4X4dg6WXM+xqNh5Rvwbe4tVZkZngZtgWZxNwgymeujqb

`pragma protect data_keyowner="ip-vendor-a", data_keyname="fpga-ip", data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=598080)
`pragma protect data_block
UdC+s2QI0Y2BGjnW3YHVu/7ZHDWVvFCdm0akpAMn0OjjBBpNXJL764RLatuEG99ERaLXrG5xMdXO
378fBvSZohyyQz3yKUzhfLIGasW6N4NyCcJSZva61OLK5KjxH0qAOTBulujJddtXRF9f0QSqLMQM
R3HSBAF8VSQAX2n+VO+blyUBhJNfnhoD41pdE7gY1cZZnUYGCB92FCZ+iJGKnNMpPRMphg0zexPe
jcEQaKhhvDj60ECOTnWfqSfDgmEkOBJL33+W8fKblePFDpWOVZamM+y71WVWunv9qis4wQCtgvEU
u2P+89/6F7SqHYYS0yjBvme1AMxVPzjo+Di02V71RSg6iA59XVM+fH2Rwi4PgRbWvt/iVfPTYeXv
RQwpxbjjIhyEAliva+/RDYDsskTguvIGJATmSOhjSxMDYwolFUtxZP8iSPhYvvaPj8QYnaOdo6dM
c7R31jpKUhKr05ln0G7IC5MvRinh/LRDRM+yjV519r+D/m/XisiV0IFAVbMzeKZr61cfrXsDevwP
pDezsr5NJUQVS9Txk/1R7ei08+JXna97XL48bZNed8hzRUgZ+OwInUo4wDxvvfRACgsRmZvp48an
vK3JutyDlAWPhY6T957s3m0Knqytg7MxnMFxs4DAg/9fcjECHqzP08luoX4Ih0bTbyenwEdbnnUn
KXT1ZwPllYNDjkKgfMA1o9KvKeQGru3osubW7FFasMLbVvNankTGa8rBFhd4T7nxlilDHrsuO/xS
8Q6QbQ9peY7OI60es4Yqo3HouBitXf0Jf3PmrhdtNZKtyAs9PTvzDb01y022ZY/l7/cM5TQFh+Nj
lxZefKZq38+LeHMTmOKQgMGLdfSicoUKJxfJXU8aIYm1QLAX1W77nm+pMkm0VCkLrsbP7nSfjiWB
hUPSR8NH8xnBXBd0desPFW/WIrQZ7LwQjbs/NJJGrBuPDv4A0Yoex0/Bb0yycZPayF/Echp/d3WH
xSd72UYdF87dUVwJvt/nI+aIjye5sVuLqT5ANbipgCQdrB21L7cl2JwVmcJ60p0KCTMbDdiqgNcx
LcF14uyUcCOA9BRqU8TFTORDbMIDCk7YNS/ZQBP9CKtqvfd4gbachm1r/5P8ngouFiyedAb2Tzwo
VNhdjrMpQYgWR452vS0crNBLK1rUKUJo17FhUKIHX/kSAjfGePM7Cq8/Ok24oquK92JTddiLP9e9
ChInL4FqlOXSTXcrE9y3XqTjaogu0TlnpW0jId7m/JtslFYlBKjSrnAio0jFDToIasA1SbVXbGiK
1UXdtXlmyJk+Ut31XgFvp1LY2VlCNR1RX1SQJs/Ablsj89siJ+tNbRLFNH/3EFs80EGN98WfAbND
b25xln4BNY6TNiYH+cdSKNrYTMBMN9gCKxIXsYccVKngC2GbGsRZSFUhGv8PyVv/Qvvv6ghIs1NF
HjwoWa6QDOsXJO/EHmKs2yNAQ1+1UE3B8Hf1WJhmjccUeGlB7WPtgUhz0UgN5HsQTpBeorZFtuhc
WJGaZGGe9qnWhtxkTfZ++Hz7U+jqPwvfkmdI42JLYGqrfUjlB+xDIK1/1q7Xzu5HyldZ249dFBCO
/khX9fWc8jM/1wzlySI3jRxc2ssP7CU7oR8IhxxHqGjfBKtzQ73771gAGqznYiiCfZIkEsTKVhsR
ukNuuC87aBoi0mCCqT+D8jnaYKnHex62iPEDzR1f2y2Eo8RsvaOp8JV3kIDGCPOY8Ikjg97qB72q
Wm2hEPiHZPedKeSeOrt53fPlH1rOvrFC02NNjbjyIeuti/g7RY7VTvsWAL8EtIYVG3g9uqMUdRR+
SI9QlBQSB9zGj3Jnr8tyQyLftxRw0p7HRbzcCYthS07qlJZ7hVa+kcJWuc8gVCnGFtjO52GhW2H2
miejcXxvQKdgoMS1H/HlQ9rGkuHSsV0XseItaYsllBOKn2445aYmCWolxmBD1djix3CkYIr5x/rE
MTOB2mXrs4fLV8Oe/FU5pxkqoWXk4qy2RNWCIQCBrYWeO4BKoUFoCdO7AqirIhd1mcW4x4HjZOiT
dqf3tXDVHh1wMttU099X/2rBPaemhEtFVkoGWgG8gAgkeoRVzQ0Cil5Hak1NNZ2cX+MjSKupmLUM
hl9nctIbQRmKQMaUCezdYr03lsPkJV48ppPAeXg7y7gI00tO7JIwHP86l3/twmNFLyciGj90H9CV
cXhtnWsdu52ynNt2wrWXSrED2vToww/Dtv2nWfCL3NphnY1swJUDVuftq6JiXjTyAJnSXgzejuMk
ju0MOcrAEgI284EWDrD4rTyr85XHvQUXt4bodi5SMZFaSGtBPfx0zezHMEOG4lpWpQDVHOpMmvz0
45cjlqmsjitNCoX9WBpnLBX5msYYeCybAGBPfxH6ogdCmMxG003lH+GiGPiq5e4wZP0cR6C1yBYc
/xUSE7K4MidGcAkYfVRi12lcgcbrqvtf5om8Vkgkg0ACVRH1f/5G6Z+E7r58fqVFAcdCY+QmfhbG
HM3E+q9LuwYZ3nWCo7mslwuwW6efejrV6X1v5dJLM+sGuNr3u62fwEJ3td8/dtb2CEReY5eYkw75
MXEx99vIPsGIo2ElS18fbaLEiFE92Jz0S8ZbAqjYPDoWHynwylAk6gVFmRyBJ9cvtMqhSKUBeNFJ
YlzBNAGVYLzqCP7j6adZdAcFm6wKMVSIUD9qASxHHOMlxGLj5sbGk9s59bpY6kkA2UA3h1WxwOZt
nGZIogxlxGTNGNZA4WtlhhLEcqDH66qQU2YPh76jkkVxRrVpvy0GHQcm0l2HwuIuaGny0nWHOatn
8rHB6IQlw1b+UA0Te+/zBCsq7/3CHUvgahND+jkgZiSCmM20xlxKkvS8bClcWVnMMhuB+W2HZGk9
vMLq648x8xFiZZ2N/qfJ+v3oJaDknkRm7M97aEjM9Msy7mtTBGEXm55MMCqQz9Rd/La7lhx9h3vb
ETY6be7St9Z9qQJ3zx4d6GPr+Qb7sn9c65gW8AjcLQ7POc0/gXck9EzUELOQDTfEsYAsqL5Cqg5e
djPQ0CHelO3Zt3pm1CC8DMSJAcw+QizYO20qfuzS5gDImu7x4XWgsQiVVTmBOUGQIMPstgqxW9D1
Aut5v2rDZuVhIyyiM/C7+Aq67aL3aDwSMtYQp9Tk+M6rm+PlhqWx50CF8Z8mx0M7SDcZpbvM+FnS
9SL0YmA0oanmBofJ8ykjYjh5JR2fOwP4N9kF5ABXXnjD95FtT8RuESEvSJFMekAL6mBtwUfDNXtn
t/pCpNjfPFJQAkutaMPXSOQl5iqwWXjsaksugKo16dVKpjoWr/6wijw8V63QSh4IY0+cxRgnlBxE
XoXU6CnaVdIltqcPA+BwfAm1Xa0ru67O3IwcqWTjoqNKd8+wBCSg8uQxXDc5p3t+7Z7oWJ2yFZS8
F7wtp9suKgkHWU5YdPPzZwmmrPQtNi2+jfBV5r1umeAxp2RNdYDfC47F1x44RNoO0q4W94UTSUmS
sZK5VmBvfxcYttzjnUV8I9Dk3Y6so0nv/DARd4RRU/MPs8QYSK4oBY3OcTU9+AVIFquQ08DmhhZy
qFz39ly2h80O9dSyzRq/vcJohXTSpY5jIh0tNQ1PfcSAMIpa1+J86Xf48wtidfql71eIbpMP6+od
tN7QGJnCpFvtvuwp1/cNn/OjfzLosK/gfnK/6RSbM/QbWqYEQrxR0I6HVscsueEKEOOHeK9K/q8a
nMxZmK3tlcdwjAOjrhW3J0ZtTOeg2BWBdAbNhUr7BzqkBlegMHiCPhIA37q0VaRPSbyi+sC+c5KJ
i+2gUM4cGTkyrLoCzjcvL9dLIxQ5SNw/+a8IxJqcZHJ4XcgB0OkBaJH7q4VrgWrEiZ9q5Gwaz7gr
ik6hDSdg5+rLFSPI44mAaiLPd5AkQR05Vo7CeW3jongi4tYB6J6Cpf8ctjB1q6604khZ6TKuLyq/
ubr+UFIF/jtjFqpEywpzKARSxW4a/pXL1IK2LHx7sIFQ4ZZ0UV4AN0OTM7CfosjyGzc8IXrNaSkB
jnrzw9GRvle1ia6RW0rI4/ajRJi7d/0E/arCEM2A/Lz6xEf1krOo48D2s/HSXie98Hf8vAumhikx
DT1XHZVVE2tHA/4hcnJwRUM/ZF51XRvC0izptLQ4wO7uIJmdlYPEuiUqiVoPYZK8Xp+fRXvGheiQ
Po7tvFEiSDO+huCo+kcmuNR19M06dW6Ub7OivrEKSW++1xw647DbZ7PtVkogDaLGaESdyeuJkdG2
YoOIjka4PpkHS4J7dQu6ZwcK+hl2fDgHd2iL32h+iBOVh6tmqE+bL2AlHo713Ppox2fjwSBj1yQZ
cB3B5Vq/r692RZye23jmwztXJV1Z/xtTrIWqktwJ4e5V/c3CWkW4fbUjtLrjEeTqEQ1r2IFXNCdZ
trewEc/tRqeVaMu6+xv3DYggDibXMxLS83eOs3nMIPU1PsHtAfimNoVsvWXyUxvSZKl/0YbX+c67
MzSWIwfKBteJlAJ80V6fAe9Oo2gxOpTn+EDggTkJpFZ1RpBCItKx9D7gz0ugRr9CrlgKOYJATFM7
J01Lj27ZHFRdCiYLZMdqnzTT6otWFATXNoNwIOM1ak28cCjV5GQ+RRrnmHLBm+fkbek2JahhIoav
MePAgFFacQ5I/kqFUvRqN0C6HysCOFwR6vEASl6UGeXmJKJXdSpyok8Qe8GGcIXcCST2fL3pFQSV
wO3OPIcCSY9HPW+HBdjv0EmBWwIKnsSNC6LJFnFvOeE2/4YsiQGJY8svWLpnbf6y/Y/12I08Dv40
UMXZiOZyc71KzqMQVNCNh00YB62EwKZD9mVu/+59ZFPjKfPIwyKnesBCV8ec4mQlufMi6QZrafgd
d0i8Ju9JxXKdbQazxAaPdwF4032Y/9iVjFknR0PLUjlUgChE574yZjKJ8WaDX1B9aGI9pGQ2OYni
eAI9SnXK76+D6JwkhpFHKGbXu5cJVwPOL+V1j+C878iP8EOrJznH8gVF94lepwZgyHo2AzMeZfmh
bv1xXm13xGhOMWUxeXeeb65ELfi0pJaACSMPKLQOi6EWti35cjZqJ0SS/g8wJNac/IfwSphe6rEJ
7vt9hYlMCGtlssL4OAOsqQu3kSAIZ+qqhCBw+/vAyQ1yGqfCmwH6SDCqoPo8IcXdZJImqvS06D0b
NpetfJ7ZSbu9L3Ybm9wt/gQZCPePcRVDusSuM4jvPze/HW5GxItvHTRpGpi3lYDQHXeU6U/LkW/G
aE7hRWct4Y29AZjc8Qj3VR0+cwqulDujh6PiBIP+0w0ldv1klBr8Wc08evocD95vM37VhYK4Lncq
KGH29bIfzqxzUSVh31w6UkI+El+u1jWvlcfThW6StejQI7sjQ383kFH/TEXxeDkk2KXz6b5HxFsn
myTSRijjAGMZeooeat/gpYqGTPp7yro9gj/fZPFNxK01r3V7D0SfWydEkuUlDBOMXGK/hBxv5zMY
3gmSQBxJxaehCiIL/mzZLcRrEIhZSb75ky1+87p1cuWo3sWcz/0ztmq8cbE3kqs/bQsLMNnykQ6t
XqU5fwuhVIVnfo6rOUdBWsmO3/b41I57Rjw4TTCkQcvROVPz3K+W5aP8seBj/tt4gB4OB1w/myhL
g7yGYq32KKvGVIcZT0kM/Wah0fo6QVo3Hfa/m5osTQ+QWoradSDExo45Sv5S0PEtLX6J78vQD3Pv
lD2k3uekiorm1QrHBAKqaFxSLQ8is4PYbOSjHodn7Hm48N9wDT91a48QJAufy525Zu/f2p/oXfo/
UoMhxCsgRfgk942EjQ2W7XoKKA1nVzP0sEStdKWMqc04QwPSv5IAr+6I8VhbVenzvE0pRvyGRNr3
S9nTKhiS0Fy9AeFLcV+h4OUri/je7jl1CxuLoMSyPYD71lzYQZ1DE1laIs8KPCO48t7rXDoNMqvy
r59SBs9GiolynNbFRjezwGD6plPoub7ygGjoyyvwSuq31KG/mAjaFAjs4y7p3IxOoBRZi4KoRNZB
iOO7PWWldAQtlcHKKPQc9a8VRfxP79TzVPDchygGgasCfFK4VM3swejsKknGhzUNa06aSoYZ3KjD
lilB4mrSA318cvRe50aV6k8e3iedE/eYgBIzgLifxqD9r3AgixGLbXxz4PyqYfqFOhsVPEipmrty
/iYvJDtd9lUl+sM5ohFlfldp2XdMv99EQ5JgtKddZLNwrF/03wranoY227Tjdgr9XTzHKOBDvzuD
SHnymTWMw2nyMoHgoTNB00lgSz4HWxRr2oNn896kDTOq0zwpPjtUjqsIyqGik1CI8shE6ScumjjJ
Q2C7ZtcBsymhi4XZxj/zjRP62EPkXynibb64LgA0rWKx1/PGC6AXB29wF+jDdMmkYL2L3ywwz+aP
IdJrkggH/mC2a2axn6AqsNNgYOBvGzcp1ai4oBIng5lDkjutnLoW7sep5B+WTs+G1A1Lbldf8IYk
Z72YHPBkzZbs6IpGhdKmpnbF/TJd5ZqxYdVFO6EJFsQ4qyOwLF2OtXy3JH4fYirTUHSayhdpJJ4I
fVEs0V7K7bCSOY/+8FVxkplkpJ/FlkDA94M87+5QtbUP8wGJRLdp2+Mfi4ekSJIeFnll6YHm0CrR
1aNDQiklnHdZDtCeZGHdlyBv5VfptUIGBUFNig6pSJk2ewzd8UCvMLj0m3G7TY+4Yq+wkmFlwt2V
toy9Hjw5K+PpE477ODPTAu7Gz9Lwr31k91QQ0LXwm45THpPU6jYbUpeozqL8jNtB1DLCnysZObA7
W9+J7BmLPbdmzysIYFSdswQKAAE7yDNuTLBLbiQj79YD+Fadz4RauPQqZ09xsc6DCYkTcENP6mwc
8wAceS6TEXLIaJBRo0q/0rX2RW3dZ5VMh+FstOHptty5HiCYOiVM4pGMHTA/faCJU653MjVjLmIh
el4oICqPM4yFwOhMMI9MbayYysFd7Kj16M/qhhdfyn9UPDwHf2kvj1O5VHd6UCeoXlt9o4l4zd2p
W+1zKq/jxkdBceHdaaVvVwNYGBfio6IbF8mjq3GDFYleZy9ey8RbyUfvLJoP/ls4BHEf7vlYM2KY
eFip2JuSWqy2Jt0DIMAITZXHIhj5OOaWdy2buDkZCe8Q/oozMPlKV5+tZpf3Dwkn40iTrHhDDKKV
cw8DrLhcwyaEy6ym2FUPMddKneO4Sy0i5HM8UPPRaj8I7QOGoibl5JYNVoZzxgX6rMKcVbJJ/Rnf
0wWiuaLMFfuFehaxA9Bnj6Nq+gIC2YyOh8fzibTQ1HSduslNDPpbdT0KjyHA7APBM8hVNmkY3CqS
ShDZ0YozagZRREek6/0wnTsoglLhN6VWCnE8S0fGGVe1zVOI7kUE37yTBfaBsAWiEAVC3WERzP9x
bD5KJneZMhF6LEKckTZTy0st7MqUbG5RdLeBoMA4/HEUrjthY5dd3sFb4PFyceWOGQ5p14MSbRF0
IW4JH+rB54g3a6Uzi4q/9Nf943+nuHqsNu+4fOQYLweNhBdtjij1hFKlmrhkYai3o6HO7ieTGJ/i
gZHeAgRubFZ/lJAYD+2KJ0DxOlodVGoQkh97bqTk3w++/df+Ppj+XfIbjFTo3NkVn8Q0Fdy/Q/bq
dLu+dCLXkCEgbx/7LpFY/jh3Lh0iRrao6QME6os7AgoavpWmzWc9NXmEgjR+az9OavWiidJCyP9A
1nznCmvj6OV+2L/ndca9YWwvzHmB1rYvIDGI9jNhQmmgjYpCjs/Z3q1f0bgvvU7p0XbiMmS4vD2N
GaoFw04vGGd8lzABKdIjXhxytZtXT1JeTFAwyn2nMyOC8MZvWFUioB799SoTj3GfttiVTqPo29Pl
I8IJagvcOVA7RShY23Ml9k1ks1NOIe7YaRmQ4n9yxpJ4eoqIfnuuTLGOhNHgWdkfvPO1jU/fJutG
MHF4w0TtO+Y6O4ga9k2Ee/RtyQSSOQHdrIqvazUE/0RzPv+Tv1M/dVD2lF9ObwOlbEsIFkMqOMv9
yAN7/BBkvd4c4eiHcrJovJuinQ3h1ei5W52inr/CEZYuvr5KlxISy1jNrEcJwfg/PSlOz63rzT4z
00dcW1QsyWChP+KXYsJwJ+KUEPeof+AM8J8r6Pl8Oi7fqyNA1C66qd8pFroNK/Nw0RdXsjCrw0K0
6L8xu4PxMwK3bD981y8AMNuK5iX18d7Wm7fYpnmtMGOgCJbTG8X5s87MbpeW00pYZR9anXyqSXet
wani+quqXDWzcxLDLVbE+rUhxN0jjAYqTL5x4bJV2fUx/i/e27NJ+Rq6Cxg7IvQt6zTB8fZXCzY/
bv7VY+m3/HDkpPAlh5niP/5NhiqmRtXkPPoigRh6/8tOceI081RMmk3x6WrJXZplK7qxEYbC6dFf
YMLn94oFP2jO1QaaaZEZktqg75O0rk6lIilx3bq1aJkWVcCtA4HsYVvj49S5iGKAy9OzLg9oFfiT
zcqQVruMCBd0GvIiv/wm5mv1EW/jE5njqtnieaJJzfyQB6DwAfIjkk7UedeDcCrX3qnil+pmgzy1
E5PU53HLDqE6ARkq5OYGb1OYn8nCll3/jL4i/W3k8Lzd5KyRFE7HkLcz/pbceNRpCC8ZC2uNu3uP
5M00wtrpUM8CFM/db546ACRZBH6Frw9kjERzUkKF64GdxAvsKpn/+5s0VP7wkTIJq1VEZdQX3zun
8BSjvnXFh5cPeNM4uSqqdrlUcSwZjcIIppDs92GOBWUhqM2pJMtonsPHcN/J3OJQByH7jZtqqUhL
sdjyaDEtm0ZrjK7zVlZUViwEGOZIGKSJ10JF/ccrDEnnI9AmJVvGhpf4TufTWXQvZriFDFhK2oLM
s6eyqL826M42OAeJ/UWGrlpfXBcyD707tPA3xupKpZBl+AoSSaqaWa9r0u/l5EIdRNKd3c4M08L8
47HqfHP9eXije7f32VdvfD8Zs6GUuAxZz81etE+Ptjq9ElqLtfgKB7AsWTPYr73GXZHkbJBFA5nX
kSujuGL5PLKLGDuSdnWMVSsgwnrEnOg6jz2FuICaXjgqj3b19jAOCTiAJ9/hKP8KpO2gcxdXVx9D
iFEkIUKIoKVWeiQ+6UvN/n5h2SNaookKlB0AEBh4ECS7LVFfmYERqDjsgmX/Hd6WPgfDUarnXzWv
IzpfQQuGCcz9ILKNa6TkaH7CTZYBwRZTMpkjo7kzBlJTvGGg49Ki0nLJQfjSs7oQIFEzan3ifWuQ
d4aHFs5ot5d+IfanG1KqAh8mr3D/nBxEt4v0gZeioA57WvHidrqE94gf5OqgTBBIAANMdGchtA+G
2PgkeusDTnxJU6uKSZqdIWHYM7ptV/YlwK/frDPb7mKr5in99DBQ5hOFrh+F5ddWfgNbvNHzJk8B
I/0TNf60+ojSvnyeSkISfCnui0oH9EPx3G7bNkSwPInzDH5mNC957klhwAQzFGoXpQ4GG97Aviu8
vqw/fO4p9CaX9lefMMzzj33lZYoxljG6jdrIxyuVZktpFE1fq5yDvQMdcXocp+vYYLaM/VMW+5T+
EYwuU163X7enUcFhA0OEw2X0lpNmWKWfRxEq7aXI9mvEqvWV+51ErUpoTzW+OFIcvnKVhTU0lAD8
Vhb/8rtGtbVNuboFhaeNo3ntT+ckJA93XsFVlMTebHupg8GRAxCRsajU6azEwsj+jn/UW706pt+x
q42az23Gu46jrTWdNBydBHu4i/Kq1eo1NLweRkb64LReAkMpUARdSW4wZX9B2sg1oqL55OomzdOw
nOst4qUBwWanK/Ywru47swF30ruNhUbqGzN1rixcYbtIo4OvcdYX1O5VZ7j/1xZ1GmIn8pEG/kJc
+epRhYuMd5y8+JUfEP9q1uDXET+CGMFC7ACD0hu7f49NuNPRK3pCuJl2JS9YFNChqiVWygvyDm9f
J8WCxzqrNsdbS4SEmzdeoFm9mo5LYOcbNns8q0WYPZtzk441mG/8tOQpPNjvkyMekVNEyaVzf/4y
2y2+xGiCAF9ttthMyE+OUWEADegsgi1V2vcOhSqFmhFhJRtLv/6UZScP30jCp9YZY3xW/KBN1KD4
RETpNQ1td8SA8Y3SGomVFukrXMyC5uQ0bi5OnTYVF7ltw3H/yZjscymn73YjFUwQyKMTXjFtBOrj
wwxzkOQ0ThmX2M0Xk1iIsvuhtKmKwSylfuI11YMoludLyfMjJrKk5N/tKmC8YI+zDRLwho0COVVx
e1tSDfpXh2dJglytxKEUmLPhEtT6j7CiebmXgcrxiNsQ8kZXHq85vJTjhITXbx2BPicuHgfBSNRm
4r07rwnznp7sJ/QgIuX4xe5zuJ0ebxs65IuRtpk27dBWpZ68a94Z/+UikZ8a/yw/1LHw1EjJwLNv
rshGbCsvFpdKGE2VLVmc6uOwKdqFUMDdcl/KIv9+QpBJTKtPScNt6JvCbv6f5l8op31oIZh9Sw4S
QMNuo0ZFAwPsBC2f3fZH6WdW+83IxCMw1/ItdX60oIp0J46I1ixTKv3wqnnwNbqEZ9HEjHW1eMQT
5PBlg9vFjrnPdbLenk5Aw/mJewYGiVl1byYO04v2Noq2pqtba5zFxQuOzdFuDqgecmHSUlfmSqXf
f2l0VeTAPhpArvjJ82gRfePnnHW6LUQLQEA3vISS/ZiCqBYlxkJi7UBMoyH2DMnwe4DoOIPO0qjq
RsIj1znMbHUHm/cuRlqfKPU5JoXu2w1kHlVtmO/lsgrWoi2NGHyPQ39exopGCp1kvhYDt+Ve3wVS
fhVNtBVLY8rOKp7IiY0KSGLdV2h66ojvIS6WuJ6XchP8jwFPZENfq2VboyOSspuskKxz6QVV6IYk
m1z0+2QStr5uvPRgkU4th8hVxQdO2tyEp2/3fcNbs21cT8xiaAAESklshaLTRtOC31rHPldLBHrF
bRzN8pZv/hHwJa91jzfHocx4URwto30mSH7fWh5dKWNHYCuLvJK1kOJ+J9X8XW4T68rsKOfagewQ
gNvkBegCMwYVi5THNy2YUc4qn2MC6a2QsxKiPGmOyedlwiZ2QxyQInCElBPI2L0Fi4e0yeq4blDw
CQlDXSobdfKKi7Q/PhKOGtFkXIuTGopJqdmInl4ZIJwbuVRdv79ocgLQfp8qs7FY26FP4TDO7GJ3
/qkgi8FR6eTnzM3tjgToevSDKvANyLFPEGnYuKzwd7Qn4KlWf2XqAqQALZ17Bi15qoCEatrgULXW
vMpY+BIoctIdEqNePQecAwj8R0g5wLTUIDU08LUkzsg7rRzdJqRTiKcq1VesTZg6aBW4ot18PET5
NGSroAU9wYQfGqdMYgq7iGh5kfmrBZ/7ps2KfuRzg+WA4REnMJD668hO3cZvmT43SY3KmilAm78O
Zer1LRoUN84WSkyRDZAODVqcMoRXj6g32z8bxuArGjGfSAJzRorO/C/K5l+bEasnHlQCC17QoNDn
R414oWjwUbVwTdwstilpzW8GmDbj+6FRb6qe21Pq0t3+pypOlfhXoSvp2NSX2ByjXp9QYwUZy9rR
Sit0b4X8yhBnd+E3Cqt+h1rHOt6kIc62i950HLGZwmKbO2oveUuQQuP3urKONBQpQDr5PpWZC72E
hYkQiuj2PEmcVQjSzW7Nsl3HAlVjROh9MoZFjJAI+nPb2AaBxp9OQ0lvTChPpU3ebddamnbAclI9
/BBKiP0+Eye4CNW1CAoRfKOxrATQepSLf0TuoODEmzM+SXfdQ2KDiNKBQ1EFcCC+OVLNqzXtwSpN
adFNH7gClngEWLqQzxWMKVpYVndHgARzaVfJyDN4ebeXBRsOovP4BNyeLHgjKIK2Ow92vAfkDE0F
3E9+fCTvBQeGfPxmRSVMKnfYjaDR9ZQET7+q9z0o3u8vDUEy6kRdSpFxjnkr3oNXTULAPUgQQe7/
5kUthvBh5JwqYxXP78888KVWr/clHc7/uI9YDXQEOYwWzzBMMDvwp/kCxR0g+8HEZQQZX7ZInB+I
b/cbLZXK2wt+ZXDVA1H1CYmGY0xafSYVNROX6ce7Go3Vy80owEFunlKyzFqOBCEW8TeGIt3sNNsX
bFGISWVQ2gZWw8unFW+fVjefIIZuFFSYfFzrVq4ZqWvGRcbVCZMUeClkt1eJddflhhmPgOMB+yWW
mS+Ox5qaI7lYmEXxdHmqTW6bXtTJXuVC+hi5CUI15frHM8yK1C6/aPju820gN/KxSGPbMjZKHo81
t6CvLYOhZm+WK0mxBdyCvUQGw7id/47HNALTj7WzRPCYe/ZGBfGP/Zk6Bh8dBZ8t9K6MT4mCM4hp
MC1/Lset4s4fsJsPjoa2yInKV2Wzeh5cv/QYAf1cgPImahdBs2rUdXACzPkxsRIAOgzhOZGtxIYE
zPcxdx/kBYGzlvtI1BtzI3kU67ggtny8juIvLNXMrq5aDJjva/Hz6qyEOkMRAROmlMybduxUgMaa
Q9yOi9CVfPaHBr6B2tPonTwbM4BIClXsna0S0MWe/IzgByDrTnHryXXc5iQOrPQlEKJeLMJ41Z/l
Cs4ENubNod/TMrq4AYEX8K1jvmlveCIZCbvWdQenMz01tRgOlcCuO2lHSp8oldnUD3QYvrO/sSzA
e/QAxLoQuBqwgZ94rjhG2ulSbLKEw5IpGjPXYpocxFKwitZXulq1Km2s6SvE3bbFMjFE5q4eCqq+
zsVGMUTK+3oW5oP7iqTQYr4gBRyNF+ZpoS0DzjJE6xiUa94HhO6mRxtOyECHpfWvrl1qpJ3j2k6h
P4AG05iEu31QasSX/x4perwWBtKJE3Ep9QKEM/8E1mffX0BURhzHsF5axiMAEPp+ju+0VnKbEbHh
Jf2nyV0R/kZI0Qe6t7MP3uR64+2axBnBZskSLMgIhWMmHjA5NX6U+C2mz0p8zc12sLWxYV+GOR86
EAwLJv7ViDWN96wmda4AKw5W9h73PMrHPRvKtxktPVIMvKnRsOO6Mq3WbI6UcPfEoOlSPHT0IfS6
mjuB9+O0dFqSYKK35mDIL8aLyG0/6tDuHEnBpVacebAWEFPXw5yJACWi8DtS105VbbIesF2jFN3p
FPMkaWC++6qPwbQ7eK/+W1bfQUf7CsSMvH3R9sk4hGhL3Tu1VZFsKp8l/pbIDlYPJAI9q1Cr3UhC
jaDj0A97P30bbkKOXNmiHEqjERxHhSF1K4imGeVEwLrjRTxJOY528WbKB73FryD+Xmi5lXQnvwvX
rdllF3o/mtZk8A1K5Vx5/Y3Go28NidJ0Sca2zczn+hX7zkbc5XN4CzDygRlx6Ye+Xz7fvtHo0hV+
bIg74txPEZGwA2gk6t3gNSpbffrm2iZebn7VE2VOlq8IE2haqL1zuIx9XHDQrzmmtdtJSnroR9cu
Imqp4s2Z36xZ3Gb1QDcOQy3iwNE5XIdLrAYKOItuJIoRLM/NnVcC5nxltX9dmmnv0n8w5YqCOKl4
1xc8wgjM4Bd5QumEWpkFTZOOC844cG1MghDbgOIp1zKYlI/9rQUpnosdaXWJMF61rmbYBOSOVUy6
PMkzPsM+sWdeWMHIqVduaEA+6xmEcjT1o7F5v1oNe3WSkxkkpOtPOnD5Fgmyc2wpq4ThD1pCp3vK
XQdeSPWV5gv70ZWNAPKbGsM8C2CJ8TXbYTcMMGVTyE3FBk0fvdO5fBeRjtPXEHUIUXAt6QHk+35C
34/EkOVRIqcYf3FSQUDxXdEWtBexnhl+Pj/Ud+Tl74zT6Uz6tFRJ9X1pyYDZhkL6Rz5Onu+Uu7fl
hXg4WRUcnWiJTfvyz1fXeF60+ACJFCEoXzPq3DmHvsrVfhkLQBYBaeJckRFr/v3LJlu4hdA5pIan
tYRvPbxsUrbH/R1uikb96wfptneRF325RVnSauLvFS5sPrjOryX0qReTMAVDwtfy+Uv91JojG0f+
k8SYhbqFIBPoqkBKgdMkRNovZ1vhxjUlnpfdJSiNUfBO9FYlMK6l2QNYuspBnTkBuR8l19K06waT
I2sPSgEtt0cR9dPXg+BFQOoMcSMfkM1Jp9vM5qpjT1V9DIcdbjxL7+p28QDHHTjMxCsVDReePS3q
tbfs/QFc/USacIxQ1tQtyFLy6g6m5RdWWTyL2EndeLRqR1Pn+4ynZQY0EDsQvVmg58ESEIrK+RjV
jUrxXI8JTcwJAHMgDUTABjVvfUQK+Dh48KwYZO7ZmpWrlIhG2ACS0OkdqUKf5uK/q2j3F0sI9bHO
iyUoHZlby+7fno8DDKDJIX6KNIwbDWY+oT2kQb+TqV9q8I4DE5khBAKNVulfCRsRNQIRmMbtRAlx
725/jxs6DU+8M/+x8xNLOmwUpxjUhyGTvUuPnFiH+BQzJr5DpRnWvIuBC7nJQMucdEouXb4IHirJ
zEotz9okpkvfdLwBui1GUmQ5496/H1k9+wIOauH9vHvhkibumXLQDCZlzrpkHNTCFfeEeWJIzh/k
6b/i5LNe2tvXfY24tWZ6MjokMcD/88ekvxgBx6QEyGXTAtyvku2kwobjoGdyYCHGopIfs95WGG6b
3a+G43xad3pJmmQXNYcjy5ZYeV0UjFzIjEr85CGmWsTgg+eL5P3f6jDstNh1+1V3ooV2ewDpydA/
xksgAmB5yVEUygM+v4dK5ex125rj9FQcbUHm0baHZzlQRjpjOXEweMLTevrWFkmWtiF/KfMeV54X
BpPdw//lGmVNyCXHFT+1Qp+0DuAcSfK+ngzzslESPZA0wVyjDJvONlpJXTaFcAlZx2N9IdeghhgN
jIqsIuUsKnjPsgbtlHsJ5GegzNZkYzM9tEkMGbW5UjTuoWGuo4qTRbuVGTOJ5Jx2uuqBNOcWVno0
WgtFnxjO0McSJeOkMqK6hu9qaRyspSzdr4y8g/rZkeu6YCDCnTctj0dJQr6wcDW05l9DpTWiIvXk
d2WJFkbX/q5FYjE7O0LSJI+zEaA6N6tX+7WrAIBcFjVLfgsf0mfbQbyD7RTDPiVC+g36Dz96andL
wzryXjfwGYch7WEgmzGrT2amKqS+9tGOeF6TRa2aea0IKMfa3EhskXksZlQSI+TWgXPDU8rt83qz
WtrpM56lpyFULDJuQX0uUJFouFeYjQn0Fzpyg7I/oWgur+k42UCOdYpDZojmGQw/A8pQOhtGIopM
oXxFW4pGm6VEuibvF97cp+Pi8np/XfQhDYcHPYueqKVlqLH1MrJVzONV3pJn3qUn9OjWIKGti4Qp
ZAJ3X0FxcVz+HfcAZhcYG5ub4ahxtFDtszHOGs9tDxAhANKysBwUK0p2kRoBOJ5ckbFzIbsvrMkv
0z+km5dOlLRFuEoVZHb0XNPVD9gVWJNgfbrzf8wora+6qkEu3iqfNX1I75lUfG8QIg8cFh0eSs0J
DIeGr0xrZbGiYFXaKbCeWmoHIA1dwgWqXRRvQQPel//xYgnNObB4aadbZ+Ca75oKTfu+Zk3dOQ8F
Uu+uBph4+GcBDQArtctgRinwNn7jQtqisbZuYQ7PcWo20fEzQBo6zyWPRVsTyESyNsTq3xmSWTMj
P4PwlfzUTs4P1Q1DISpAeKNRYea+tu6yRqFJ+c03t3q3jrOUP5mGXdr4/txnJTMkkeTqTWjvc0iW
ozwYa6m6ih7/N4htsXkZ1K3anN8m2GRIKftOWFVOugoBecDNzcTp8jLt3STk0jgKd5SfNX1bWM+H
VxSeh81lovubudeuMmbX+Q+DhB1IqaXhSWSTsddyJPs7G8vhzxUNQe6eYm9peDuo8wP45Or8QehO
KyXPdolxgu2lQEBhDrCTyqpKhcDqmmrGJoIHMdDVFnNYEEF0TcbBQbR20t2HjQ11qV10WJZM0/15
lju1m55Tf70Ja/QbODEKM+3N4ZflK+RB7OfTWmYerb9Fk24gE+PfsonsCKRhUl4sRgUlH0iXYeQF
ARf7O7qjycRGfioAlR02dxoAiCE29lvXaK/z6ApSsFqEofIYg1h2bczGP3xtMdg7E47KlcwTj/8O
LKoy+7QQhs2KGFU8FqF8euCtvMMiquk5c1irNpTfZk0oC0gp7lTuDxyw++XGo8SINhqi/K9gNAst
Q9qXga8RRrC3DOlTDe3vExyVBqg4rRh0BZz7ggLB05r7eqXMkgpXYxBiYCw2zvQ4VXgEfLbQ//ws
EFaXxAoY/MCW0khUZDfYlf3d9MYTIuYBKu1xB8W3GUqLFovKw4oMSeoaGlDSeQI4MxNltlMczT26
YwYyoEkHKISmfkHZxvS6jKFL6oOLAr14v/b43p06KQlAW6Jq+6dTwSps9ChcsmumX1wEY/99Qm+w
orfQ4/mKyK+o5AN5hcHnAjbt+zmxwUq+eDDPYiZjMzoWBAdSziS2OP89kJNEnvIV6R7fe2U7VAcC
L3LA3Uug4wMWfAPhlvHGxd/jKao7xNHXG6hJR/AQE2yUJ40X8JbTRFM23LuZtZHztY+71MTGAl/z
W+roRHeFMnUeojR4NkCDCPV/5PYufrWFRhD72gngjWNIZ13KOAVInxQyYZ2jxkG35nUGpwdCackK
ePf/8A8Lv0k4cehqS2qvU5hG5Hci02NnVSONTEB8Bd8N+Pf8UhnDEAyiS+zYP3vUFNSxGKntVlZk
8tNbB0RiqhI1YvhhXhWO9SCbej/Arh5aTZIpTHrmQHL1YjDx0dU3h5sJt4YKa1nzlg6bAfdlJAO5
BQeM1InC/EOVLJu3EYQB1SWKM1vL6odIBeqqYR8x2C8eIlcItEvSGXkvYhhAjNG3GIl7AE+/OQzy
gcvlOFkwzHPrM0kL96RH7VstP8WO2WDV7agZGq9zzcnipKxVR9HHqGej0RFhZBoNP8kTokCX/qZu
tR97Lyq/sxtwTe0cI7qg0GrFdnBFB2C+MqptnO4esd3HgQRjSXxf2d0HdJtUv/ffb2VZPqJaJEFW
kS+KA1zjiphU+R+YdTSrY4yHcf/dBENZ8QcbGSbRAl3O4jewG+sok6eqVSaWt+njgt/oQH7B9o5t
aA7Bf7fw/oIdtjh/S6Lix24vXz939xNcoqt4Z6OLQZHe2O82f+o9o342FMqhRmQOFtZeDMpDv9p7
AH1uBdBarRCUSi+2DGUwe/3XOFxA14p3yqqH6z4G8kfNg025zqdbfV8YHJdTxqmbhUzclfzEbuu+
q24CF30WdGb3EJVMXYoGRmQ/f6kG0c9rZv/KRM1yi6bp7bOWx+Zl0zUCXKVsLdyY/Vm3R6yfR5fn
7sJC4Cl7WbhCBxK5ECsSsZBalJCL8BR6VSqvbDZD/Eb8rYsRuTdGsR6RJy7il+nA5HTaw6ysNDtV
7zLlgy/iobf11UlpxdsdXfxhsWyNpfxvhCqmw936W5DxUhurcIMLAgw3FOmMA9zsCQ0IL9+9J9JW
o07293D3VXfHVMnxsDF89o6WOTO3vlNCc1lKzhLdJFIdPX1C3kflS2kmQvZ08lpMjRZ+0DEV+hfm
/xjWVTW7fwZm2fY7amGMGDsuKBMk4qASkfBKzbQ/SabFnLxM6dw3+viDql4bB+A8gD84N8vcjUJ2
IMj1B594Wws2iZigLvq87WKz1UVM/sXzIspFJvRqyD8jvE643C+U5cqsMTczdP+M3B8uGPc79MWW
1IvjzZtc3peUcAerf1crVqbo6z1qDTKPC7pW5cHz8+dnr/K1Xb+/PKMN261Eh4242e4Ok5W61UbT
8P57LxQ4EfW1a4vswpCkOpfUxGFhmN4u9H6B/T8+5mxjigYagND4NqQU8hhcf+si3b4G5zhy36oK
3zBVilz6atiuxe0vL+HO/lq0lh2AIPzR9y49U10bgdNOeVRnsEZtmz4m5+m3iSJABqbnH6yEJfqF
QhCaSP/DC/wAOpUjUpSHnyhkY6W053ynL6OQg6ExA3+M6FirroAjMulhVMlcDKVL1C0DBmUyGoDI
7cxqu2HS+CDaI4RYzJCCX14ZcyTQnnGLbdDrd2Ft/iCdVe9KvPMX3Rpuso9ofW2XrPt1y8TgaCCp
f02019raUV5NxDD7M1CrLrAcp3AehGZWVpb8++8Bk+Gsdw1s4/ULgJ97shnWlJrltH52hGvgtT+z
g1WQd3ORkF+QRQOch6jvhVDkJZwuOVRCtl5CG0vK3wFtEncfkTiUHH1woBktzXjJsTTHZv8tNkpm
bwZH1x2Oo68cIYePmvEQPeOFgeimVr9elf3F3fTp6Dg1N8166BnN7VsqlsSZFE8jHU25HiwcAnC1
yWDd/Anw85ckMOxYdqN/eHK8a4yeIS4nF0G4CuIT4PVhzliL/KThiMnKknjMeiVR1lIggNUxwIhu
GdNJZ36E/eCcOeGTrXWNkN/Dos2Mys8s5fcIm0nEnWx00J1WNZLqsiw8PXE+nIrUEH7M8VGDpm4/
vuGpa5tIkJUhpVj3U12QUXffM9g5rUJpiiIHPIPs3h04RiKPwJxgGt5RcIiXfHgv1S0s8a+iZvk4
vOI+wbJyEte/Kq6HBvALUgDegWir6ZK2f3F1AyG1ZIMyRW+uVEvNZxM3eZNgI7VzhE8RF4ukVrZZ
jV/MR0EPCbQsz1pTFtF/6ASTqZMEZRjLtMFuKxslRk1X7xzsFf2z2EnNYUoshj2S/jh7FqG2YYYH
LAEZI2r8UGvpd4rq7CCap9rs3gF7Ovi6kGdVc3wbjWj9/8ArtbU6OiCakfMkhJJ7R0XRIpUupv/T
lvMyDmyZOvFfUAhtXjFaz5GosVOXX/2EoBxFEh/aFXWwAKMbGYUCiuY+OKcwcq43oDVfu3sc4dQ7
hb1pT0N4W0CvQ3+ptKoDGCS4cYQjgXwR9Yf7/zrUWI6xoz1A+kC6H81rSlFmzqv1pbuMsQoZ5s3S
qODC5Dqq/E5Sf5cCbvT48AyTE0YxKU5n+cWKKSSF0GAlj0AqfWG2Z3oca1utWQnj3TD+rhRB7HLe
2wHbeF87MHLAhAlNo3Ta5mxUZSbGhQwEixF79juUKqSM9ALASkjHL+5h+kqTbHSgj84/Eo1u5CLr
yIzKN3nkxZVtp86zMivQaTZ4hNNaIeRJUjHe2zFGqjLmNCv6xALt4EZd+oh2DVsJl/A29CqjoXbv
oSgjCaGe4tUOiw2TNLZAXUYRzoxZtc6FjmEpJeEPF4r2vq8J88vVVx36k9MgyOACwsKTqSZmHiVd
L+BqjBKAnWL2hzm5TySKesR0ejUyx8N78yb+XcPipKTEgsSG7TCx3mvSSBsFZnsXY14hXvP3WPtu
iqz2ejAtuIOwSjtDkinVqxAoDSxxR2xHo1vtqr4LcgophA8E7ortvmmLNcS+sO9WdNzHlHvvCtq8
w88RDzQ+uEAh7+FsPQ8pFUfhL3isX8vpEQteTRK5mKCJNPAGw32hH1RY70/e0ZfH78rhHqK0d5GJ
UmoKKk5Ps6mfFJnVHAClZ66s8wawUmn2r5w0ehKy0nkscFUkCL7LgZp20IB3ApRtE8zGddkaqck5
YdiUhY7sxixQXhMc33N2ZHXuZEdJuC3e3OlmShel4r7lXulG365D0QeM+jDAVg0pY0sW1TnGYUqH
xq1ii0NoYmCDZGwjFGbOQPK6+fZBj015vK8R+EpA5UHosrl/MD10c0L2Ambd5cAia5gSq+St7Y/f
+TdJNdhlrooKPkTE2lmfz+LmxZs4k9hgjYZ01j6SpXtHTu4663SaLariaMwbbWGssHZ6TqvAX2pm
MDYpzKKmJZSHt0UC+11V+ukx4R07PtW2QDQP5Q8zwS0JGrnAlkO9s66J8oJGpa7JgYL54IO9Aii+
CEbKudU3DgqepS3n1xYfSQsM2oC/apgfqNZpWGzoV6o65ONBrIu06e4cZh5FufZOsHxKGOQa2eNw
XSoLCRtl5gkD4E+bD0hfl/1aMkHTSCN/VsU8EuslggqcW1kFiOVrZLZVfqhv9DM8nAA7nfhEf7zw
TUP0/mYajRQXYtF+cUZzjDIUgAKrTWTFpAr8RnfMCy7X2Jl8xF0F4NL4OuSSi5lr5G02vortVxPm
yRobcpwN2SvJ/XfdPpi+ltYuW1k+ba0Pxe3/Oj687xjpWngmfTQB3QtuFRL1SKguTz27lBD/3emY
U9denWk044qdtddVjpOmVSOHQr+L1k8AHMmoLRka98By4pS54d8HY3ZWWH7f+D033di8Fv41qnrk
OaOWlM/64QpJ14F9UVMGj87G+6FX+eSH7Vod+SmOCKmA/5mg0wiFP4OdTOz+zmPQ1+fkXwBxKu+9
1bcD4UvzJa5Ef+4IQIo84O95WQjIo+6EHP4tOKxaQHd45A4buvSZy5evjwb9Jx6LcBSDcmlRO5EI
k9/sq98xCt1nv3/gEpXz0lYFthmqpWlcZvboWAebziMk3dvRIA0xlk4jodpnw1vfz5oQT0PZS3QA
t+hDUcDEmQwcuub4p6zO6I4ZjaY8z7MzkjUBv5ysyzGrlxp04Ydg+Xf58vZR18Ts0V5LlSzn3Df2
cle02vhkXt3YGGxOcZGx9+xJPD6JPix1YRQAkrtjTuSJvGmMeQUfSLDdjebLzbX9Q89C7odgPr6T
qhJFHNV9CrDFQPyBaghG/9HU2axhW0rhT7qoE6+yqmDSXdnMKujx3SYHzE77EXRYOB7hzRPn2d6/
PS/kp2KO4OetfJtOD6XsIosvdXI30o6QJ7tsH96Ol3fDsBOC4wyVA4JKCw8OPNYX8YNuQ2pxRYJJ
o54z4DCUIKjwp10qgAZa4/1L/D3sSGxCYwMLj7nSYTB3AsZORcFp2gnw0AhgGk7rXcWE4OdoK57I
1ZHIbfnPcEAgKjxGvG1z0T5wUaT+TmbHshYnv6ba3AdezoqCZlmHorlLsfhD+q9YF3blVASKzKjp
tBVhB9X33y2kkjP5jI9A9hXuBdFyRmkDuME9orkC7dUmIZbvOMbIAxNqRv3Gvlz3mJNIh9S9MpQ9
h/iGCDRNN0E54oD03GtlJ47Hjhh3apHTfL0+i8xpRPHlHnDonDi9v83B869hd8Woom5OKLMaMF1w
8Xd8I15r8frUjMUHs5KcnTTsQVHMVWknOmlBMWS9EGfC14206vHWPqAC72C+dbUFsRLl9FnIKwy/
7oU1iYlgELq67id423HNHWYAUABIVUwaJqVjvChFFWf1ZlvSCy2sdp/ucjsRtZ+WIgwooE7lmIj3
zzZcq6F1gr97YLjnx9UxGDIjwi0zA02/LHt1jCL2h1koNG/ew1HgjbU0BzbFRHF3bHik5wWvo4Qa
azAzsjiRPRWyXqagOfzkKjZ7Zj/7Bxi7cOqd+rO7zCPvG1iFskprLCjctBryeFKr4XieHGVsrGw2
6p1gIZ+mm2kKPN1acyrHu/py2n++Jr+h65dsD6g76OygNHgj+aIMmqlrGWgT1uWeeLA5J/4ux9eV
4dwD6gaPspJ9U4HCaZRiyHOPzvv7JvCND1ckU2dy2hBm5eiEPVrn/W6G0v0HR48+N3BwAO5qeDOr
y5Olxg/QB6eEE66nGZFuZa6nzWRnMazPlmoLNg1IYLshS6KTZzNp563a5doKqKolAl2cy3Zqg1q0
0gA40ivKIqMp4+Bxpz+mrodlbEwdXiEBFfjTTBwRnvzNuQyc7h04zS+tK5p4XDnyV6gah3NYe6WG
0wp/DfklbTi5qUB7mEs6LbdJH6aqK40LOdCIYOw+4xAXE968bsIHo0uaDbxMZdNiHWqkK80zwGl4
5VCKNMDf/MH8IrH+75wbEjwm9l1wz3Xe2AXGsCf2KQODSxNDFg/OncVrAvSDDbpMcAQnBuwOLVOp
5XFwn1UkXGoON6C/xbxVkjHZ+KoJTSr0+9qsFbX7W3BrdbIrnGQ7YB/PcWiMNslaVugwlmtmdspC
m+EFzbxRkmE6Gjr4gQ5hp1wPZQqMBHf/4Wb5mQqcosxLNOlw7OsvRLl2jFar2638DjeNgVDoFc7Z
f/5gNg75umyJzItY9dPWlKToT9M9OLt1gPX1vvO3Yuo6wdg/lvy60eiw1Kfi0praCebT/qMn25YJ
OOZT2+NFFne8yB3oOTxbXEKIh/AtsUwu5Bke7ghq0Jy1+eOT2nq2aDLKrg28gE7C747hZHSzMxhW
tOo9ARQaaxV6TCN8pSEIahrLNt/Hm7JcuONS229s3WwYQT4FuFutIXSuy5+pvs0yzyv3gWt7y9k8
1TrYGxJE1v5jCxyHOivRvUnMTod4eBpCDumjqUjG0aY7TdZe7aQFn9NMLEWVglYPM/peONQ+2CpJ
5se4WXYhmqO/9Fuvh4OQRt65CiKEwAoghZcofpVzytMUDSYo4VbM8gydkTrIcMv5KlKN1dU+910Z
yNfGis7jljLTXcoaiIoSbPfHjY9OEsfz9m8miVv1CNuTCPfDRqxRjVFZ3o9D+17glc0PQ25JESTT
tHzhRIcGhMI6vMGY8yPKOFaLFuIpore9ef+PzRq3rRdMVa8OJHS+d7Z5lfZtwcBnM6zUbQnE6lIL
RNWylXNDzfMiKEc8DedPPhSvRK3cKbx00nY/j/iQzki3pv3Upd+RWbtJkbNrF/1jAUNEuQBruzq+
aUX/Ayku7U24pMY5TTMbns9WK4Nqn+/lRzh31cUGq8e6Yb5V7YvMMLfPJEyDoegi3gOmdUPgAxoU
dUqK8apUqyuceYNG66ykIVCQS+zgr2BB1wVJat5dqrysirz+KZzKmvPNgpBpp9gGvlnSpv4awzj9
pbTcBALFOjE+7dK4yscQ1yjMRtISI14Zx/qX3kHVfwc+4HpZQjm0yHmrpZG+bajEOZNxylD96XYD
h57ERp0ymIKOaMyIWoR3g1tmXSJWlhhyJiaODS8eb7nZF1W8VJyrjVSmngoAX+VngGXytGarB97J
oR/xG929/YBMu2JIdMO/1CEqFOlq6oO6xQf2nnBbr3HCSRV9aXcDPTdAGdMSC5NQFWINtodifjy7
nHoEEZ7oHkkdf7xzkpFaz38ztGK3+BGP7zhTTOQSpWVhD4u4z6hxeRUhLkg6O+APF2nIdBRg9svS
82FcjR9eJVoZuBxdyEd7yvzTKoQqqGMwc5VdD1fzbCDbd9zbXOHavkZhuDweNWUVB6KFiLEHWcO1
u/qb5BzTPqTCaxH7SaeY35j28jfYemr8h41BO/z9QKRwR7tbZOSelW6uijSuHLiJ/DRrJlnmURVi
Za0TBvds/dkNnSxfxoRuJ9wM7XsfVLV8MgVAoRFLBfb12zj82JJ5HNOxXiDbTBpPj3OOK/mAxaZu
OqH8CbzHUVZVp6e5Fkn8xkXcNDtV+pKSYCwvrRBN8hbSbxTLU+maIVK/bbvbg/YDY5qZDLOwTrU3
Hq7A3UuD0Suus6fbN4Evlri7JfysFM/TmT7Rp8ckt91GvSFEHfKa9HAfxh63FLPm5Gst5J/6xc6v
QxtZyO4xIZYHILkWBe0UMjZz6zh3cBnyTYv5NqkotHIZ/4/Qpxb1qfdG/cwkqX74pbIEndZxlfvt
zEeR4Q0NvzVz+nXp5GR38u6OCeRB114C35Baez9mwUXHOpb0efHRLuT6f91TzgydyB7vqDNh+m1K
WURtz2rUvPB2vnATOaB1Psc0Ov69V+Y/Zk1aHOrMK557fR3pLBwW4TqzUW6MbELnaPbLoLpQe11y
bJRtnIIlrj9GCSTd5X/2vWhPZ0lhzLjQoWFlKBU/QxVgSBPRgXllZN7SSBT4OgHoEC0RYbrMcTOM
mO3bOJFdardu87kG85kyvsZZsGqSLagpyWNUtztc9FJea+dYisHHNih5FNX1kcCIwmXB7k4UsULV
8X0OFGGpw8vc1rKbzM9bfzkwNVmcj9zfHN2ouSmuaMci45in2Vt4/LckrLtXhToW+GecQXlAl2dJ
RdzMk5u5lrVhI3kby6KjItjv+yTICFcDfixzvEdvq1I9ZdbrG3qrQWIU4S6LbLDJ5HvYrmUYWTiQ
NIg0/ffAZvdM2aBPXMEcXzu0oc4gSyBt4o0RSncqlCDSd7REl+V5x4Xh7oiI8rMlPVLGCRnkV849
IsJecUuOfe/dBq2bmQp5O7HQLhi1QSoMc5dRBGqTrxgWSR4z3BP3YKaFfEUU057UPAbAJChCGoGl
W/RnO88fjH8rgGioRSJiAk4/4/qQ9UhnHd6n++szi/Mw93vtLYY+CtLUOMaWHbprYAfZWq7Szgo4
o8KEBZxquarNjrNFFGUEOiG6BoQx1MbnDDcsc1yNKfpiBH4gMedomdoDR5xjeuj5d8OHi0OFZGsr
3EqR4Se+g62r0C6/tS8V2w/FgUB00TwOhkqltIGy5SW+xR0AW2YkEuapJsG/9XqlOQB54+3fyM4w
sEqrUAvzR9SK9WOLrxHq5N2bwregllCX1GjvmGuRLuz2/F+bJgOpXwyn0XtYLDJGDzQfrXiX6zPx
ERdiF1rf0Z69z58W1MAH1qiRJx2jjtDMZ9TBgQi9PGh62GYbDtbqoWCdaR93ceXepGM/a9n/B8C5
XN6Z8TmYm8AKzgXzDdYKczIMbo5op30oI0QyoJZzQhVdZVYRAKrZHzkzgtT7TcpM2aI+E7+E7rRA
mJQAkZ7YbgIMAGp55CCNNI/bCrRdDiCoQMPJSI25zRxiHeIH0MDRUXqhdsOiNzxo4U1aNHAesBjR
jcjtzuR26RhPAAywLrlgea2KiEH3BjNn5N3mjL0W07XN/2mvOD1zmevc7AkJAYjEzK2wlHCCMplG
Rx2zgpWN/wnxJUNyssu+eMKa3gagH/Jeev1uzBsS9JXxMEeCISRCmgtOOIWsinrK0T9uLdH/A4dr
zoXzmXUtTrf8hQBKssnipcbMc2bXCC0a95I8UU3eysEs17+SG46Rr+ejrcg9MzC869Kb9NkKCnuz
CdYY4Zt2PZ2xH6+j+6/yWhWHQ3lRPwSrOpd8+jEK4BuHICdPtJ/W3u90D0hWkhLGiig/kdBdaIqV
nrf9TRcI0fQaie3SPoEDb7N8maiAImtIHFWcHB+trJ3RTyWbfVdwlkgsqujp6sh6WsHI0XvTIXW0
NOXY6pftez3qWP2kkazu0FIWxULssH4tyUQyb9cqQJUOxK9ptvltKPXPsbSLOpPXaAOTsvaEgkYB
zPmQJlAtDprL42Htusxi8zstffiRMf6ecLCZnjT/t2SQMwgJmKuaJSkQuCR8pcxVPr+hh7iXIl/X
w/TtZpLSvVuP/DogT3aDXntDPcOAKN5kLBUxPVlSVxBEVEcV7tEphidBAOl44DCHfF8pqqs2R6B6
1lOBZq+uI2fbzD0R6T4PP4F7zjM4aQJLJ3dNxq2/qrj34EljGzObd8KZAiCRsxCD2R54KpHUANw+
KzMc7CRs6II23bwJYYJIPaykWF8oBFjCRbUXXWL3egBPIBN3JJiYZ/5GB8GntpCL5yusGHpgVlds
JSsoKKa0tpRcr3ojbaD1cKTjKH0GLuVGGm4e30A5txSoeDI9I2ZA4gaeQivwzr008cG+PnQ0Gs4S
p49/kf9wQppEJvWfoEOkajUrXePl6+7bWXMlSHpmwGses0N44NB2zsfqNwTFRUDxI+kosxmIHPfr
h1r6++e//igTTZMOCaK6trcf67eVA3WE1cbFQtohEojAi/AsOChoQgAJ45pyyepOwWI6T9SNn6+/
vL/olxC8eIGWG81HeuaytJTCtJKd4ys0M2irLHL/oenXMiJuQOwxFDVfv6h+JAKax/hNcPKIMHbQ
lgUNZGfzxwxEJQfQrW3jjB21eiNytHGskuUPv1bOrGqyCZkhrDVAKXPWITbgDfxlNeq7dOmDL16N
JP+OTFfHxlUZ+peJXnawl8JsPrP4vq+RwOh6jaFcI8Z/OFrXeq0ozCQkV2eEx0O/K0U6GaFGyQpR
F6Nu9KaH/2d7Nc5nTBEcgf0rQUL+DOydRG44ZLHxfJ96on7SBj8xA1FI99bqkW2886TWEbtyIPRj
uwWQBA5HsEeZQi+uIYkoofHRpyyEC1zaUBZzoalHZgaAjTDeCakut6QGzbtZtz6vYAGUQwv3rFr0
FnHTXqubh3g0LW4A9VPbeyX/OpJrQkOfQqQ4w1t9Z0RMqsDBkxWZtIFyuLblW5WarLfr2pytCB3o
KgLRdm95uRPXkBtpL6agYld2Vea1KyfPj2rU/7zwAs+nnEgd24dfAHb//2NcZz0zMphE0QVlJkt8
Bt7hl051zm97SbSYAkAITRCPIJjRSDnercaY+G1AhfPh0sHCVMJOnx1JRG+qqXPdnhFctJz0O6Dl
mZ1k5rB0cxO6DMTehnjWU7+mzp7rg3dd1fhgXArfaWg1tTOpriGxRuvjmuQBHW1ljiA6GYnlHZ6i
Ie9xcM1FSc3LdqCwv2jijEqEKKxh9tlq0Klv1huwTXgkwPn35GXwgKDYradL6bnAEhlx7s3euHhR
j/W28Tp81M33MNsjKWbEM6J02/N7+AVSgytitbyTLjeT1weWl+M5g8gC77ASsIEIAqI389iWZxgx
EkqNY4+Ozibv6lMqJ2hig40E3Go1+2+KVdhRengSBX8vPdgBvyxve4z3bJotYyqApkWj7ik9omco
WNMR3Tea9bF0vU3drL5OHJSE6MJqJXJIHX53GwaS1abb7yMI7CklHelGKxaNjIYR4ijthsr1ovtE
+SYc2oaBZH7o0K2BhbcyIbcfjWFQyCeQknbDB18D7c9DvY5T+DEEwppbEEkpgiVd1MGd1gdWlUTY
FqgdZDCM2zitBqEEsmie6KvLjIEUkIqSM4fFjOPlHSIicqxhmyxA5skakeRDuvNH8eHD7Vsfd0YY
0VomfdOiwOMHWaBGBha+mrFwhGxZuVHPYo/eKiCwyhQMH/IkG7pUoWf0iAwmuHSTEjnzc8KoiIq8
qnBpSKJO1M+6BVAeRei2/SDl5mzWqSc+Wvm72YbtiBBButErHgt840/QzUxKZsJ5ZC3BppxxLcbV
iMhvv0iuGqCKro2/Kn0uo++JymTpxcSvKi40Jz3Ttq0CfNR/9Xn9PgZiSeQZeKWwqM+qjoLMtevG
gV6nWc7kD+THj9Dl6q0fOm6/JZJUhHiSuzwia473DN5Aon6dG+TGNQV3OGSqbM63PQMjlPMHo51y
/PLcWfhGqnee8XrSiVgpEbRREz2HSP0cqgO1i3O3G6K83MwRvCciU89U08+Dn4EfDL0pJ8Uq0S9N
JeK+FJrJ6qkH9LOkTXJpU6lJaoHfzVzBEHsorAbMMCnD0Hb5m/4jKVZjevTUdP5e3dROtdf7l9BM
x6elrq7fZmWuDd4ia05v7CsqM7lc5juCzQaX760p15kQkajh6xdtfjMXDjdDHOBKg3kBveT+uzOd
g4Oj+2a4XhZ8rZ7hyh5eR6aj2/muPT6E8WFAYRcaxBo2LRod+AzH8R9hgq6TCQEn9aKFLp1dVAG5
fmr3Qc2MW4KeotYbOxS2U2wLGKGQqpFTnq47GYD+hpxYbGql9S/oDqBfwmFu958r22f5agLTkZWq
nTx40GjfquvwQoVPYiPse993Cd6udfCt8rrdbm/BhR+Syy4D/zFq+euWFU+U5Tks+vk9k0VH6RAQ
emP94408WNJRhfbpnja8PzQMQF+n8aSqyb8is1ZiUB3SVMpd/nsn/l1RCSFQXE+hunqdox+lWIVG
zndMGTJk8X0NAl7ROV7O8VlBYLpIiaG6JkL4y6JSpFlgsXUvrJtpm0X5vvyDpeMWpsf5aPqBIpwK
ybALit5fbrcFq+5SmI+JZl1VdukhvMP/MeLd8gnABBeAeKgL5q0NqE1Vp2E1DO8MoOh33+dcr4dV
pV/nbnSO5Bn3gtHNUF7JE8zkhRKnkn3JUOccP6GpxVqgQiOt2GWRfXBktYcQSGYM3ggGExiyz6l4
3upPC1NkJsGowiWumdpcjKo2k+2Y5yUCFBeCXQ8UM7jRawEZxfpnKfzA6mAa9cFOlrp/5bVgkFPD
9rtK+gXb/H2OfHfInmXUgJyqhR6Mv8iddL4mYge8cP1Y15l43dcaHnuN3h/ktJv1mppt4zvhe+no
oWDvVtZhmNVPd9JQr4D8hzMmDnYOmJaUToCem5marCjvpBU5LuDt/a/H+IsMTDfgZ8Ahaz5yryD2
DWGsYxTwT9g5LL2pl0tUo2pEGmZQwXuRnFl14z3OE8JS8vd6RoZSm1OfxnRT4xdkBjJtnqnwLhGr
YsZgi++c5MTzQvs3yX/TYEbclhSfo8W80G3HeWUPPK+Mo0OCZ36M3hJmstmINlhhiRR44GFOErLa
hYluGMidlXkAYb+MRTuDuENzc27y3NCTjtfkI1oBOxh5QjLBxOEgZs2D5mRTamOQisBULjy74JK/
NvkeT43TxR7C7dquRb/X3ZJUfq5neJJTtDCEJYaDhm8qKIwneJryxKb0ExVFlVEVqtHeIXbAb0z8
OOByMXH41Vf0mwOYqqIdt3jGiypo5+p0CIEZ8kbzjOelQezaDlXKNHDxkv0j7QidJdQw9QqbWdOD
WeZ1Jg7cICOiHdV+iWbu+l6kXr/pHcKOyZs5LoXg3q8OJ7UAccZgilshDrDodvNkOq6slzvUdgN1
n5mv9ru7bbkCAaJto4jlJi12ERJ9TvHkxF/TDBA4JJxg++IFG0Z3k2eIzUxyvxOqbu9PDDKdRBDj
a9Mrj9Fd+VA4O/5x2pajRAm+Aod4A9YRFd7poRGEx1Aq/7exujNVg2N8xsL/CCrjk0hdnjvC/Vi1
D7qrdMZ9M+4bD48yp53yZUwymxG0zvwqMHB7WWA6Pp/41n5V3TJAb5//ZoDOoJxH2pWDfE0QegU+
GLwHv6EpfwUix82QzOHAApsQ74SkO9/wqTc31/BJbADgI1ACXbIic1zAlyRvs3MYGTBOm8WaZNfp
oCi+UJT8dPPDPxAA0BsVX59Vu+oN3lU/MHXVysIxe6+ijoGzRxUD2UTTaC6qwx76cbkWMttC1QXc
pYPgVSDVa09/LkYPigx3k0T/ym/PrbXBAEjw6c78uabKOrkMiHJjvi5jYvitsYMR9Dzx+eTM9+mB
hwamCoEIf23mEU2IgK9a0jIgErao+NlB7x3hwQv3D4NlDJp14FYk9sebSEhy/14s5yKLGxJ4jKaP
mA2F4lZ8l7LLZhQuAx8EUN8sKZCqIi6ATi/7AiTsC5xfVxO0vTUgatZzLaWAw+AWOYOaIo8Wk5fY
LP8UkfTCK1SpErrMmRzYIqAquzULy2rnsdmZ6SoPdxVUk0zO9VJoxOQI7RcOiE53Qm3w5crAnRv1
0cjKPXZZKQ1F++QZQbywYKMs5lsbHvycfwf0HHMCpiaBfiMbP1VI6SErS2i4XpKZKwSOrt0zFAlL
GjEIRL/GO/Koy1h5qJyiwp54mH/NY6h+rSPCdYqcm0VnZ8654X80EsK8vttrD7Y12ZJuEq1aUVUN
Pt4N7iWgXrHVaTTD1fmZvycWM4Jwke3uXh8QtyoUcCGF7og5ql9AVujnj7hyxmZbnIpV2C6bPhmn
yev+ZsvrjZ3TrzhFDWOmsIMe1hD4ep/3re5KJiBuSRjBQOp9WfgE5FhY42783wnk5lAoFgzmIdfj
Gced5Xc6+BXeGoLg1QRvO6EkBc/koGdXB2HJtBj/4FwRLhH3oBuCojSLSc6hTrbnatHXsl9G1rBI
2U5WfDOKUuvVEyZfKLMMkqGZ9XFrsdHaau/W2juYIGzpJz6thwn3jK601gaeIEsfcNHsrnVUKbvV
D8aXf7s5iYo+u6ywZaP/wIFu2zXxoDMQUmWbO5fKjMNJC/G0LDBt6ZoKA96a3QvaP7pPBXC95c/t
L3ByR5R7M4qgG5k/VZIS3cVlsQ2urv//TRfUEJty2+CX4bTydjPAiHFjCW63LuRYvuXNr38w/PnH
JvWpBSvNQHfn6P8Lgb2mv8gUcG2CnDSAq5Yp/0UTGVz4YdMGRnznPwBtf2SNS7rqh+D2hmJlJiBf
FCbcAXu6MAZ0oekwQ0rzIQUaBXPykLVAZb3AZ1PINnO5MExo0rwGY+TNjPq117x2r/UF1+VfM0ia
SOjeYyUr/aSnIj0Kr7SPlrdqWbJkoWX/BYGOGG94wdnMrHlF+qklrJWXrz7NvKmcIAhuriDDmd1D
VCbSpS5NTTEf64d5kp/HPSdaw543YG8uHZ0/tmgA8h2x6A5osAfoFVTAcYvQ+1P91WvL0BcVTmzd
YsP2mBe5NzUT0z4fz1F3agdZBcxsojBTC/VIBGRWIWdowReWOcNLY9mE4OO5viymgCVH2Znuzidd
vpT+UcYk7wOl6YT11bDF/A+KrMMgOUJmU1xTU3osyKL2gj2XhGRlqBGMULRGTrjDWJEWnH7g+/xq
vOo3wBroAVg05LyaSFLOMCQTjw4+hqAHGXaC8atOw10BdfEXAlZUjpLKxeITVAJ5B9EmopE/q/vJ
+kidC2BD5U+u496W9WtDcPofGz2otZPw7yYne4IxOHJd9V0N2QWaFOESrEzXTOtPvn2MxMCphte2
JMDMQQEiOGnV0wa4pVmP17h34HCulpxEBAOrEaFeHGbYEqB00dlcnV0Qhn/AIIuXs5dLlGxJ2g2X
sj5ycxZVL5ndKD4IEz+fX0du+erDjpcRiZIX5T5c3ZiCp0/iVhVM7uTxiJOCmKpNpLZGn9OOn0Gw
3vDSZUn48csQqLk4+PEFdIIc0re/7+RAi26oxgMLqpEOKqvbdUZpqad6/u25dkIoBU3WNTclZepF
l2MI4Dec9RgpuuTaIudTOJUsNNZcuGGAN/K/kF95pF9wFKJsil8H+zmUP7pmwM4wwKKvM1DMIn/J
pygCZt+efy2ICqQstlfJWLIRxm7Uk69bfGsPhQ2m41VxkGbmq923a7UhXRN+813lTphx2qoxlerv
b6S/EL56cjGXO1pGC2Y6LIREjoBp0yzEksmEJSQJW6tVPd15DfVVjixf9QftcPV9DSVNe7SonccX
9S0dr1Om/8ltAFYZMMbtMwRTqj/OvQKq3qGufaSzIQmGcuVHvT/rpXNPh8V7LgNO2rLllMazy4Z8
HnHoMtg0Ea+wdkeT8RxBsIYwst6BKFDpAJOybLLcgw1KpHoafoArbTc7YRZ87b0b+8i+N1rFL53K
q9D9uQVxAB7SFtqXwGI2UzbIwNaOAjc4HhrjtGf123jfJo1t+GkONksSC9WAiGSEi/dszcSWTeV6
ZmCK4+Q1rf6FJZVe+ipQ+KYnXpZcOsvFNpwAjKdWedsQzWQ37s8erNQehA6lyHHeCDyew9AGBlfY
ar+TeAW7rbN7vkx6Z0RFXt3gJ8/EPW79+2zwlWpoHZe+U5TYHtChbgmIwfqLRv9XSxctXUJBczB1
LQ9l4HUPdjBvjjEo2cdy8loy4Vr14oabUlNnZ5jUjlQPJzwb6n50PJPgYho4Np8hKlMfkwmZX2pZ
f+CMx+fVpJ47NVsUVTRDxMykXhV9vtC94tY4yQ6178/s7ybnh42sqPjTGKto/0a8fem8z0QTEmcH
hMaNOZ3cxPazJFTW5qGb9VtBG9umIepoVlrNdYSxULIY9x1e8xJ7UvVMs44rcqZsGuEM4OjVer+A
ghoE0LHcT9+6Q4krSBu48NRdvrfHMVtlM79pelMRqhGP9GLBtRKNsTskf3KRVvVS8m6Zkxpw4NoI
QY0HOEVSqLEFkbRcyoOwK3pKwohPFTJ0NAlZKgXSy9DymamNEVwDAfS798pJfUv8SUEMmnL/dWmj
TYjtjwtcoR5RRrM6M+53SzFPlbCXs6kbQ3mjtXmnxX9n22JeYqMy37FUNxzOWIdLIpNfu/m8SMpZ
Mky7v4gWZlVplpJtNRnYfroLp3o4bEFomhwzJEGG2nuF8tRNv8mh6Oko0h7vEI4TIQ7f7N4NVCzS
RXscrgPzHZoeeul5qtHTPZr6D2y7MwN35WGNEHr98f5ij0WDw8o0CtrNlh1zx9AZ/UmAU7K5SNR1
hesiDc8o8Oc7+5VCc7quyusWwCx+mRKKL/d7MruOAIO5Nns9McwPryNffLFOuMZ429pz8v3hLfE2
sIrzJ+zRxsvmEtRg2GQ03HHi9KTKbEuIo84OY0wRjAlzqL1BYn+XPHnNvmeWjfPFn4nt+HgJeMdM
0W/EjJN+GEezSZ3A8yUwS83SVYkghszXKL3XLC8CgIs+1GXcDggQikkaQRM2i3f7BqETKojNgAu6
UiCB9t8oz6/R7DnUVpMgFI2AFJOzFmK79LkS7O+71FdXM+Q+3kBxFfOPvxTImRm0QRpZ3+aJagw2
2WyhzuQRyDZrIqjLHJV0ePzbs+mi/ogJJJhcYufAQ/rU1trnl6YqrkP3NJ5SjzFJ+M55TidNUWlT
a4cih6Df5UTfDphqJ6lzHGiavrYgwciZJ5l83I09rHXUAhD9NRKOUyEhSW/7Rm5acZA2j2QsCgOO
sA4Oes9tUPb6jubvBqm/gTtzy9dM2SOBBysCvc/CpQ3fs6iCeAb2P0yGwNfz0a5Nsex7mxpUfBXI
OqEoO1V3VVTYMekHWp3Ezx1m62zdCVH9QekLM8G9sK9TfJJNArO7QLzBcAWacidv4kc92FV0ktQH
d/IkSPhVeI0wld02+MXwo1IRPXUt5nehyiF0hulI7SMOdCv55dhOE+yWf+eqETorpBUNDrAgSE9I
0CEwcQMi83tDjNuBeYBCukvhrRY70YNNFv54vwu6MuuDPlE7d9pcqQJWhFxdw9F1+rN1oT23H6gV
kflgD7M01YaJKzeoYMUkjxNAcQr2cGYxzf7QSUhzE0YbOmB6Jk8j6g9nKBDKXZe7X5JFHyuV/mbo
R6v0L6apcrFoAmPvEwb5WUi99c8Ooy4LUakxuWrrnhBU3QOx2jZYJd0iUjMaHEMw6Q7MjM8TiHeh
zcftbKPBAEHZ6crlR0LlZT4nJ/cyObq+iF+nI7qntdspBunfT9o9/Nh4j9o+zDFnl0Js7xAvv7yF
lH6OPWH7BBZQQ+gkZbOxy9lEAXEVjn3ntoAg/ILCU3jzVbl7xyher8NvB8sXdiuoskgJlerY4Kra
tVm8e18AX8xWUGOQOSqTfqRdPdfk6BehNE1J70I/PyD0foicRoPW7ZoxNF1rayCOdoN1bWA4HwEo
iKDkluBVHOjGfbsXg6LYqSdWnfvjPKSeeXlRDEvLhE54ScukcYwfBghM+eKXwSVQQa0C6YEYCr0R
rqunvA8NGtVag9qRB41K/b2ZwQ7yVARAtcRj/k+jTDwphI0fgjG84jB8KFMdqXoSR/Ev4BhHSPiR
H09e3YcIkTm1Mx4sDVVoywyft/wx+nhpzRQ36vOdRRmll4r8coOYA1yJhF0KLeTsIeY2LW0t0M4+
kGpmstLP5hXAjzlJN8V/4ppyluzOpAVZlFNHhlNrVhRmtOwZa/YWShWNadm0Ulh45lOFHQ3UR3O3
mIPfEp55vxFxgBVDlEUZVCYVmLXD0fTXdssCyh/n8migXxk7CzTzC23JSYQtVoOfHxxJ2XSfvBR4
Qnc9XfJiBlxOjOfTIRzN9LYMMTrIQe2vBraXhKAO2egkAmlIs9yV4ZXcf9xCTxtpHoMXNi4XHFLY
GSxrTT34WAD6LeRZw6tZjN3FPzCjvsKTBZnNCySmPc5tCljUKNsjL7jrxRe0fRzWqoHDJmMC5tDo
PU1+/sT59I8L3gghyI0MQQY/tdWxjdWPqrbtA6OYt+syuec/2UCf5SP0uRx9rPglSu/nILe0uwPU
EQOUifLrgkttMYlYWp/+4uhtgYXf7KG332GXKqrlmg25rOsLGEjCXmCQkamp38CiQc5UCCksbGYn
RCUlbrS7JZEMqUnMgKyLuh4NHKYjoY8S04IOemztCzhDTj7nnFMpoSlQknoEEwFwQE5G9UX3N4x8
jWThKQJMwL+Q39LML+/J0/CrgRl1LCgOBVjwr3G8O2b7ktNoF7YRoUTEGOX13i1iGB2Q6+CEoFie
JxOa+Dwo6E9n2TzMXooTyI2shWAhc3AtFJjVphM3eI+7+EAs4oazxIu+LRk5Tw0ZALWvbwwu3Tz+
wDRfjFYCOqrdjZpwJH5vzTNnYS3QoyISaQph/+Zje4jupzsHJhPBomGzEVYTtQqCQXEBMAVjaloi
wP2xzIT/G6fHQqnZ5MNEEvRYdBN16PuCb1p/Zfj75z2cmWP8kedT1ugCuWw0fEDt2P8amdkTnRk1
1mjx2JgZ1bXyDGNMnHa/GDr4bupascdT+0a4o1sYaLSV92zdPmCammavur83PPWSsqvB5LkjTPOK
Mk+Z3iCZYbHcobklWBj6iA1saUySJwZKx27eo4NJFZPRhQthZoH8Lhb2mOcm35f0n2Y7nqUI8Xbx
UDdKnaHNMXNsZC9swPeWU6jg4sf3GeHposSeNCYrm9+SYDbAu9lAUZkhRIc8SzoWfNMdYs8P83XO
GjKayInizvpd3Oir1aEA46vg5zBkAmZGqdNvCzRA148ZA8FsEQAK1AAJdyvAnJEskiaTNy3D2hry
5sZu8vIp+VdelFasOw2zAK+1sE6BTJ2FQXED87Yt1hzL9+WSAZAvG4fBmDJrcDWELfpq7v9aI+cP
bEUs95rOMDCOVGVgE6BaIZPjhL7FFOIsieQp0YNqUrBqSX/iDdE/K6tyic2IMyUaEDfZEb4PllBt
MTPOoKC2mn0OLJp+9ysBMRTGKhuWPoyGj/4/PF/Ae/8m4adQufi+Ex0u8eso7TpDEx0IlxoJQvuA
qlkkJcQO/hVP9hr3dr8TEw+w8Ooc7UvFAWoCumpS1DvFcJ6+oc74yRgoz8KqIf9gJJ1whu7pS5G1
5LWmseF2jT36SMuBniJxEAmsgP09vhqms1ZPZZsNmr5LzUeL7f2WxlRToTK2OdrSz8Lzk2b2vCBJ
dBRJr1Yv3BHyW8gz4iLR1SrLG4AXxJyt7Bpi0W1utDzrpZtPY3Nm/GDzy+pzIjeyaZJFnDw3SU7B
0YnNsDJ5wJcPI/FCESDCA5m+5fMHN49+9gvOZTNptapWSAoa3Vd284+Iebn+MJWmmNA4DzKmP8so
0bov0K2a8Ell/TX0BglEuYEH0jUFiN+Q5qORu1JK6rRhnIXikl6V18vkDbL435iWcPU7Fx5OGXwC
JAUQf9x/YGJ862/Tc9ZdjlbdZEVSFGY0qM6+4vpAoO/b7R6Bver65AgGG9ec+wl/16QilGqiePZe
aN36P9YoorMyeiImEYseq8WbqRvdfOjw2Y8NGXeBgraP6OuU9cLgUrqwFWlrS/xus3JgfRBOnKnc
3VkXzx6nlZ5ae5LD5OMZB0ZfL9uIeCpWg8wmJfgfAH6g39rQJ/JRNFRIE5PZPj2LaUPJK35VY4/i
/dBc/TXXm5hA9ojmM0q8fghgo3zx9LPSwEhy2o8hFMEoHcmxHu5dk9Y5N41XW+aIkdS+kcIlCGTv
deSx5wcVyALJbxH1r0gL9STPVll4BwSGfBCvcDV9so/wUIO/GlJYq/aSmAnD+lvfW+2i6YMpvMDr
PXEm3rq60zhxluupYl4FYitJKHy4d87DzNdeHiRuYNFmsFEyJSboUGD+HZR8Ne5VBpckgy1gS3Vo
1fr/RWlfvASr728jrYjul9B8TdSEBYzr8ddN1hiksgA6kyOzUwhlsUDiyi9rGSF/wu4TpTSGBXcu
5qXuFSNT2Qog6ve+lJeMIjxii4ZXsaKY7LawF5xj55GVgLe4T6WFqw5FxUkh6+w1TtAK7NRnlona
kgp7pEXuKlw6QLUG6uZu9P+P7bSmwoWSZ1Vt8CPr5FnjBLZOnO+NiVkofUerjo28OkmSpNzLVUco
P8b7xA43H/amPxQNONvbJWHvj/eU16ar1K7gqUiRMenYC2lMogGquMGgvMtqeiWa/Qc+/8IHpRHv
z7SyR/P3btLAt3Lt+XML7STrrpwdOL+gD3qGxpM05j7PcKY+G95JheadaEYrl96MtMljXRqoLHfR
9WEK5meqp6jwbJDhqNi8pFRv43O9t0nX6tA0djh5xCVcHbbl8AcHlDJwHsONa2471nc2qnIviMoa
O6NgTl1lxy9niCT4Fuf6zt+5sbNGpkDGgBf8w9aZ4Y+eKag94ifD9Yc19+kLfimw6rVpzAIlWawL
CSJNnBYgF/g9DwJ/Od6nzFWsTsZPMoiLOwSy1OedxKeIuqAqE4NTGtSgSo/pc3Np4DHhpOdWrQX5
xQTxQxF3yc1N45VCx+0z9oZ7RiUz3AP1IgUo9JekeLd2ZLeTeC5cAbzCektlV0VDYXiv1M+Bdv8N
W9gqxNoEISDkmjJN7VmywQmWSLUb590sCFSqRg3M3AqDbBMB74JxDgGFmPM3jMxJY9Zi1blnQD4q
JHFNgwTXvv87G0y14y8r+QAPxLUDQ10Lj9wv3eu1Xp5sCPSE7PqpEZhbsx9AYa9EeP6vQgZGs1Hr
c4RXwgiDBTHgemRbOC9pha7J3gqJ4RxXD0Lx3HmKXXcMOkX2f1kpGpjO4Tep3uSqeq0iIZmXDf66
jeMsz3VqaDhB3nSvDHbGWwmdjpeR/+aM3t1yu20ntFew9A6DuK8o1V9AwvkmReDOLkJOyDYa/Fmn
NCk2w5zkEnjHXag8VX/niJioLYhGfc7w5Zj8HdEzxpw9U9Em4SWR3pg8VUY8NuEgcC9SPCfZnGmD
T60pqvNrt94TnSjxhXX5hzFsMPo164MBNJJirahxFkDhYCxqahpIg9iiRzav5UXbHQbfUeFjpuhX
OECDnQcHH8tAIr4oSBtpHnFJ4RSpDEyihwDv7zEdcHWVkbaGJFEHo/t1UGILRZUXaoYF79pKu0l1
Nu7ZYWUaaEyfw6bhArlCB+0eN1ruFWl7yg8bWjiInkQ7HE2UpVAb/jzucsgxsMohlQPbbI1ARvui
kiMXBbBplqDVHy29wrLhL5jXKK0acDrRHEctXGBOq5APRmvvG4UQH+LKnJ+CCPSfIHBsdADUeVOX
h1DA4IS9hzp8bWFrRzDh+PyZpbFuKuDd1IGNmmKJeTyyZ5Z0rT4K6ldXqPZe4rAU6mJ5GVQi0Urs
GHiz57XKoynxmX5fYigDzg0/gJSaEi78MJo9dgm3ciDGLlTLMES1bUfxq0XsgVpUTaQ18m9/TZet
wUNIxd0MjqzhAKsAf3Ak1A2D0//n3G/0/BziMxOvoJ3TQafgBaNnc962lt/hRKVAWZdtFwVxp2F5
X6dlX+Xo2CNNnJMEmPu1KhbOSgYETwM2QwM+Nf+GkR5Nx2AiHHdM/h31KdFqwhc/MK1ALvw69YBT
0u1PqIr13o6WFc6mRpmfDAN27LwgW+0Fq3Qq7q1XFOlQRtTTvzz9SkjuKHTy1HLcJWspFBpdW4IN
jVw/HBSQBg9Bfr84mqPyAf1F+mPqtyeMsQCsEhKOYnTe3kYnyGU3jOEovZ7IL7F3GnAjNl0wWvKj
zjZnQu9LtCjykJVYcN22sMXn0IjqehlEKPuPsgxvf26KXh8fuBFJQRHHbF6NGT3JpS1PoooF9Z6n
B3rqnHGMZu1dfTFdJIfFfN10jdd/rVsPBLDYXyC7aPZy9Q8zNccSTQrRGQJipGFcNCarWYyWLi+K
vsKq5aEAIK6rdHlVStcis+Y7xSqI8na4N9voZl/A9val1kddtZGKl7swsfX2PUtUkRxg4i1MtkCn
2CM4M4WOtfq1ZONHTKyZRbG/spW8TKZLfFdq6IkIzjuV2N/IFhiKBuAd6Haax6EtIDn5w/NAa9DK
uCMusOgo1Dv4dsSgk8/76UOnmnDyZNAFENiRwDh3rkWfSe/TrMOJ6JQ8B8r9CtGmTz496Lv305e4
O4d0VZBC0eTxo33+o0jny6KcNq+S0clb7utAlyQWbULTjWZLQxkQHNqGIq73TesH/1ENnnvsFALU
bE4rLhka7mj0aUzF6dde35y/UKBVqRWIuDvuFuc11TAPFOYDo+yu38tY1IXkuwSgmZSAjG75nPMW
ooEokQtv4GIedb4uk8MldVmBL29rOF7izGUNiYQLhu3tzjdLEj0i3cwukqB9vVzQf9EGeO8Q0wkM
DHeYkVjKZ+4TIalATg49p+UYNgQc1g+NJeODcfOpIhx5yYvF8hfJR06P/790VvWNuIL9Qw6Kn9Rg
fdlwmuj5jFekOiFzzZxz2Dz3TJ621xrAtGctv05zuwkDpnmmkTlaX5gujAM5pSZENxapLxTI6a2I
oSE3AzRu+Mk58hrRN4J7VYSsf8/NthsK3iv30wyXPSktP8X/qup3ME9E7NWmcfaGr8g8qpR8Tk3Z
5ut8nY9susRQr16NwHvbkk3NsIJPsRmICnDuAsSM2dacalhZ5qIpa8g1yWgWaeXG9WxeAqIKBn68
Ik6HbdmrFpSW2wVq5x8R7nPGqwDwl5/ELPI/AC1I3zoTLGWweSfB8O8Iq+LJCgGm7do94R489XGA
dw7fLPyJqzEiKXAbNQg+elqUt+PNx/17JnXz9AVE9qc/UNXMzu7GsEk7sqpiL1WV/Uktt66p4bgw
oCtMUf8stgy8rtJcTnj/bddUfmNE9TUqaYLnvOdTI2QWvHR6iDsDNj8Z5r2zBiMJt/E7ARoswVq5
j47KhaM3nVwiHTpyr5fD+ahmBwbEQReE5WnG2nGo7jKjMA0BVIeU4Ke+ZQ7UjH6DIwZSpMxC9TFx
3eU/mbAJPAq3pdDq5KFYjkMLovIsY1sOLwA6l72S/gDtKTLMFtU3LpBbGoLN3fPlO4+rxqfDVApD
Qigq9cTxPHHQuR+GA9mPlZVH6pT/vZ5JXq0E5q0/qgJwGDEcZ1DbjuHrizxnHUeawEINAfqyj68L
5VyQaMUDaGxW0Wq0GOZ4IklG0UnzIjHzSz7ZDoqz+mgtwNktfqQH2KIzh38SHY6AdcAn4JJXF2SL
iHQLksoAxfPsM/hYUQYaxs5mgHY26lFbcpmei9hLDQIEej5FAskE1Rp6W1pNu1U6zrL00YOsFthB
DEGt/P8QHs9aFeXbEPrOBvY8U3Ob7bH85bM3YUy3ofOV65CulGNHx0tXW37TzEiLX7CN7AXTKGq9
+pL9OlbBDlCpKEPKq+puwKoEAJWAU63gSanDVAGGDzxjiJy2rgmot8k4RHiFzbCHDEHm9Xvwz/O3
Bx20G/Mw0YbGYKJXAe+duNq+8pip2dmHeS9ssJXngb/vqVkuvS1JieuosyCW6UriBXAbnJAGaWAq
Oe/P9t8SQ96YcTwNRVODdDLVfhEuvR6pfKZbRs7iZbY2mikoBathd7khxToX5ySysEmIPlxj4Vgz
0gcDsgdrqIj8pC9lM9htOCJ1c/VjPpXYCkjjdTqKUsQvlabVD8qPpVQptgff11X7/KTG4zZyDHkt
/bE4LuEnw77a3UkoLNiL3q7m6cYv4VX6AmXcZ2MvHhHXAoRoKkaBOuQkL7WkFIqAFrZ1LsjIo8Ap
XG/BvFVV2q443Lm/npox8lI6pLk9ScWXf3WEV2RytyoTNawn23EqTgXUaT0UnzzvHxYJnVtLy1En
p6wRaZjtLNq2Ep984hVticDX7rD0J2RuVqg+4+W5XbAy13VA5PAYC8wrf+onBthnT3RSOSXdUS3h
u9jX/Lv79xGMiOkT5YzbzciFX16/rXT3Kd9vfJ5m08qgEwmQdF5TjA14vvQ/ZCShM7uHrdTXO/Tg
/0h5o2ScsZ5vmDgwCDke4ZkPViAudU1dyCU3mtYhg57TG2BwYyLItC51uBKSKSavY2uIeSyWtafn
oVUrPnTr0Xq6nQltqsQemrDZ/Z32vNQzuiSH8t8haifxdRzPxAgDhnpC70x58jxAbZs32WKwT/jY
DcFHjNCyR1EKyAeBMhd3VeMzSEk45DdEaagXQwrVW5fsQfXv5SEuxK497LMfq1yDKkPBuLAfRWZg
i9Sv6OsziZfCuESJFdQeHWtIXaJ80U/soEQz/H9BQ9ZAW2cdcUP5XGvL9KScvoiNWBaAf+9qaXiA
Pk6gCbMRYzjN2PP6n5R4KM6fNyVPfoiLguQBkugGHvm7v5eUGT35YMkJU69NE3Z2dOUltwFtY1AM
WDvsWuuQFD5+rlDqWg4VwUBtAOEe3NdN5TtroS8keSNizprg4wnZB7Qha0a0ttikK0OuMCVe4pKl
kHg1AcZpTw/tR0r4bA8QkVD0rHN7SovF23Cye7vkhdkxuwJZgTEEaJSmvNk6BN2aUx71xoSkvruQ
D/hV7I18Wp4wOABw1+5e4hRS5VDgcCIrROEj/DFJZ+1LV0K8LUUMnnyKCZ/PM5VX/dOggJH4jwun
jj5gS5a/CVVNrjmEFmZrb0qwRn5Mr4H2AyTavuOL30BKquf/NlWPPyR/Kws7Qy1YZEntyrnw2Tvm
V0lwbx7to/Asyd1ELbZFFW0JrxGxNKrDZYgUNNVaEuuvvnnmVOGE84vGzF5FBjWqdIDGPjX5K7OS
WC1cpVQlZoa5J21opAiK7e9IB+bxbmtOVmBI7FxDmJw+G0EPt+PCtZO0hmmQ8owxKDrMFyRM4LpX
T1oQ9/my8jLR7FT5xHMKkgww23pLt7wULIT1ABqqJ6OmbmivKssB+0SYADdd1smtPemc+BrMnmxy
scA0k6XbgT4KNNGxcdHlxI3s/avkBwu62+qk/bIm+isWX7EeyCC5HXPjQ431Uo4IOPJiRQSXZsCa
wHvk+EGqP/3Dw8GncS+yYwZSC9I6SShveU46UWs+C4pKQox1qBJRYTc0yFXTDbP0Mg4lI3mXff7v
Lb39eyrnR5VYWCzQiCJIQ6IlYOlw5aEF0jeccI6DqI7NQ8JMGSD8nwX0br0phH2Na09P/L8Q1EuT
gSfu85/ZEMTwOuQhL4SR6/GOX/wb/gbHd+kIAy3bxFbHFmP39uNJv+U1IrHBXi77eVxQKhwpUk7h
AfoGsrdwX52noIrmTgYrii1gTD0FIyyoyp3OdXrDM5RL9Tw1tV0AKcapofb85lwyKxbE57leO3tm
6W4Jl5x2rVzZcPC5+2+8kg/8UJ3cCdSPRHPJmL8uGtYjIYYqzXZXSZBeN7mXPaw0vtD3gUwvyRaO
4qSrb8e+H53thfSsA2Urjbv1GZpLMbzD+qMrChbBB8S5by4GFGrh/M3/5HZTNZG58vDgTgjS7enz
vVkL5MTZbRlJQMa4G7HCZCo5/Bcmsb48etAxKUPNwnAqm15TKIs16CybH7KLIjwS2MTxbPeipOCi
EERBos9lS1X76ND5290FD2A2B4oDJFJxXr+ARIU2lMaWg/GCXqT6k9Q/5vsjc0BQXawRxgxo1tfz
YkhOGhdoVObQvBEq9/2Qls4XGRrrqwsgafIyg6YTO5DUCEolW7+CZnMlrj8dwnz29r5QM0G2uJ96
rGmyOGfFpSNXW/3wxKxkH6FMWDTFFxkR/+K2er2dXuZplZPyRjYnGmp4DdFE8OAHWyU5p1fYcaGs
dchlFpIkUArn6P9vaQVUsEcjG3A3hZmBqt16CArj7Ec9qXvgiWuCUbWqHdxsIheeCiPDh2MeC7en
5w8abyZBjj6+MtHCcDiq0X6W1i4Ah50WbVmGHwtvWOVMCWzUWuv9o39E7WOWweD2nJ32aiWX7UyE
ETdKSjZ98fudEf2WQrhmOpSF2HibYXOHb80Xs/TkKhvGFBbWCouTQvJpEbuttHlOVqm+YrlTK8q1
PyRvA+njey67Fn6QYPM0dWGgfa88sIV1SmVBOP0+xsM2FX/j8rfjV6NLXdJQZ5bULk4SY9wCYPXK
9cOf4lbnHIs2vOiUCd0Kq3tEPf5lGgmufpwiffIZGMGu/BX8kvRHvaTF9uTtG2SWflK1dsAfrev3
khK2lUI80sOOsE8ZwfaAkX5nfp/JaI49frjeVpAS2v4Qd0gEa+Rfd3j/TwKvyJ6sCz/hN1vvEjcg
BQDyGXfGJvyTbxkBuZgqPLOpsbcAG1LwkDNVnWcGsZYLRKTVv/drVV40mv/O9/WnjQQRPXok9vyw
c+FwpRSza07zDztVEElSw2HjorShdN83lXvI0VHAh4ijyTKgTq5qq+QZeUCS2sjYFIWLicc4kJFt
FM/6LxjfmAzN2CbHbmPzP94yGB6Bhe8WC6T/o9zw3fynASxv+aiemP/XELD5TNxG5GRP8WQ7jMeg
iDZLts3xFh8LRBaWHhlzP/dH+7khAPRAgcALlU/ds9Xufz0bdeb8KbeNUSEfRYzdqjGD7hezIeTD
vdt9QlKcj5cclkTvnAAG9CMZ8ckKn1ousnRT6VLoWp7HIerL1DuVqZkN4/kGDZJBPHabliUY/dYm
tSVKHU9qGiRtnYrx0vVCVxfM4IMg8+ubPR1NJLD/4X9PzPMfELj8mso38mq7oqd8b9UjgY5UWE76
uf4pAP7nSDYytC6mb0POf1WiHVWrO7iAdZGDRX63K2nXz2/bgP4N+/gR4GtrDRNqfFDXw0ZpovLJ
k+5PWkzG8NSqQIkOmS/nhCcuL3C+MZFHeMb5XHJ3sNfx4gK8jnM1Z2y7kr2fRUsCiy8y4bdbyEdn
Cu8mayXBVd1c/A86T/RUPbNfs3SGusMQKSV6+tGD5+HVxoPSbyw6KVxbaMsfQ4zqPN8pFOXVDpAF
+mdoLo7ez434gRlYfqlOZho6Uh9BC3AHIZkop0iQ2UFFRVuL1uCJKS1+CYuPRmIEA93ky15FK9zJ
H5+l9lxro0kXr/l3fkaKYgvIARAQanzF2+mwAuJSleuQjf3Evtm1BKYUaaKEJZAVc9OkEF7jkDV2
+CY84s19fkWp78a5pqG6OftJpiPvwHX2HDnl8xQkV6bsubNeszyfUVqVajpPgr2ZTpPA1qc77CoQ
GjHAicH6Kb/emmhocGj6R914VRF+qI46vQOW3xVmQuiMmrKs3jqn/uZJEDcRAMoxVYS8D8pwPNKR
3NgECRG494KhbT2eKB+wCd/JNVqVj8sztFTdFMEW4bf9lQ2L6hJ9NFvTP3FW7rl2yHimhoy5/uY0
4mYjAo4tALEFtyBQ2bStFq/phtM3QNOdD8ih4NbHdIVzwJmEZpy695RbcIxnTt/W7qig9g0dOaOx
KGGhZJvd+wiStaoTon/qEn83sacBRN/Rls+IpHSnal33K7earfMArSav4M5N+fm+8YjeoDfBt2BH
reKeL3BkX1XXmHVLgmedsJPImYuBuxPuIXiM/b9ktMu9pBbLiO1Uj0vKndCZtlMDYyxfxy6hh6RP
vTQT3DUShPwvRwn8WE4HZ7CWFh/mcShw3RtrYR84itri+flitgRBtk0YrJ4bVgIJReiouX0uYJcr
FV+L//P3OmGiWm51M5pTA9+BVww39wOXF0NBHp1A8strfPEL1IZwpmah4nMtPb9LiVcNG+C39PcD
uA/Xj3suYaMKIdPQLQO1jDTT1k07jafiQHDjuch/c6FOZMjRnSi3uAzr1VB1ueCAyBza5nU1Rmv9
mtG5WbJqHuS3QwA5B1cAMUye/qF2H9J2Y6PGFKAQc5RijBS04/n1fD07GkTx9DX9H/fFIMAD/vfk
sEowH3rkGqjmky78rlux41Du3yHwdt0U0icAlPAB/b0VwIZyXa3iQnNhzggTsLo+8EsxZb3odMnq
uRnXSl2SNIVzTZsz4FHCap74lJKpRivhnztpx3R5Sa9rnjs5I7h8dlG6WRsKzMlV6f9S5sJBM9sS
zmfRfMDyd47eh7QQUQCt5T4JDKW8QY+5SlnloGby76S48b+t1EUEEDcs2NftgzFo673m8jE6YiIz
dC1NcC3qICjCPl929PSXcBmDfe5ICR1GeRhGy/OpMWSaK8CzyFCQ75+Xk6Wu4Pyojx/9p+24e1zv
OHJVnEB02RnguLkmqmQ7HqRl4EkdH6fgMkHoJqYS60O1soeHSPJIaDLlWKi2daFE6oDPadmXoZbf
PTTM8BUtoH81l32Wm/3dw2jFuhPoVgfmU1uwHv41TEYY2nVwmLR4/Te/WTqYDoL6kRK/s+ZSSzNk
YsFnvL1109GlZNueFj92iyubCHYZXBxmkI8O+22A6XuqcCGSi5Cj4UYnBCel1a91dbmdRogwfNOp
2UklyYjdE5xf8Lp2qRxE2h33fe7EHvsjqBTZzSj0npFdej7qGa/GP0sSlQduRtB5aDWZdigQ55FN
qHNbrmn7m/KlK3nsJC6IabP9PCLId+MrBQEa/VSMdfVMCHLKJ8D4uG0IR19WvAHzbYSVbf0LXiNm
N+SVEgLV0ZMfN/sKqwb+4yTKus59mCP5RsnTqd7FIWErHZyyuq3uFof8fCFTq00BPjy3u4RuShAX
ftQrPv5aH8mmpZe2MXAKo4wLCrWxn+oxlDDTCn3jfWmniDqqUiqd009etgLXxHOLVHzBBZdGrh46
l/upmrHBqNDhC1haZM85a7oMHlHjkqvAgWqFRJGBtLaf4iiHVsNP4uCqI/n01xlxDzuQ2RvmW4QV
IHj6HnBgSCxa1dkBCgM2nc1Dqtk/5Is3dzp5Zy7jnpu3um/6mirw4q38z+IIBuO8URTznQ72PYaX
8iZAKFcFZbT6fRDwpgg+pxnO0e+Vmg6gQqLoes/GipNZLXO5OcatjpBEWBkMmWyTosW5gePT0dEN
KSSPgth6o4s3v5Z02/L/JL9N9j5au9gvXZzZS5y7w8R/87NiF8i5IlnyiIfz/r786NLoj8l3mHvo
r3++wlb0nfj/tUpn7IYKaaMB+jWLuKfidY25W00Cjb4vsN0bAnvgQE+7AlLMSOqtFSDjx+c99jPl
EEDBrgEi88+ewyhhvEpVTzxKimHwaCnaEADoWCAUugMX25qz6yn1r2VwGlDZGpu0sFLlC0OucdPx
rWHjS47u5y6W9R07GWTSunTsa+9vuaYuj3bD6Dowh8iD5PiTB9Vn6GcXf9vnJc1nUDc1l4GdnnW0
xcI11syqZxJjy9/WxLXCPFEkClzgrmxeKtlUkBTB6m1tH71ufJ8GLDGrsxoX4FGWvMZ9oJK1/FBr
5YgRqyLnpV6LES6YSVG4B8UF5LOmFn+iU5px7UhdFgQgvUSW6hI3UlqcWKjEjMGDRRtLFXj9l2dQ
gHaxxdSTFJtXYXwhVd1uURNpVpXog4eW74U9xtuc7WXUNvrQNfOkZwnRrx0P8JhDGeMeLm8BNl/k
GqlSxZ8HkqwmeESeDv+nafohKAfsHUIObM7ACEHx3+gYzrVZb/seEgD4UYr2hhy5qDfbirT9l9bD
GH98DGZCXmULqDWdmtNSj3s6+xBb3iebn6KvkX/QWt+pQkGWMuFmyoSWEtBdCG3fT9VoMuPeDiur
hB8RrEfz1gXS0eU3WrmZe14qPScs54xgaZyH1bpbLQ+T79KSUqqup7oYPK0h0utXl1OZPlRVeyMT
qyVJYwvFZ3BCRal18Pe1u8A0f8tZ3P2gsh9TYUFnSMvOXitcqLLY2qSk7CJbX1dDutiJ0Kx5C5qm
x8V8JIwtA95mW3c6SN8GyohqMcazgGVTvOJpj65lWvNJrKOYyrO2x5PA8gU8QImlY1kqOf5rYjkv
woW5J1aaETfT0WF8str+gx3I1GMMPUIMOm5gOlpPfrVWiOolfPaz4nwEFSWhcXBfEJmQiUjOCCBu
6F9fKpS2lR/mBLgHiSDsiJQXO9Li+QYHtwAi2TP9EEmnjWryWBR1bL5i8BbkNxYnro+8Hsw6IPPt
mxV8ZyIjt0gtevxGsl68VLzSRtEEZNDS8J2JlL1cZuBCwg9JG12Gv54g/rzlPN0RogQ0gHyjj0py
rbA6Uw/Jst+iZy6jskdJmQqVxwyNLnzt7XKGaa+oCCdf/pmNQvqYMp33CyDkjBnX2B6KMX+A2pMc
wBIOqkV/L/rRMd8o7Yy9+15Gfy6FHQSMGm8gs5agtBEf+/KtUgfq7JTz/g6PpZQTN5T2T33thAnv
IjCg2hJ22Ud0TrbNr2KjxZjFw7sjXTPGBe2xpwJeLwjYFEIxX3HXCygqonPhfzI9TurULVthm7yD
Og5wozj4cb2c4RJEVen9jsUmm6T6m3Daxoe6/vP3+EufcM87ggn8AFchcV926Cr7madtErHNVZHn
MYvqdmBGmpcO/Gvju2jeduSgyLJOl22JbTt6BQe4kMWCRajfciywz0gr1SnymkfN79ferhmGVeYW
Khz7Z0lHjqVnM0lHRg3B05nwTnTrMl0lxD8QFj5T3RXhd5vQEaq0yKmZSxhiluwGIsqy0eNFWz8D
R51Vrkm9DUCZo3O+QlVwzNjyIEN4y7Nxw4SxOfend6Pdn9D3UOucTNimBsfO+PsJ5hMVgjJzSmd3
v4HdxOeB/yKI6A2cUnP/CfbMbAMztKizH9SkbcwPvxTpcm4lNXtfIF+nNUDPIPXqD4Xsi2xPohcS
EL8ANGibJFdkHQv7oF/C5a3ubpEcXs/Kw1RV9f+Az4d2g1bgmcAqFaPE1DUtbuqrkgijMhIzw4co
qj2XvP6kKXSryn/5wSY/RqMpLsx/3zsr7LuWlgGSImF0wUTq72iJx5ZdffN+yazywc8v1xAxrOZD
4EgvW1yX8UGpnAfG0LYXgdIsP+3uVK6N9UaeDNePP8eDRzRiqp3oySKagHutjfhVGCQF45Jou4ks
IN8SYXChL/vscQgp+HhUX3q8DTZmctZdh8mUngUG2+ng2F+xetqthBMQd3ohN0RXJPOhloCoWIu9
weju+90x7Xmscg3lYluw02oNmLckwVNH9ylkVUOVjn5Z/gsiwK4ztRkMF5PvQmgJn20AWof1DaZR
Q64O8Kr7+E5KaUDQC2ZIaHm1RDOX+Jc6kYqr6MCdaHZU7f29xBVqpEpvkZFFqnT7+W1ayN/qh0lc
5bZZXkkaWyl51rGw6tpfROaZR/KDQ701+uu0UefW31ilGoUI1DPt9lyMzjBfMwGdaH9DBHyc7V6d
tS1Pz1W91KITclDlbMXFYdnNXuPAOjJo5K9A/5FdntpNmEa42LURYcKqyHNI2XgYqJIaPA+/h+1D
W1j8QEUrw+XHMZedvaxfjAE8sjfitQhqkQktNPQF75qlpowoe9ivMSCfQNCTTmT5IgeYgMjiqQls
KotRQ+R/0yN5xfbt49Y5vdth8vTwxMd75Y/lPjAKxoIoHA2B8SJCMwPv5iUc0fhDqghZ3iMaeQxP
X0kCgnt9USSBlU5seoFDW7bmK+f3+LrCuMfgs37HpwA/+r0+b1wWphi2bwrVSlVeKMGbjf2SbFOB
0/qjrglyW/E3J3k8FykEAjq0HDosayZABK2vo/A/xuNCtD47GeGEXW3qlQ8as31E3fI9KU5uinxA
i4rL8fU8mANucQ3rK8WAzeojQ09nC9SsEbdvASTXlUFEizZKwmt0WBvczHCU2o/3dVmMAbtc5xZF
GyIpBR1AAFC0lDMPhTN1KsRCH/1Hpf6SYkfSJJJUS6602on5MKEISGhIwFg7gnxw+k+yEvRv/t5g
YltTBenaadLeZ6Kzo36FGDbOcOqzvMRoBJqXywiKq26K569R6kAM+kiJJuYZ5wTclUudmptNSGaW
eFd+PQtO1fASTxn5FJuS6UxdXu7fkw75XhZFpXIOF+NyunR/CWWaw9uy26/amhuWHJPV0QniHiuj
eTn3r4QHLTib5gQNf53ta7jLT3fiK5bJRriNAn/jZbOyal/IMxvCsEZPWCzf/q0qRaKOt7hAC3Ws
YoFIe1oa8Y1VoGCs2QOgpjxHrd0DmRVwMfWM5tVdnkRnnjA9ZMKNGneiAqIiXZAYem7PDYKe3Ps3
XxFRGqfMplHQ58ER7ikOuuqjQJbLLVYUyG9Z0+xNiY8svOdkluwqHMKMmdisU4glwONQqKyfWexP
nhdVAG3PrWFApaAe+vb7aeO9JD/i0zt+jX98wBpw1SuftGe7n6Ci33CmjQcELI8By+je6GLzhK9v
bL9h1zoP1oXp62L5+v/vi3KmK45EvDY35rAsV3g9y+FmWbF1kvo/pFMyj/E3yMacrtaxU2C04TsB
uwMiEHKGej6wLt0EYeZPKxSeuKsZVwawb8SScDEo+uj0TcJ14lweA+9Nz8vP8xk862+qIFrgt3aI
2f6DCH3VnJBG0TZJFBgMZjgRTgwIpFxVCc/PheIQmWP0bu6y6sxx5wLR04MIJ8hyRFUnNh8cUoKB
JLtvLiuZqL/YpOpTzuttQvJwqUVKIxyEGr5B0tLgZivTQjiRpAw5tuwl65GbNkoTYXmyw8gP9uhW
rGCzKYijONGkHMSjqBrj7cgdJ8bfOMAqUyyKo6WENK5FS1wlYSFJKyGHo9NbaXEJQxdlGQLLLM4a
VPQR8JWNUJpceGfe8zdZavmd0C2yjnaxHKxeOsenUpvVavUc3NOqC9s92O+b/DVPi42yspJ043DU
f2kjuIMEujMIcHi9qi3esoI/eTpypDP2UkNdfhYItx+O9Xer04oRPpTtoR/DK5/KTMe97XHStTjR
Vok8omGm5D0DJFoxl6AHMq3aUe5JWXNJMI5w1qSKhYvIrcoMWeS9UBT4iMqfuCYyM8X/g48nvs0v
Qwk63TDsryToaxCtz1euTGqjRtLI6IJSY4S7jarKBVL9z269f1+0pR27aud3wLSgYlmS7fW6J9Wi
BPIxOvthN4E8+r4wCVH4EhmJVKS2M1mRnYBcyyOiPZtTLHp7WLJHQciqYOp/ABB+QULhE8t7WAPi
mOFuCTGbx33X6X3LJXhRGp49rfElhKEoPCHQtQSO4E+qI3Gi4hV8zwhkvuaPuUDTxHuLo5AU29CT
acmO8HBmWlPJ7FvpKW7fKgnI73OHqRYybT+hDWgpg0Dkr9TSMrrHnZyk71qvumWUAQfPajpiMLUp
Xff2AkWlAlqBEEMMz4/EuIK3R0G7W1QG0IYrM5D4wvxjMyJXNKoc30Q7A3vpKgiTJyxeuETwmRPk
1KRI20yBqtVM7oRQ1+XNEgfnkOO+/5vPjpQgaVESO/guOOGme+w9YMmJMhlIkxOBa9tDkquvOMRt
JPReqxKLVY210B4m7mvdKuZSmjJ94A7/SfSEtXxYFegOECWoQPukzRFWrKbgpWl9poeCa0v/Laf8
bf3462uPsKpsdKwYT1q5kfMQCmksIgl/4aESHVxZLl/40eHnOLNmjBwlAN8pqiZhUyE5Jr0BN30C
8EcJ2JKflSKdKRdy63x5ME9/zQU/Vk7w4ql5mqi2Z+110P8kmjlI2sgQ4CgqlMerWX4PILv0ZVWY
dUCLYutvrUNcqwUKTNgUPXMGzgWz71+0Sh5nJJxg8WHutrBIq4BGJdijVbT6uKlTbealJaMzfyU/
4sMxvSGLpnQ2Z42cwQsrMHWr7RU5wc22WcGb/ygcs3IuJx/Cmz6G6RXSCv5I/TD0bOmZ6wNDpofJ
Tc9ztlLRvQLexa+mBCgm2cpq4t8HCTFDg0O5UKKWyC5xQEDr134pjTvl2dbuS0Ws02ERV5rDG+Cw
PjJ0sJ3Vq4d0RQ5DBAgd7lqXYPA4q8xhMbi5bYjepYHRyWUPS5Sjqw7PyxKzOk/AUbtsTz463B4K
qMTLq7ygjj0BY2MAlXvHzS4n+BoFgsotq1KuZK9xoNiIqWzm7ywJ5JDYU5ZJ2JcKdKjT597U6Jdc
7qbQTI82sda+tHBCJTCXk8nhypN+HcjFphdM0Pnx35E7kVkwjthTUwoRhvTrgtb+quO328QY4Gat
gNl/HYkTPBrCB7+bB6vxKErSVFc1eIhFFV8hjQsncIdzx8K5+cU+OMKTQx9CiF0OMwGGS060G2/G
YSK8Yt2MB3ZeFVuh5H6NC4WJ+3krZRlXg6ECrvM0hBYI6keTStcT0XEou4h6K60UkAXnRsv2cGV2
txv1WOOezkF73bebvy8XZzU3ernTNfR9ENOR+LVUkC4VOCWXAXvxM+jYlWL2wUaRuk11f9XX+aBs
H4d5Il417hOdk0yahpF2dXkhTWodjqH0a902nfFs880aVq6NzlsPQAbcs1SfDSrnxw7C3K3RBLQM
QrllYFfKUWHfRtDiCC4qhFD58gxvhIgtUqOV6bdQWnFreWkNtiY9zPqOwxKtDy6Kn+M78lQhFNbR
RrGqMrl6JQzwTSOjFg4dNQuWEX0RCyBeR31ZBdPW8eyvfQdbX2corp8aCFQ6WjGhXKCnR5/komzW
ShF96P5uM7nHtbvVp7jEIcXz4iRx5tGObzR+dNWeRLfzZwxLklvHWPzM/2mURRD53uFuQPcJmvx7
yNkBTjMd0yaAcbbw7AkVEL74A1982Y+1wwPUI1ZYf8N9KkjJ5jF8NpT4z+eAqo4bCocpYlOnns9A
GovxzvI6FBEeYM0/1tlGp3bejLaDvYxnPpbJyeAlJTR6UwqlGXejpFOgSgXFDBrpsNiRyuaBCJpP
ZdN+2RGK8SLz6jWe/1ayH4uvAzHYw5YT3yKKFSi8/VP5whxeuQTdzx/we9iF/3ruHeTFXbLMcE7n
hN0l0+Buj/nRsrp8ntFmyFRUrJzjaK5XWvB47Zg9//elXibmhoYs2nOcOhTzqDFqpdyU4bpXboNp
hb/OHlni4N/37jYsB6seAkUu1qz0JxICoJum5p6h2v9kpjevSPY/5Ztxe59WybG0PmA9CJbFkpDY
qPI+mjWKUjmlGKeMYOML7RPofk05CS8YuPltWXGE4dccPBT4icvthmn9JNt61iQyHnDBFi8HcaxP
ST+XG2KtoLGwrDAi0xt7zZhrM2sphpQ30PY/QxYGR7hjh6dRXYyZr+GQCTRN4D7J8WY9II59YqEU
W7V41Qi0yzu9tqpj21XPsFf5mBKYEaBDhTDa1Nc4x8RW8Qk9XJbZk+cXrgX75s+eZaeLmmag7ema
D1GjbsBbLwusPzPf7d4ASp5S+iSOjlINMJccnWycFb4Cox+4aTxPv5BwwIHniZZQEj/5I7uMXQJd
c+pHNrK86bXRd+hyhsH8rEpfeafDETu2/54n30SfX+KwfKZnqrZwGNxB/7BcxbiMXuJiT1FevJwh
/b/JoQc26h4EH6GZQKtyJ/FjO1Hr00QwvTJ5b26v7XrgBnkSMcgbVjbiwt2Zeub8IKik89wX3+C/
E7KUYOkLlhnwUFmRdMcyeraTkqmhjPohWqBvjTaWkg4bgPL07juBGz0ojXgJ+6uAci4ixVRBOLsT
Z1GsuYTrI+nrx7Ccq6QSGwyNemOSkkPsS4SZUVJKRwMjjvkz78BYH7IBkQ6WGioTq4u/LBKfmCeV
iXNAlLwglH5NjFUOCuA+KvkbIduQ+QUbNagXRfFH9ZWggEFmfy3JnSb0IQ/RgVGLqBMCobC/u9OH
TV67tGs+p2pJ3hnIcVVJfT6gxpnBC5YlZbRH2NYefChuKigQy1sKdhOV9ZN8vHw5ELtl7UlFL1AX
i8D03C1EFk55uwG6BLLTicsBSsWal850zIi+dFnM0MDZ3HTUywaWFNB4RVQSCjhbD51W2PAZC8F1
UtfV4qSzZmDSLl98Ha/358ZPyuNiIwXodyKu430/IhPMcY7a9GsYAj3WM8sGn9yLOtMb04wOBEj+
wXPJfNSHO3zisK4lD6kuNw67AqSnvH88MpbKId7+D6+kjERwVby2pqIBdkUf+WBwQzpbdxwnzCHs
Lr9Uy96qDMTuxbYbFtFlBzJm8AtBip8fRKBjquVgpkgF1SrxNWBFnK3/91P3nj4Uv/hhfPevkr4y
srHiaWUxGkaYCyFjfJGv1oKsLc7bgfbLx/Xh/nvYaxEl6tAonv9vWNkYZ7PV3F+8fI0qFWxTY/Pk
des2JBOAYfz5/sIayDcofT6Xpj6cWfz527KdjXqsvYwks0gIN4mTMf4Xv0nEZVwzQb4lH8/Y2rYd
IEiFxU3ClPGnEI1zLk4l7lENWqoeg1JILJ0pmbJJcrAz9Fp7rbd3BKXvD0N06xzUrVNtHZj8XQ1O
JCdC5K2ta170oMEkcZfpcxPpEru7Z9bMS9aSffxPGNy5lI6gSPO3+BPTExBtugpe3k4UeRDpYr6U
wy6mAOD8bRUL542uO/xLqJPFLQf2be8MT2cuMgE98EZUw+UpA2BfpmejK9eAYfnlPDum1/bpradh
IBiJKZ6FBl/EEG/x17ST1EpBcjEHCFpgpDFPt4XNwtV4sUrvJQKu98Cc9LLpYmq4rClOsZjPVkze
+YI2TP/epXEnAJ3WMnN/KFsNMRXP/mbBTVFVv20JZ73RNltrT6Z4vB1k8b46KxFLcLyiF8odYBrj
Sl5Cd41nj39PICrclfghkxXCjIqDPVGwU3XfRYfvHcMAGkGCJ7UdSlmtX5+g771wtUTMx7F2yYah
YtEm382isSiGXTyMOmp7DjXXtZ/uMUbicPfFMPfVbYdHZjCMkmh6M5pvTg9794iTubt2rB17NpzF
uFHtTGzijAKJxRUI2znTuHxjw4tVy6CZs0KyJxI9mZr0X3BktRXXsCfKyr3jy/5tXpeoZhGK1OwI
cSHYeBwHI1ElPJxmFBlbunGGRXVA66VNICcyUBqS5d4ONFY5NDHawXyxUS27Rk3l9pFa6CwKZj+O
oIYehCuov/e9/vmiB9jj8BDUMS/T2BsHjtl1S4H/7ZxtPKKGrPlQDaMEGZdoX1Eiz8qc3PuXQhog
b5HxVmCSdhoprtZF7JLLgxdooVLwmiNeWBrTWIMzDm6SWWmKavxqmGVJtx1oRUENVJqOcKNnsunX
WmT2fkOHGh3lq356F8km/MZ+ZRZhX46gH/q2prelxCf83B/5ndkZORnBvt/qGnpLkZI/n7AJAt1X
X+gbHkZuxg3UVPagMk5XnK4vKsTN9PDpl5MgjBWg5YrvFjh+7V3RP4JkX2bla0OwSfpb8v2hqIaD
SAjIWA7SQWdoym4yReZ/iR0TdqhIKckN+Nv/pcHuckpzl99nY7FB5qhq5hHDPX8brx9/0LaDz1/R
RbCt38vpxEjY+uJ9/E2YILFGHNaq2i0CthOfzkdP9YcovnVUvZtr15s68jfVuCwvFHO9DSl6oG0G
gQ/MwVck0kWEC+5WA1YV/GL+PisH2iw80kSh7B0D6vFvKy1lJjwD7mBI33ZslxZpSCK1oiLTHovK
iDpZYzNshtViV41oBm8QtQbfdfpNEaYHdIGzTHO8M0oKjufhiOwHxe/TwEhZDmjPC/xIw0L6fanH
tgpbBX+Z2CzhkOR1rObuw6Yr/92QxtOjPRjz/HTTON3fupNNpECmS+ATB6yTPYPblVmcu7dS9OuR
+lp5wzYT0VFOYu2soXrY+F43nTSsTOSufLrN5iWUicLO5pnCSvjcgMuuRwO+DqHfniP+OkGTd91J
Mh+ap/GXg5EB5JWiKu7NX10KNTE+g9+7yaNgx8sKqbQY7zp1M12dasLfXgJPHy/pPrOUVQSHzJLe
yXCfPu4lsvFcGQcFiEXI8iKUlWjYLQOIEKHH+VmJ78NlwQRQz1SCuEbANfCdya0DhsdwGDpr1Uiv
Kqem0/xx8efRfbXRKkQuQh/2zadUpp08pm7VjN+1R0cCKS5Vvnm5UgQWPexuRcDDBCJUd61PPfOV
mYnNqtCtpE/SAOpPCqJbRROonHpzW3ltowObqjs6SG/2bdc91uzBnzNqL3h4kVRcP3noRroMxV1b
cwqfUfVBJpAVj2bno489tf1UyWova9EiFzemyr3TJ6I2vbet3wMpaaw0yOc93YO5lZILVHP7Z6M5
czGv/NtlNVG5CpwmeUn/prsPP0/6v+ITMKFVzGmvDPkPUA5G+DhpyPtZlxkxNkmL6v/RUjqnW62y
5IZ0y7RrdB4Bz73bp1/oVDfzO2jj6NhrM1NifF3YrOHPpAcyzQ/3DKk/h8lfmjd4kuBIi/8ruRt2
hJLCReUup8wbbx5FlGWoUZCRCc91lJN1iFBOkobJU2mDlet6DET4nhkFL1/5O5Orwu5cwHHUOcrn
ZL0TB7EwIqABBfyE+sBGMawpHUK7QHc7Mh0reTjt4XEwd0lxXOV6R5ZdUdv7jILHVFGvfhVRiziX
cWsfHyX7TfPha0kDDvUuw2pD6yOBnGjw/Q5Y3Bx0tOUPbAgg75Fn0N43GGNDcul4ScsCRkGqCNCu
O3pLIfKjKbxnWHBZHPJCqaMjOldnpjBQBWkUOXRHDIgLJVh+k6q7/SoBOQUbxpkDZWMvvcr2VaAS
btHAIZWNrO2DhGhxVywH/io/gvL/SQIzYnesGuRc+3tIuc2Bq0yOJOLTfZf4rX3RVJtaDd9lJv6X
5BhnKELSarg+p5ObVeABHhOwv9bPioFjzNeGJMjrnwOw6KZuNZ84hyjUPie0sgEJ8cO7LQ20QsiG
ZaC5BpkAhXAtz9qy3YpfEc0s/KnM3X5JcsLAcuMaxynRrt30zQ6UotZhKgHXnq3ghy3aYxagF99I
QcWUoEa0cBohqwHzy6YqpJ59yh+lNWX6fdTXHA3SZ7dSxmxzU1CR827NYybVzFfbQqwa+2k0tFtJ
+IpAQUtM5fygBK1sQsjKlcxYzH126JzHuyq6ZUH/ygVQLRNl5wFe3WjwzN7hOP/LGjaCyiZywRGI
rMsRSpGs52DgFC7RP8Y3DUjZ5c/yHaAK8R99z367cst8oqam0aPrK0BdCZkJvse3gyyS0G4XhNFv
BoakZMF4uDKujzop99wZczoG4y+llLwdljDlNh1PnVHAOl4trFRhwDcNTtudm7Cyn1Ref99ekMG/
X9iMmUmME2ga1uuOctfr1Z21qeAFwFyDwq1f8dEtIOzOZU7osCHtULcpqJqpYNXQN6xNWjMOWmOu
pcIykQgTbD8vZTXpX3B9raQyBV1gFpuAlgBIobzhQOGRt+vYscC5uTsYYmcgKqQ+EDeGssNnlJCs
xk5TzTUbRbpKf7niBnUhVD0QdmYRAcnABpNyrLRbVyDYvXCD++4SINt7H2/gKN/MHNyJGm7E21nd
3l9g2K2571D1FoFDVZk3PYSYq7j9b4iLJmm38wgsm8uFSNIwhlgGEpZCWV2qEkXlCk3k+q8hWtuB
RACdW1vohbM2h0OHbrx0MRQMMkXdKTQCfQ1aSo3dpaasAC7GhZNsmGYi8Y5mbN2deVIAUcVw9MLm
t3pChuV6NewOXcMR0psIhI+zz8Xm/beuXfjm+ix2priI+lX2iEn/llgc3X2yA0K7PGT72SXtpKpo
CZwoxkykQfBkjtzQYnnMSN02u8/ZDMBge90x0hMYl+1nVHAdWrT7yyGlO5BfHltOgdfD+E4z1RsZ
4fVhT3YlcpI1w5cRqJc0cCc6jx0a35w4czXQvkqVECSquPP5NeWxuF+OLJL78Uy3igVHKqulW7c8
Kdkc6oOiiEWEHrTQX/WGCeKerx8myCwzNpyi53SEdDJ1RgFw7vUYOTZgVgLq+vN6vd7wGLABWRWN
XjZLLUkYkOZBWWCP/jQeZN3zM6Kk9Av5OqMLqS/8gnBDnT/S8djoZWw+LImSs9n453cE+bGlXjlS
ytQnEwhAJxaEzteM9vrOcirCvoA66g17UwCacczIo+4UDLoNocec74s1FfTUQT8N4bFn+ME3wFgz
0TXyd40o6PDVE4YqxM7pB6/0/1kWDfOGwKQAuDBBavgZEa7RN2gxZPE9kMr/8B9EdATPEW7eh5WO
mqkSZp7WGP1Mh0U17osuhgh6n0KkyWAjNbjWJxcoZtzFw8vq6oFg8FPCNSZBcXUsfqlR2khG3orr
qzS2PXnCNly68ZxwfClhaYdgNIXgKS2JsdiXaY5NtW+AxH+lzuKoygPnbmYS+IeD/5M3az8FBuEC
6yWOtz/Zr11vgA2eaQoi/u45wZzduzxvudB5KGtXtequgGpbrNYQ9XHnUwSTxPd0QnyYnXip0ExY
xf9x+G6OzKRmky91V5/TYImsfTEO9pBfpF/3Fbwh0a+Exe9Gulvcq5Vqrskp4SCjKj8MlTGd2P1T
fgmNTJ29kqsLuQ9RPuB8yBMfoTUTtiJi6GGKF0oVPEPmEeGiMMjgo8DLx11EjZ0LKZpf+EeL3KFS
kienekQqoZg9sIL2n1ceBfgbJp1/TLEPYTsgI6vJWAxb4lIyTuyeBKa5IqfcRDjUXjOv5/99kYg1
qIo2RY/A8nT/+OgvZZeiLM6GKfCmpSwFb5zGBBDRDrL5cTKBRtQE/NcWpyAFJDdtzAx0r9JihCGi
qxznzcyVfggsxyYlV6XH3fYDvIdzl/0DDljFJWV7GeKqsytYLSPy+yD6iE6w5Jd0z4ZgLUv5QSzU
BxZXimQIQezUkV8pF/pLvyJ3Wf3DAe0fk6uadh8vTCz/WHivEyslPxNaZe0YdqpDPa+wVraA2he7
EizRjebPwVBjbaCYKmQpDurc1vrdEAKxsFWcijhB6CoXj7WREr0/qv229vdGXMHmx/SreC/oTWDf
Wz4tusIhXw8QUxhkTzcZOJsvrs02kw1HEm3zmyVhsxSbEmxvHzq2O9LH1Of0i21+yMk69P9QVxhW
4YsT2m/XCVBgvWjyRr9VoGb3ujhd515hxUiQXtRB+Xzm6y4pu/7oCi9H8ShB/aORTktuPbY4pBic
8OmRtw1O7XIFbKNLM7/8OIfg6RAXhzUiy2TeNF/LgdzBTEYhZHCZVY3pnA6KgI+IKhaqQEIlVgIB
iF7UrbcvJQcvStRYrFu3H4jgd+aFcfrJEminkBxU8dwQjqaqyv7vw2nzSto0LoHXQ475mTEv+S2C
5h41uoQJsCcPBvvoB21yjFyYg/0ZMjV+kVqu2HMnMVpMIa3d0JyGByryKNS9xT+3oiKXDDc+Rmb8
uJtoemp6mY53VgQHq1pF74x9pXhBaPyDGqugvkH4tUiNoeN3TvF60QJIPRNgmajt5yZAP7jnCIQ4
97TquFNYdrXJ3RL462YJSQ1a6wVdWUYAvE4LC28RGet6V9kh7I6keuFItnF4dhO+C+EfQxaVYYlD
5NjvqLsyOM6xK7w396NEFgDfG/omE7vIgabQwFmc12txGwy+x1nHLYdh9Q64EnaUviVbSStBvU0r
pnHgzswdaTUbqJOYL6fLdnc9FEkdqLxTkNVi8jer0uPG6V8olBvbLgvNQCdZQBSXQUr+oGAvglg9
QY5MwhuwBpTiBLnK9AOG0CPLDBnokfCsB3kvyubTN+dMeXU0P0DMlV925TcUR4sjOnP8KTXEhEms
rwYImyIiXB90WzRcmhrmJo3hh3EGdwv2nXgud7OFtryljS/lwcqqfwg5cWuTAglfIvRctnTZis/5
qpPSiGYXTrhErG/LytufY17tjdUpUrcYWiw/gtxcg9jDR7L/A10DRZrNlqjzKjoVQ2P3u3OVAGOf
osvuDguFZ1ZUDn8M9WJabuD/OZSOQs2DR3uZPmEDvJoAslYHpDh0ueRj4AdQ/9ZQX3Le7ACHOwHC
70AG/rwpaKMGR/KNuv4mVPmRnGzvTdiCou874SmUNO6tyPzA7YVmYcxRWdq6CZti+KrkaF4rGmBx
ddmvd7F1uG2gWqxlgCr9/9FHcgR/d4Kyh1R9NKumy172uK+T2Sj7sWn7QEZPVAZnYX7d95tJ78ya
kEhev/YPxOy8EudocRfIAuPW6lDLi0hVraOnP6vA1/9zpCLJtWmij3+i7IPTC/fj4XkyegqnkiJL
sFgC/gI4x/Xnw5jsn2+ObWEQv3GPMtQ8kD7OyGhHPB72YYLIG6nAENNWNmxqe628X59/J9hV8TUt
lW7+h3+kpVvN5WBLgJDJkkxuqf5ntt0SDOqnUXv8sxcRacWRyVZZcHMh13Cqq8MLpwkiiKgVleh9
qBaKvTxYhb1E4XPIBoosn0kWF2Ivk/r/7P10WdRfsCffA+3Qu+EYpzT7JAWzkxZLiS0ND2QqckG+
lqHNXtWZ23SBSZtlObwX5bOe01d1AB5pR2wfK2rA1phjtj+VnBaBaFVzoXPVuVvbfrHAo3ypazdL
KCwGQaK7L0WfSr1MX1aKBqnf3dqL9bafU9PBWO3Hufv0weIedv2Otl53x92YPrq/g4aKDKkg32FL
sCXRYkBvVaWgnYqLN9JnAHLfeH/y3kDO8UHgnKTiLfzK8m+/5FfpLS0ZDONrJ9HOdTLelSg7+U7i
pyVfit829XxDYTL5X5/YkCVvLKwUgDBVhv0N7E9PHAS1OGDdsBxuwQfkrtCYSeIdI2QhfXH99waF
xii8LTAHFMp0zpDkaRTOd5eQygzmRf8MUtAO11lWUKzNVJPg3HdhRgKDd9YaTzQ31y9RK3h9NUea
HKegSS2Wgfqh/Mj/IKqxXgpR4l8p3MXIvuPpNWZT9AJfqi87HXyClMuPAB2Ht32HilJk9o/+vlRS
ISWye+HKYJ4KZDWWSOgX+0+3XB2iVIhgJp8/Ovo2bPuNNv/dRqt0iGasPhzywhtT0JPjpYaZhxuT
K80eBeX4FvSw7qjioBH/VpGrKhMhWLzdJ5y84/7ivrL2Rx8SRlq8rTfbPof9X/DcodyO3MUCbBbc
SkMtkX2KjnA9sVuqrU61jThMH4Al1j+OfOhj6jIhW+lv0LcAYS10frRnEN+0fOwTqEDH9SoeM0Om
lWs5aJtWJLNouwJVK2bXfNBg1+Ytj5WO0HJPZcl2kZCHtm1qXxvRUbxDqr4OKEJ0IPgk83gmKK0d
iMkiOX94VOLaOE4+lJ5s14IHTP7VE6D4D+gobL5YWLJaSeJFygZMj+0qnRU7IBxrIW8Ot5y9P+FC
90Icczc1q4xjnm0gf9dB7NpJ+nKqhc5mjVe9rfpVEgJ5phdw9ZLtXoyMAL/bY0mW+23V4xMV3vOp
xaGpy16KW2sw+Pd3rDig1JO3WWKjjDCGp3KblDrMSXZdaqRHjk+rzTclfzc3qPsEAsZx918AWxKr
nX5c7IfYRjlO4yEE3jltip1iCyVVSm1cp35pjcDo0yiSk5vrvS6oRmtRCbjmCwr3m1BFsqr5Yab3
FVRZIJ96CESMvxxGWPO6lZusLEHqxe9n6GSWYU2JQExWEgB7cJRfnV+xRENGhVaabptwQUric/XD
rwLsKzgswUGqNJrnF8NPOCSWvI1/eAthEH1E3Cl/GJmrqFtaSuPwCumXoB0Gjb/ZFoJoFukOXi2O
UNK9gp+EBQ3cELsb41LVitiCnKymSkv5g+FHLTwVnPD0TzN/hdr/MfN1EIra9CP3mhmm/ZAIj95V
puTVuQfDh8ul77w9JuXYRa9NgnYPVBqNSNUTocvGmAvTIvawisAvz2QmRGkEkPzzxfmmgErnBdaW
fRigU/wlVEA/qIUp5+Oa3CHTQiatJ8fB03EX/hUuYF9K1ug1GL6AdSQ9Xc06vf0Fve8DiVdS8sAi
Y1WxpVW4oiAvZzCyCTiwlVQPLrdIiLjDiX5O6d2ZdOayYhfi4yOa2Ifz+ggtUYWZG1JNYUR4eBYt
Qd0m1bnJu/quRAIwDT4s8lVrivk35Sve2fGjFNmEcKtB06ElJF0qsAR9TT8wIgSkfFo50nZ3FfCn
7pDdkbNdcE+2AUDZTBB4iQgjpE1JpyNh6brDZcYDWFKINfkBfdHhkCuj75rv0Fhe8eV5a7zmxdzG
dcONzqSd1Ar8WmgqTBxvqsYa5Sccpvusx+ilaH2reK92sAYmOOLqX/RfvNYgJI5mSkCZaeCQ4hrx
8ps7wGve8eQLTjz2myyGVu16wOPuiafjriirJ9d+Y6e69PgaVA/dTKCdwqkb/V+S16UaSNvtW+dw
wbT+RXUHmYIZZjjwaAAKeAlFSXjQf9/Pvb9zkA9kmc2J+mOQhKO9xlE0Dm3TKyOIYV2rIYeqcR8d
7sHkB+/vO5M2dakdcG+BnZKuBTa1AvjxnWRwNjImYJrai0m7ZeJP+mjdGLXIwRe3sYS0trSqD+DZ
usvUlg89c1OkVsOk3eWPJ4BWk3trYTh6tHo3k1viATcM4ry4IoWItogBCghQ3OtTDFvCd5qBssTc
6D6Po9j8Zd9gpaNeqVWdBbbUdAwRzjd2OP7tWMG8ofezNGQ0r3AaN+y9NKrx0wSOfVb+rn/yn4/I
bRYVceanahkOJD3FgEBjNVEj3onztQsRtcpUeueea+WgL7DAGdzIUQfuwf7zYWRYJ6CIqNOFfJNe
q/j3j0/vzanXmYBHn85wCM2NmSD8qVFRjDgfWbMofZEKl+dRZaYJcLVs0huPTaTUWsE8JmyOLkld
E7dlHM6r74sysHqoqE/oOolKUaVBuRrS9YAFWPVIFnmG6rKZ7zkm0R8EuBs1zegdHLEU/r8U+ZUl
OueKM9X+3JgD3bgw8umUiS4V40zkrHkKEhb/aNiKWzB4S02Qes3om+d+mHQINUitZ+gapCfnS25I
MJPWx1pMcJ3rIed8dq2dmmkmEeHrLjaHc+unZ3AjgaTbh0MWmwQ5w+ViTOjGDmImezCTmoU6GmvR
/NFE0YHADH8HZO4NtgIe3d7jus7oHALs0Q5Hc9DZByVyQjM+j1miQNo8ERMU/YgAEK2yw04BcOtx
XGtG6+CE4RiXuUaXC81h1uj/IGLrYvWK3RHDK5ZLQvxLb/PXj5AJvKCPZ0uLWQkw2ei1B4SjT6lS
H/x6JacnrZdIAIyLfBdZQu3etPuiUItS1JHdEhikExv/qFrTihKzJVSWf6z+8H8lDl65bM5xJRlg
xdqiB8NR3IuALEtrAprbMOefbWptUFdju8pjA84Rik2+x+WkaN6hFcTs5fyczMeQA89sshbgkdVW
gadOGB02XCRfcL0IQtJMSTeIQbXuVx7GwjQWV/fSHL+w8huvFrBxDhxLooSheyB9UT7+PbfjSkA4
MFk4Zv55YyLdthnU0LMiVrIIs3IR0iBfHovfeJ8rXK38OlRspnP0YDMT/Q7g24IwWF27Md+woIaw
W+wYh4yeiYWtzg5rGDT5KFjTlZyG2Aj3p6CPvxr/Aii62Qn7A/b1fDY9LABidAU5K7IfrLGhUwgQ
dKxhALy9zAJzQsoLIsYjQpCkgnM4nn1k3bDRe7HyoJwXiFagMtzyRXyDy6mFaaP/cqBuvALtIlLK
zODiAb19wOchVV2ENllCyuIuQEDsjpB7p6M+AiHC4/ltEGZ17LKVRuFJgSrrhTtOpF6rE6/DFfgt
8lVFLy9hrUQzzx6QIbYeKuInQth9jP72ylGp4ZcRQwEs4yKasQyauj33GQCEkgXVIuniuZbBAQOJ
kBlXJO94wa+K2eZENDsJm7wQ8Mn9hG5z9CmNxvpLOkV6Oi09/pmJN4IwQcwQgir2z1eDK8OpE4TH
n7UiC+lxtDHtoNQlvmX1jfP8xhQ7LYHOwTZxFiHMRnEOV3GUk529LF8dy2/jMazdmb8r0fp3FUur
9cpfTpyq+TcboFfOsV+kRaOegutNCK+8K+lJU4gIMNKAMXOlcbujJLplRycssLCBBdlhNduhc4hY
MDK2+L7wxlLSD3HKEfhM47ZI0DtYKzimXPHnIOMFCZmUOfyGOnK2naGh10kBoWnzxyJTosRNsKxC
+6F+s36auaUQvg7kfTUy6a62TfaOuTGMdyeEOHlLdGBWEvyu0pCmdcHZecN0vl8Rt4Q/tff/iERP
TUD4ilshPgWrAAQsaop6DkjqtFoNCAdrzV7vEsAQBudNeKZpYr3gFzlaY+GCAioemgvjebZYkfQ4
DdM63nkwdt0Boq6LEdzClJGRlLSSe5XODprY2gyiGvD819sq3mYQW/X9HRtCMqkggX1V5BIrC2A1
gFEa6UnTwsHpEB4MnduaNOKvuQjAidx4uBtW5IDW5iT+qBM3krIwmYIJe/0AK0O8s/xfjQeEZ/jE
5D2LBad+zP0AjU1wrIiWOXMAHMN6MDIUgxxn/iAR2ZFPnYHwRDCbt+9aKRH9FzeTBkDP9Ep2XMdz
Xexxs9K29cQccr6PL/HNMsTe/kqavcusa0f83GXigHhDs4+Sttxwz0LjQ78srWMzCuLK+zF5mbPc
mv4MbWrmVKWFsRhl0+jatn0pKvOEOjskccClD1CUSdLw7DDnPkoMxalUWITe+0d0dA96CQ91wwX4
pip5Jktj+QiY7Kp02RnErmgcjC6Maq4KRbteQExeCcqQpBLKr54BmG6nBENtJFDkwjU0aZsDToCW
xP9M8sN0P3qSwiS5D7An/58s1J0F+0jqDcMjvRdLpU1vhXeTtEPdCflP3QlanwOiaND2tmHASvkz
+BLRbZkGJyCAsGAp4Kip6jbgUFdN/qkyucZUv8fmnn7X+oi946QDGPt9s/eng8ASsPvtvPRnUAhB
CXAF4boYenuyPTw49y7jF0XAywOV6BrRkpIp39yfwspsefISTnRdxLn3IKMbsulyiQJqIw2WrwdO
oR5E1OSRW7v1jU6I+gs4ceLq8R2HUVyMhnegGG8Pff/rXRCdqfm2tZkHi1eWOITR52w/RLd7U1SF
3faja2uepERynjWFr8Ezcqs+TCwD5rFHGB9xTf2jS/wsc1/ZObGhbGZWnnwCZYH+9Xr8v5hDWH05
zX2yseYI3oyYpZh4H/RdOCr/GicDWDNNXlKKYO+mZAkyRf0HFrYGoJKqe1NM4KLGOFGxJz+2z9P5
cfjFdwl4TNi42SHoliGGL9Dhk5UGozsC5Vb0AU2vFM2pQR3PzqRUsZ3DJHrI1kmLS0O8AX6eybML
WPvBYEsgqyyGMVKCirAhJcswNd00rh05ISpcjkmoh8iNWfonh1fwnEfm1TrkhgZJczAq5hg4zxW7
tIeBRYq0Ygs9EjTZTp12pGRIAe2K4yEJXVL7F4YLawTQsDZsQmdgo1IFiEk/oGllGZEdnXjk3rip
0KtPNhXecYfF46mYmVSCFkjXVOh6ghBbCtaBU7dFd/LyqZxZ2wnKipZxXWD3lxP+yOjsdOqg2qFs
ayVHU70lr1KYpDkmUEH3N8ymG9eBW9AOqECXSjZgibUHyaRg9EUWt5r064r5MsCi2lKsA8DU5Bo2
mtU4YzUIul59mekHwMa2mHT3WPE9fskvhYl6/fI3t21P7Yx9TTnhxYB1wOCWRmDSnj2NBin1dU6E
4/DY+Evdl6YoaxpJ6Tkrsddbo+m2LyK421uDJQhXEoyVGuwgEMxdQaMbSOmg+8Kt6VJvCc8SlUhm
T2M5PMM3UHXe+qLllLJl7m9ubHgZlVvXKaBEAmwv8FTqowEbE25yvYcXfgit6p6simo5e2VYTYZY
UM/jwbMuagezt5kyYSMUXsQTsQxaRsuhrTcCxdiwmjrtKB2/9YqS0pUkb1CIPrYPD2Y5cNknxMTJ
LtY68T8A3AuPruG8AXGcQRLXtmBzkMelZ0Cquv/el8sLm3dBhXvHj1qUzk77fTBxdRGqMLpJ+4zL
07DbqLXFzKzLp9kRg0dR0DlOjmv4lnZiNOhvE7dVcM3frlMZ+rMQdTytYJW+txoO0Fql89Fcv1do
3ozp3jUE+CFZviv4BD3ZCuJ3kCQIihShkNZog514vrcAEPZdZZ4h9O6wY5wa22M4pDWqwhHT6yUk
JeQkymbTt+uMEVk8W+V8wl7ioRzstHborcgZ9vArio6IYtvDm/JP/W3jYpzEdQ0XCyzFvfIWKg9B
E4v4rrmEGga8rWv6m4KPLV5Ps7qlyE2XGgcMXn1h53o/lI0wGf2Xok0Z+YtTKEEZIestN8sEKvZn
Y6W2my8NVXxzrhOKdVIFsmFM5SfUxtIAJHPRfLQumB8Au2LMChMruoE3pTEr1iYW//i97mbfQkjk
ydcmiPK6KkiHnDD7GY2Mlw5bSkvXUywoukyAuljHxWWiKnwra10K3UR77/JB5cv216z2YGsQqU1v
c7O2JcImZxQt5TaTEJULuZUHFzD2kTvuGmckAHOb9gDNBGmRT1B884AG2OQcs34R2WPIu/IUE/1p
L34VwwqpoT8kE+1w5YSUEEdt4x6rUFk9GmGe24ZloxYqnDkjP1pUkrQh2rwYDXAx+KyjFBLDSF3d
qqmHXiiEfzBienmpCeY6+cA1+oJg6jiAE+/yHKxGOh30Fz9mjobgA+9E3vxzrgtj31ALwtuuHMHp
hIa2ko/Xtb2NyM6AuOQdPylTsRhyk80NQrzBdGJZJWCRLnKxPDunITmapdRF5G1J+3NLhKp0sI/M
ovNiizx6fwFrI5EHdu56IENEEON7mT/kQCIbIoeuDHQkKoDx/j1019JJnAWQorpf8pjq4zXCsl3o
TFSdrbueoH1qdtKn9FDmksnPrY+nOqe5xJ+d7/j0tjXUNslinER5Fjy+inc2CKRr9B4p4Ml2VcXs
RBEHlXVuEorq8U1soY/lEv6k2xx0jVi7dVoux57xnI1huGuZjEjNewbAJppnZD+l2C+gbGwoqSUw
AnJ8Nk8KpHFBcRzgTblsD2zgah2ZIO+jZuYbzxzisfbFc6qL998Nn3WIcq4LN1vINXfBVxYfFEOt
yyBminf4IyOq3luOPYSqwZbVuwTlnUUvVedb9WnMSwpYVzj2mQjFqXL5wVDdpAxqvJAp8vAXS7kS
3jsAUUshaoXBNheeMTnR12j5y7XwNZotREFrtKQr7T0VXoANwLHfLrLDLxitXISwB0FTXXstsLNj
q1SrP9tKvSCI/AzjTpydCsERerONE7tCaHcTdFvk1KxQukJ7L93RjpDIN/hvM5s4nUE2OXx3T74K
HadY2B4AmIBKUq868yZbzK9UGRWz7wEg+SqQ8smlnYMR8LrpiHJYAdpuWdnJGuAVgpMV3HcDILdA
FDqvbl670QR46ruP/XGrnzgohK3I4EC0Udy1QehQYTFcui1SnyeGI4X3MnnZ8xVfxBh7jcuzib0J
hhonRMP9DA5p5kkEeq3IsaGl2Qb47lpbaSIBUSyMMUBGeiJYs6URFl8+HYyUBU6MgLIGRhyYaacN
z33m15vsobeDGrJZBg/ynLGAXGufyTd1Wn9D/GcLYXgxBcsGAT48hRu0xcT2ViPNbFbVvvF1lnlG
o3X3EU1R7Omf6+SsM6NIxLjlGJFf8jwx3XIpX/4ewQ0Rn7cmkwGqe1mPI4OA5IbvuYG+jnVXHN4o
tR/9ZQWTqPrLs82Kitcafy4D5nzP/sO6K21VDjlYxat37tDcYJvyh8AgIeY/Zmqu7mTAjTjmJP1E
W4NnPf/gvdvc1V4l7MX2kWvx4fEpFK3bR8i3eg/U4kp5ZhVSN0X6Od/IbNpGpqbi3VGqJlua3v7H
pKp5Jy5vqAaOekNH3jpsQqAXrjlN0kgO2E++dis1+bP4LOResYoqzYFNKytLw7idrFOkJE+4v/BJ
vPgtiibYW9QTG3zuQG41950j+hFrIJV1XjH3i1y6d08Kox9f9BVz5sCcOxDBeMEvnBIs08zrN0iL
B1DTS7pbaVA9LWTCmuLNFdMcDvvC2qLZuqP8fXHy27MHBYW31MbiFTdNzmVtJqshF+y8HW0ckjR9
Adm57SM3bBREBZCVAwJXrPccRYSvlbH8ltdFbkyHq896AAU38dxQhszjEVZaq381SshctostJIb/
FAivKUyh/XqX3KS9EtPo30Plxies06wWEtzOsGwcW6B5x4D8XBuPUiFpy9KYyhaNZW16dcm5cOGV
mPQwprz655ruUZUvy2sGdbpkk8lGJRheR98qpNyRf29XspCrP3Ytk7SgZ8/Hb+bPgfXR6foNjSZk
mMiVjGltCs2mnIJMidK95faCce45nBsUMzhhbwM70qD5cDZoitm/1Hryl5ZpxugGlajg0zShk3sg
IJkacRqhR0unpsY/aZZcIdoRkV6uXyCKit3kr2kIuDqTtXcBBR53Op9mn7DERDtLlWb9Lzokv55W
3rVhrWfEsWGdrJSnbS0tww0QTD/4RLDbDwOrvkVHJIOpk36Zg9dmyN97sPsGAOklTO9b/IIZiiEa
thSEAuERONk+4KPXZ8b5up3ql8ULTUv7Xfu9rHazHJyQvpJEVVyoH7UJKZ/OjXipZjlL6jUYN7Dj
/WB4jxeQZwYE/5DRk8B29UxrGco+k5aF7oC7moH233Oy/OWBX5DGlPTe9UgbNz90Tnemq5EpaTxH
83sX6osCYM7jFEBWInsTNzOKcVImw1VIUOEcbIDMHl9+XNfj7ZjbCXcc3D72EOSUjWAnMcT2AEqs
DMWnX0+G3Dbm5VFBofXe+vknNNlEwVe4jh6V/yeDBzI+nQj/ruGVtQTUZAp97kgqGcw0h9MwByLf
mAsyGBbWAhKNmdw9fRmyPGGS2kD05phcajYVb1OQixV7Do2p7oeN2D+2DxGi4uxXwZaFqt1ra1Hh
Sz9xqTs3NDZ1NazpZvl9/baP+TKCmOIET3QzQ+GuJ4Rg7SOZrTmz5LtSZKcWuXBGJIvCM2bu0e1n
DQlqHlRKa2nmYsTp8RNPPIGgci79vjW3IIn5BM41fSTiaCieaoE7HSAdFQtDo1rXCs52q9gxa5Gq
t4Im3ToshRuQQrxZtI7CuvCz2dWY7OzhtcDB5fozYtFgRn4rRzBxy/zHTINxpplsm0EFcPORb5BB
3OS/hlrNSqjW3YYuPQvH3DiLS6n26WaK98RjiyB8ynnkB1LHleDqG8VMHZ6Xsfzf8lUHiiNZ0Afa
y05EuZ4Z17Wskb2yPybgWN/0fnWBLIilwVTidceWmsLk6DEH5M3p/Tpo/CP7YBjEcCSRbVTTgSqv
b2f4RKs1C8MYxvmMDtlXmpWktNc0R0CQRW6EmofE+GyBqthKhoR5ZHqt9fHaEe5sGFhvTCIMnxtH
GHdAkl18Soqib5b0qKdpHPMHGbBDVNuITlV9Kmpi9viZ/7gsqNd8znU0PvLiRpJ4ktVhj1xQtJkU
qzPLKQXykRTEBtK88tIy4z/t2C+N/lfqnkW7bSZX4gth/OdcZgJ9sDKjU48jL7MRmt7WsZPiw7/Y
13THbugGr2TWSgwAnAeZFiCQ3QL+mH0VgN5BLiyGsMQJ1ICwgr8VHr42vyLLU6BQIhf8nBJqrzaB
B1LCJE9EQk0FdNkcWKyR86E2uS+WWAQr3BvVTcwyaEEtU4ENWSAnwvPcErJG0D+0W6WETj4ZYJJ7
daah/ZoDoLEUI5LG2kyot/L5TlQ59NYt5bdve01ceDkSZ9shx/o58JvkwCgYW8bMUVcdnqepOO5F
ZKj7qdwJi60bV4DIu3p8WTo4TIO7o1MsBmvmfqDtgJwie/y2H5yer3g2BGJjoUCNj2Ru8+HHyMem
hxRKaLSh6zWO+vNcWEUxPwFmxtbgBEVCJlQHZnwT4qrOEj/Gc40oaNUz3hs23bMSv+PHYp2WmYzc
fFjC9zDKzMeEKl4MSG60SgqgGC7yZCJqa/AvH0yX2xe1XtuAMuYg4ywVJCSdvBXiD33w2xH4znCQ
X785Dw9+gaMzqayGzqzhK8J/Ulf5LJNws/5wDiE+k32DGivvT2bma75jhC0tY4662TQRx6OAp2OI
eG0ouQ51tbU4eKxzi3z3pvlv4J6+v+cdDzLb06CBBScj271H1vzPmrkN31cQNbY01DV2urRF3oEy
Nioc9iXIzILSgmzNJARqg+pQ3cEX1MVUk8Wjt/RiIs1XA1O4m4qiL3lM3hOu4Thfnt6AeCtWD2KF
/P/2RIQ9xZo0kTxYBSB6COm9RZ4MJr4voAZYd8Zg71CEljsdRb6RblrAj18HaasDR/ymECS2iidI
4Q0/klKSmoUvlCpThpM5NvO3tXw18ThHT2QviRlt+NROs/jEs9kSbhCfnLBTiGAw0NBeV7IpSSzY
X1P8fkZvSwus2173V4b1icX0n+Y0b2W2KVLMNAvftvuaPv0p/2+B7kq3w/1jTLL7GrjD7Hj7X0+o
sV/S8v4iHLCxKwh2WPqiqpk0Jnbx1RlSnO5lFrCYR7zi+RiGzVsPeC+GraNte5PaCcTMDz5yKSFy
9aRdv8oTYqhjpIHVysAnnv4TRLifn0oVA7rJA3XQPYD9FyW7gK5ui9X3D9ldF6GlmRQV6y0O9BjU
jF9gVyqzw75haeIg4Us33Am1tnkPJ+2x/PFHttnqO12Y447Ky5OxbM5pKpoX1F/W2zpwRQ8Hawz/
JfF3+yfZj0783d3DN0OaMiHe4lpE2Lbqll9tXUChkTpbvv9qne/c0eD0fXJ3fviydak3dXqjgJPq
Wl1sR7HyUcRY5nI0IFo48iODJBPTR1qonCn5hE4Yeq/wadFVEW3B4q9fu5+K37dqn3WOVe02/o6Y
gir3Lze4j25QpLJauxNDrz/lwh9ghlmfwB2GnmVtiaJUB5IcVWkwqtGRd1faqnHg5a9vxAV3E3TM
97bbMn8NFuGOgII0JxKKAV7/XCuILuD/NaSHgN9ZwnRd1dvPU4cXEocDRMu9wF1h2OYZ9lbQErYJ
CCKD6H4+nDWJZrKq54s9msGt9EfksVmLfm0abtvb03/I0j98z7kR0cOoeS+mjV8UkJh91m7Fb4va
flz8QOKejyMbkLRQQQ0awvCAs7RMYIqe/JwF3VVDMeJ6Leb1PEcrov3atVAzTLCQxVDZ1czezn/X
2AF1wx3G8IU59rtgOV2cD/fAYdNbfDChwhgKw8qC+4T+h9/BRGyXvwdvI4PjK39ggXxOzqAHHXL5
1oMC5GZE0SD/J8fLkgstFb5RTz3hWf8ojMz+PQddcniThUgZg2V+Xjs9z/idTqg+5JzDCjY7lHWD
1qeYIxI0RPBs81+sAOfslVJraGVJw4arWGEl7jLi6Tb595jASe8KPo7qvut5xY0W87ZjO1RBUOuy
sDrcFrpTYGV+DkbyQoRsbCcgOUsMZXeJc/19UGw+PieLuRTsmndd+kwnr8B5JOI1CwMljwkZcLGt
OnN/4enxnoShG6BRfeRAsMTmEepXX7UyDPpBShySHooA+UlY549w4V2N80LZvdZfl2I8Wu3EPK8v
qSJEbbai9uQCgQuYQ/rHp/6RMyII45Qi5KQerNn8xFlrc+PO8RzufMNCTHsh5eQOvOvdaKkj4AM7
OajCruQbdZe1EP71Du9zTvQ/XfgXLebWbbMFP0QKrxPJWtLk/1cCnRFayPf9UyNwAGfzaAPqa+fz
OF+7otGpBQrm2VR8CB3QhGG0KdSbxf/RSwcrR4EVc2bJmm8xmORLgfVl1ejVt7EVaxeBWnYpQJrn
+hgt5SAZCXAXeOZqoYNulDyw4SWvu2HJxRRq5UST79RgXD9gbi4MuFXhc/yyi6aN/XXgJ6f93GWi
tLO4iEx80z6/AhUGRVs3/f7kud0DDw/iPMx9h7usXxLhPEXd8fXIYMgeubWAjIB6SXp/kQF3O8ff
Q+KQxsEavyCJpzno1qdbm55FeRIi3WRfko8Db+K6oq3kR0/c1cOmqYd9fp+kiw7H30ZooDrScR3b
wvjwh+dP1zoSXj6Fqth3X5m99xxplypTH+njAFgJJX1eHeDsmnUdOB7HUubmjAQKU2LIkHnJbURw
b7lEzLUeJevMMCyB5qqR/2erDbP9ZgfDTXuQynsP7FIFfrOKlW+30QidVZ6gkLvuLF4d93tRTYne
UpSh2sObp3KsaWht7nmAIeTG2ZVCrh9j6NOJrAjbftbsop9S+QD7nRQSGL/tvdbNdM8ppFf3oDy1
LqR+LCT3q9guqQZXE95WGwrOwgFzik6/BaWbIBKEPK6LFaTMLW94KnNOOb+gAraU/mvUcY1gWl9K
3hbWKVurEh79WTQgt2JC//yPwrIJB/x+gSmg8Oek+x2a2DEYrWka8yTBUaeUFa1hY61eHzy47nkd
JRtICOO5g4/mKk6fVz/S0hedDwQ/OwW2pmGXN0YU8y8OJH3+31uh6sr3sbIcrA9pCMCa5Wq9r+yH
fcGDDF044nnmhdRD6kO2eRh45kmkU0Rwu7e2YGcpV/u8WMAfq5H+/+sKgt6KyAJQDTdBby1xFIpf
vrTPqdyxsRVSo+nRPJBKt4lpRwKaWtXky8p0NfQNHIvTHS8wtCVqSDi9dJ8nT2cSk349yBT0Q3HV
LoQZz/WOaENGkFiBjlcZ8HKsZVYW0F4zp0V021plp0zucNWtgaQmgbICTu2pNKlJs8+lFludDuqi
YdIzwn6mGa9eZrm9wXkPGQ1jAjw6Q/5teAc0evFnphJllxcnr2YgSZVjop4DeN9cHSi5yGAU5p8n
UYAzmATfmqVI7002uw+ZN5DS1/K3K7p4WF5hSF8sZ7b4BSQJaAp21N4YzuPqSalujX9hGZzMCc2t
Yono8KjHqGU4wRWk7+tbV8+Wa89xDrV+XAW6MHmT9LOPw8D2p+4PD/3XlN1dSm5SYnbOqSMFYGny
VbQDPOL8u0jXA8zJlC54GwFJF5POFMrr3Sjs9yDHW4WYpDrTETCLil71ZUUBEFn7KNN9bah4CrU8
g7EIW6TxxbZXwkWz3puS/SGC/N+e/l/nqUE0Oh4RS9hOentPGO4Gl1LskHoxdOcL8bT9V+e80LGR
KktI5yG9NCf6BEnvxIC/1grGt9XLYgANFeRYVbQye0vhANiOnJs3PqiXYVl0Bj2dMxYMb6w78FrF
2X9amoXC0Pmi4teF0bva0CxZMGXZQuXGQhLOEo/nDJbE/SPGOVXYGrXB3I36GDNbakfVlxOmlBZq
jBpiMs5O5eGFDZeJjtbXE25rf486CfWwRydK/AyrkrAalzosj5ewUhRyO4q2Huq9zReCL17bZ72t
e+VzWa3FLJuE0cCGslREoVi0ZWk65HZRxBQNMtxXjvSijrQPxvJVESwht8MOFIUlQ9Y8p9/nWaxI
u3+Jp0IVq4qjE0FdsNXzfbBEyO+xflZ/b9G8iRdrr3XEUasXT+XopSts+M+JIKvVxyJwm2igyNEF
U9UfQgBhuW9GRDDrTIFbJExsHw8uKKP7zFt2ByRCR1Y8WBsVYOXRRWPvUrMzYyvAriL7tf4F+Ybu
nYBnYO7mCNQL2ZEVM5HM6fkAqpnksmQCtSr77/J5kin0sbD4bFW6edRn4w/1SlJtw/srvknoueVW
Om2+5cmP8yvl0HnDRaKTjggxcSOuj/bh7+GywyxL0NyiTFhwY1qVCEPjeAQMhAIApu7qs2dTL0jc
lpbnbWu+DPcnHNVmKo3If4eiuuHb6Rh7blwUDk8h7Z8ylBdOTzyOFKwZOoS4YEjXMYjPugYgQ0Mb
++MDieQWaDAxcIgDTZAEumL0G5JNTxO8J0SwcqnC2yy3raFaAwxjKmUlV6zZIWur/G1RrVZJoUe5
66Fjl5JxM0Iwuvsc12bSTseNOoKMJyy7u3wEOgPN5FTbt7MR/fwbhAKADGOG+KzWULrdupL+FpIh
6mJUsmh16bFri9uV5NFCHTgAIpcPlqHK0Tf4e2gpfQAbeARzqLQooiUH5Jsy3pHKN3u9ap1Prhy0
o1Wd/WmVUR/Exutu0RfwpKUTuMxPGXDnUlITdDpOs/umb8COPiKqB3Klz4F/Pi+icFGGAGfk8eP0
b4bSaoRlkhiIVk126K+osyXMdW1aIjZbwZJZvqoGqI7K/G2TKuS+6LP33L6eKQ6Ir9M0zrBBEe3K
5aQ59YFD8ExEBoVLl/JFGywOoXnf7e1OI8JwCtheWnXVTq2ugNiVf2t4cFjkrioNqSlAGav2/kpJ
9YoEOTkIHGrdFVkbN3QiH4GGE03MsUHofijXpdJpsrzVNjVG8lXL1JHBSeSJeC49sxgcvAw1dWQ2
fmM5AMZIOTrIaUFPKeeK+PVTCcPSj2DmYe8xf7DAauyJmUNzfb16lGcQROsTSJRG/r/ej+SYZF+J
XMNx3zpxQCfbEDYH8VytOgMrThiN6g3GvMcNcRnlJM9vjCADbe+eDj0gTzyK8CtvsK+e6n9xJLl8
4TGlbX6fvF7UwrYON18RjIsBuflQ/e9cwNFZbCbCvDk8092eWYXvXeb5YFpf+utABtvcpVYmf/Hj
URuoVkd4Az6CTmcFV8qt53PYwNZ7YdqqFNh6YqXJOKGBs9D6Rc8Rq04s2831KTBdOrGi2jiJUPqu
bsFMB5WmcSV6bQFFasHKmCozS2lslL/8axLOwGH0UVXQvHXkMcDE8BKhdKvJSVtv6TY6s9oudkHO
QyCXsRFwHkZZ8H4Ib51C6wQN8Gmw5LV08eACsQIu6Q+puwfUoVZIt9qrx+cYskh3ttPhR+JRNffO
qCWVFpjgUMJhq4zTETZq02E/EUg9fFZnwDWM5uWnwFz7bf58T1271GtbVt3pfnqwNj02VCErlkWP
Nv3oF7Lm7YectZCzwlEts4zqwhltoM4Qls9jg0mMjpRe6uMncEAQSJq50oq9PQlUlGjRo8q+5SaZ
QChBJJynb9Zj/+R2J3mGbaKyEThYZloV00Wz5jNiEBqpRdHWJcnV9vGKibgiE7nTysr4I+arCFXo
OUUPntz/+1WF6Y3SC8f95O/+z0YKoT7nmHLSMDDXmI17DJ/tQpHfg2nHWE61qnvEBlneUePv5tV6
jZ5q93fk3n5gS3m6CtMceD7w0GlIifnvB4iZa8lzkh5EHx5UqwhBPe94EVIbAITwqIUsNFXfiNxe
F0Dk+Bp3ImGLZwHJl0JaVtik83o/h9JCrZTrOHwP/vXcRNF7uNsfC2BbSCQjbqUeqnKK9DaLZ0v2
WsyHamwGN2b4DlfYVD09Akl8V0ywBqKSolLvz17JD0AgPwH8zm8TaRtxoXfp394IMBCvhOOkd/zo
HFxNuf/pDoGWOjrgditXbEbUgEIKCZ/0I0P7dZkKDz5Sf+jzF9jTlYeV3XmYG/5Kjda3r1IgzIQ/
Zod2/28bxGGhcD81tk0ESPXREdd6Pm8AwoJW+zWMRBDXXwhyxDoSgaPa3PAB9Yq1UFxLFvGi+AGq
Ba121uYQsgiCI+n+tPaybiJtXYz4VaKLGddnjbXMdt35d91JBiDDxqiJQdMHynt7Bi9ylYVZ8jOR
JRXNv4hA1OES9otdTn8eiETNQKX42YqmK3ZiyDajenekVQTwmldzUA/U4YQ9sRuM5bbB80UGcCdV
VSByw/lR2UzAu/qLk/Yy/vfS7zpEMW+hz66OCqHFZnkPCz4/tmoLQAMwaQ8s+PT4qIE/d8lIJpKU
NvoXn45HzYon1D6EXTHBG+PCaWMZIjXRB3hyc4n+5A4XsN0m6Lk2QuCXFehHlZnJpUILiyYnZhCd
XVQwcNvQgxP3JMZT0NauVMlHjcUu/s3MP77VaDryKt1DycsxJ3upeJyCZB25o5DakvKvFTTm+O8+
MTXSy2Ex3hAyGPGdRMKLbzYn7pQDm6DGJmxjRQvQbvnH9eDYgrQHRIJ2pw2agCJN/gD2SkhrueKS
Ubz+h+rxwV42jVE+x9bKnJch+AIYxRiLIk8inhrl7VUDDn+w21DlAgPliALDs3DAFf410ns4isgF
rh5RAUYiSxSKGLGcjcCz6mqBJGdqRiTIRE7b2UX9EbmYlYvCPdGw34Sbp4FWhblbM33ki0daMU1d
qR4KNcpnQ+1aXnRG80iOT9WPd52RJlUD75tsRv0Rc6AzVPnC85HtYK3IWThQiztyDvu/Oq8C3mMf
qRqQvNKCiTUJw+gkwWUnR/Y2gD01219MLK+bwS6Ui0Vy4eo+q9dc7MmnMHC7t4qFuUo7M0ilXLgI
H55ayQr2WYSqYRg/hmzSkGiSvNGwByyoT/Fza8AY7fgJ8v1L79YCWyHL9i89gRdpgpOSXVNUijIX
rMFOhJKWFzt2TGx6rnYg963pxaTzKbNtaoU+dPJFd9DqOy98DPWuaB5ZyS9CF7dEoLRt5DVh36IP
wNJVZ7nTBjrM/7mL9qAiC7321sK078OtaOAqShjuXDUUVj/KXOsiQWkhUzXWh2faNh2FmjSjfMJS
uHMUrTZ91S2xBwPrn4eM1FnVtkPWkHm/nuEUIVzZJnn+87VvvVuHN2vAI+wqBd60C3h4S3w7rIqe
Mewf+u3WFp2TfBPuqBBp48VcdZNT4dWKI8BBY5hFbCG/hWEjcs5wX5eD2r6Z3Yq5jmP9aTASj7Ku
wdAbLPU9ix369K9CROkBPMeXFdW4mfzst7owFBjK148TK8Ti46jyFq0ic8KzFcSprblfMWlUmgjR
NUS8idO1jgmjWc6lzPVxkXo9N8Mzfwe2zfqYfGqhBPud5ZUS35+1SD11XosAN66ZRrq2YkVrL8CN
XpXl/DVtGsDViFIgQzlCW/8Patw7XUghJuf8gqpesubP4jUohLGmfSI+Z5hSf1mMPy+9K6w7V9xM
GnR/Esznv4duRuoU7ojrO63xaW4IUCSPxLnqGHZkK3uNhFi5bw9LrwiVXl1ZGYjBRRKFLQ6bjH8l
aJ32pc7QeIb9JOdERL/AAr/gc8zBPnXYR7HGWvLH4Rlnr+k9HakNp0C1rrwWIK3gdP/UJZfDUwDA
W3d8+zo/zevesLhiTaBxaJQjNOBUmwEDGzNTUCbpTUkdRbvXDZxgaS8+wm8tdliSMv/XURVze8fY
ozOM/mTPVCniKbWpBlSI5X2Tdc6cZJfumFhrXTP0K75ByyvTKiVSU5hawRO/3NqHkY6OM8gwC18l
hd0IeoET8VQtftCyvzR00EIR/BoTgNTNn48jEzIi5VZQYihGjw1ARhrry4qMrbpr51BCfQt0oKgt
WffO4YQ+TWoAMC2eb85eddx1FopIKHkzhz8bL+pytHvtlPgRnWo5uFrzz+IiJn3O32cF7L6oiUhV
dz6Iy4WB7ku1vicR7wE06hu4F7wauiLIjz+Nsmox2v5BFvzLqx/0rwHBbOwdCHXX3jxQH4t88Q3s
V9R15BA7eFBzxZHByrz1HlDrWXCrbdgoXxZ1VLj7EMBPz+URUy4+fw4f7RlFVdUxQOGew+/mbtf5
4kU4cLDU14UhRZLH5iAkvL1OKdlt5eKLCC+Svs8QfGCK87LeoCfVGjxqvihVhNUEAeSqSx5POecw
6mHKtl0YNOxl2PsiMKOubchKT3vQit+Wcd5bDBeRoe2Dcngjsz3qA5bSGzN0qRdefc8oPHyFVS1J
MN9gcGG3/c81MA67mv23K/9lqid5YwJxf1AwXmRv2ZTgcZJH9nW8hCVvo/6Iw5SZQVWjTdFUG/43
BrgGkd3BgcukpqqQbwsphvelN9kZL0zqagjPdUEg0UXO6MIMPYKezYCB2m7yslzcFWdCN9LgPPVm
ueBttaZCyVtfUQCSlKBJ1xZIl5Jbnvdc/45dFmICDetfxVjvc0/3Kl7EZU6aJpd2KMfGwkzTG7xs
trFnYcbQ5QN4ziXKMgFJuKb19cbgdEcKaZP6YMoFPvhWnfFlIydQ/2oa8IC+OLDuFpBG6IZqoMfl
AXkiKMDIUPrvNtEWB2uTgs5EsOvw2b2/sdkcUWTg5sygrBmTtpuqm3Gay/Q2Wmlml5Fgje/4z40E
qYvI9vN6dCF9D31g2mtaBymCCSFXdXAXDhVWZdj3jdPAy5gYRDZj9gynujCzNoQNlSI8JjRJSOVK
yXMjYME61V1PY0b5umiG85O9eOCLTbBlpjHkwFjuENwDxgIW3v1PqrUfFd+ye2hqvwRT/0QuUaHQ
gkiOrIPRDepp2ftm1HgurC6JKdJWzbDYzCU4YN5Z9A66W4ju9wDKbqasj9rgRxbb4thWpRN/Pabm
nho50Qky5EI2OKuLoNcwKMVx6ikWLxZE5dsH7AA7BS/hl4WQeZfJQev3Tvy7cKTQwERk1aAhdhVM
F1mJdKq7SXLSQHGjjuRSHUTzw5gLduytUZxNmMsI2MTWxvxL+1Ne8LZzQimivnbIKyb+fZ4gdJD/
iExbKnWjtHWYplj101cCJb4DzkSashtVZpQMxRoXCllrczFa82qcRmUEb/ZplZ/Z2/nWzaCl7FgE
Ml12ldN2UjVel6oEEJOjoIng8hYY+CdPCF24zJmhWabC4snKQUG4dfb/0zBao2E3OwFUoBIvya7l
NQfq9mNrJByLGkJsxG4BP9mwG0WKfzU1fZC+jUIETWNAvKmgkYH+wCXstczpa2xvtuZO2GaJUiId
3l244OK85hlOOE0geVlFUgY+f/m4C0MAIgA+41P3f9YXhvj0hsbXi0oDX/6sFimeDn0IqxsZk5Cl
Juwu6cqr0celMOs/x+wLyHL9H1GiqKnzh1NhnVO8kf5z43tpxtZuQ/9rcansK7WogK4DEDqGZe0C
L2XFuJTjUYSeehj0Ul3ny0dQpt0tsG5uKwkyRHQowajDI9zo6B6y152ebiLP624u8Z+aWH7T7B2l
GtPCFyml0zv0XaaC68c6E9sp2ONtj9UxBD8vFDKlynIEUe6c3Wn3SAygL1uQPxyobg21+vtRysQY
ihfFWRwGqIKeHVmojz4JbZKD+OwBD+5U1TY/SXAF0zWq+qKKFIpDgs8Njx26xEVQm4eSPYmvx7fL
59Qu49FahaOTl8YwiaLoxej5r9EwV097/fFz6CvWNPReVB/BxTLQTxKsOOeajvYY/fg1Yjx3JJAr
TxxFtbEEjii7c+G7fMlX6JmMdQMQCRDhYbU2rQLYHgyAfBfjT5V8A0Q5U4knhXggRFxJfisFKMAa
wUkfOE/t58Lwr4AFMgwrP558PwC36NBN5muCRDqVxZtX2rcbA4+nAhJr3RV3Jo1e6GcZ9qZUMQeF
28dX4lKbwyHECKTFQ9U5zvs+DOw22UG4IMr2m29IqRgOSiqrzmC2EMZVZ3pFnCarvqTEfUc1Nroa
fyoHT2kddtDlwPnSYennY8m/YVNGQr4oRAWZFkwNLSoqnll4umq7GMCT43h9Yy6OkJNMZzvc6RYz
SriB0hxmfgIEeUYMiVBr64w8eUpps2qou7elvnVbJlnMaoSPTFzT8Hw9wDht+UMQ1JeWWYQ0t5ve
JiOpJVIAYLGN8YPR30evWurvBrE2yC+FN1GN286XbRAY2FEr5HYAAAnKUVfqpYLQNj7lIYyrxydL
eD3xmCZQxK6PLlU4CXGAdsZbGeJIIhxPIkP3N7SO9fdo2iMQZpdQcTu94OH8sJ3uEguDBNfbIHBt
eIEoG8zo7/0RHgqgQ+8nNm8q6H/R2PVgZjdo/KXJG7x9u1rh62W4CsUq7xU78vTORMSDNRj5fuEd
zbjbieWG3M+Kd0VnRvFegrl0sFPgCRE7bVTg4hRpug28iBmDqFNBtk+1y8wOiNvz/bqpXBwcVic5
uhKvl7djDjaWuKOqel7b8ut4PZqxWA1thhKfshZYxxYm/ZHiEMDwlNSLBleMBk/kRwFyz4EI/rRJ
uEiXF/yqXXXbDZv6OnSmhc9WQAYiITQqxu6lw6q3Q9f0utYj8oq4dbvmfK7wUJPMSOyj3hxsQqda
EdHWlS20MAlV3GGLNHo7oHsXfFThdjMaWSgnjv5lUKsl/1Gnodd4rJ97x5ejvvOkHh4eXEMaroCx
LGpyWnxl/sGvu+ZMVl0aF2T0GcDiatY2JZPpi+QrIoOt1yh7RQy2N8lT9w8DXduz8zU1Uf0X07Pw
KtwnrU+Xuf+h1fj9fnh6pK/w21Q5JmW7R9haClAbsmzdkoWePg90g4PrDOPOGTE3+AFiff/9eg1t
Ac8w0MESGhfY8FcxMNJBLEKJoCc+iJV+8dKSdGFe+M3T/5oY4gO594YoewKZua5ifL2ELYE/DWDx
zRSYv86KeEvr21/M9d9v5aBPcM48wVC22ci5zaQTsyEn23nntIObZDBEVIP6YBVzSkk38CkInwgY
4eYC052o0k771AfRB6d0HUgVGJWUSyakJCoogOe3klYihuq4RgLGsv2J08I0prpV6aN80vqryPBL
RfNi1BMTA20uR26rwOsB1CBMiY8D8cwgUS2CQGr3N4obeY5YLp9/If6cezfNwXZ5cEYt9rxgnRRC
D4Asdvtu9rFDs8DBd/BbJDtxWL40pApnS2ZFw/Pqe+nAlgEINz4oJhetIeG28b80tp4jQ0Qjqc3j
iyln7T3SJfRfs86whgjhTuguryqiyVQkR2pqfqkB24vqO1vtMJtkbKCI7kIsZDMJ5aYK/LtGs13+
/msiWBrlF63ZvDwjyCTkbnek12bqF9/dhEnA+eH+tDL5tTem10Wsqo8IeAZWEgtLGu0gUY+MQF9h
eK6cYvSe8ddS8OvLY/ok/Ly5YBkBbKX7Yb9lknXVF8ldHJD+Ua99X1PiBSCmjeT0v1J610SfFGSQ
bC1iCekcFju8S06ZXyCFVEXaT322glmSyM7VcW0vQjP9o7KvwO3UVGG3xcLPD31ee2ObamJ3be5e
okowbb/W7oZ2veATBV+l9bYeP/FYEtaNqhrM+w4ELcC6QT8dXQyXT30sJg7wBgqjS3KBMGMQ4lQb
PbWUqhYJObH4Vi+LIpKnBkzjzGWssj94+gFgoTwGahtQUcFzfFO44dHkKNU0homw/R/JfvKZZXWD
ofeEsfcLz/OPJFTiKAPrw5H7H3RAWUNM12Ddu2TcFf703dQRpPh6Fawz4vywNKXboYIE1l0j8mlT
TFknu09IOSYWrkr0wNEtTWa/bHSUQ24w7HNTwJw6d5KFULT2evB+02qoQl7haL8h5Bs2JwIJw632
Zl+2gRt2CPpyo4wIWcqfyLxVB2PRZBE1cplKWJs86y6anprdmwW1tnwAUQfnNm90IAblSA8vnZC+
QaaOEhjejH4u/Wqwuq+LtBTRFlMMzHk3ajrzFMA1l6oR88xWu294mSWzAKd3ly09Hlyw2u+to2cx
/DWsf1w9ZxK+u57HJC3+xGQsqvAPkSCxecbN3+pZtKemNN2AIXr/ltkcCUselWSPvW9UOCd/qmgU
3AV/umoN4ZGD4vvhb2Z+GCpZPQQ/t+2onPaHWp1PwqGvn1J7YHkQWBBbPL52nTGFpxhvKozMznkS
u0e01guhA+ej0+74ktiq1HdviXzDqNhAtg9z6Xft+E8M4uVeyTrlIo9k6ydMEAhz5GyYeRxE2Tq+
rsFmcgw8zfJ633Ycu1ETe87dDDDCXOjxxqCF3srxTaR2otH5e1Bda3mE4Z8nCbTOgaOi5TEWl8Dd
ByWqamKqEJBoXBYQj4kvRJq8frnyiABq49lYFeo7p/jOPysaHbz4k8xR0NmrhKFuw5F4mvIK3XrT
aUrY4dKxJvin7xavlph8GVWKx6gLLHiHhH9cfn2Udj93VYcm/QCxQz9d7xnS6qWzKd4ibBoPk0kn
9M0jgTLqMN9gZc/SP15pt5s/oIA8I7eKcLag65PIdV+DQMh6j961iYFA5I+pP1u2gKzsI+NeUS7z
+HR0W/3X1FQsLgwRLyVdC4XGDcXh6NW8w9GcGhyAAAThP+xURHuEhSOlMHX7jSwJduutIEH73JLF
ZOer4mWDt1IDNQZMDV/DqMrBMlqaDBvEVJ/pe6NS2F/nE0WitvRc+6snZnIreDRnZF22wmPysOfJ
gRFt8+ANOIiaVELE+olUarcuHAqlCZQWAfQ9vHptbt0jHLZj56rsRdyn2SaikCDpwirzXV8m88lO
QvnEYxMs3U+InqIzCgHEhgnLTlgpbBtgEWoyTqGvxHLsriP9aGw/S9nWUgp1BvXG+QsQutDY1RHb
C3gXlPkx5Jyn8GamEGasloYHyBVmg+65+cKU/KZw5ixQzPgaer6C7YzWNO37yCykCaL2LXt1+xk1
2AeQfJmzrBSsplPUhhcuMrku4kPZtYUDucAkEg7slVvhE60EwDWYob5yCfZnu1ILhRVJHBNxHmL/
YSG3xnmA085z2hlOYyoZNdY9/UbFeBPf6ZHLF8qrRjZanVW3s7IRiJn/+k7pJbPuwJ7HeXR8O4Pm
dNXgMPjxrNzeQvUw/A/vwIukVb9RTU/hJLaclYE3pA1A3XLy0URHZ1dJlcXQtctSp9fgpqCoJbXU
tthSKoqUT/0IeaHv2SQjV0eymSW5mIgQET0SFa1m73idB8tdK8zXi68F7zkCUaOLrCMYoOTWE5mX
oquDNNAzE3ZGVYnNydy0Ps/Js8TE/DSShUmOfvzjNQPLhbtOCH1Vkw7/Jk9ItHfa3PH0f6nvzbRh
+esk6uj0uSKDuUiybKGTFoCEzEBr568kCth+VqHPVt0SFXmP5cbI3fv5axmLVNOm1FGE29dfSuiB
Mxe4e7tcweG5djTCSouZ9SAmpl+Ig4m+1YOcFf/5qjvKlhbv9QRrhxI31XvrqptG35KOG0MyCH9W
8o5gvKluEDc00J069yh/wBhVnS0B7rMiGBtNBJkofyH3OomrRy/lLiZJVb7EacjbRu7WRVaJBNMz
ktvG+Wl6/XKTcjbswyGPGHSHAwXuO8zRSPIcS49KbhW8cbKALFPL4dBprr+nH10e+92CVJn1NQ48
XZWviDzgrPVuJbJvLaipGc57n2y7BMrHPsQTqOlMfkuRc3xa10YXBsgjIdCQhw+RKA0mgSeQDEai
hPrhI5OKkUna9e1FjMxLshBjstxHfLZF9A96kIAKSZffG9loienSVEnU4d/jSUuLZpyXti0Ehliq
z7znslmhn6332uOzASRKtslkL+mLfncTFYbgNNGVBIQszKQb4rj5/32dHv31v7e7wRkiuLR4CnVD
nbGCgIOt/mDdOQ9QCOns/InvGtFo8IIL1R6eZsJu3ztyrm3o2qsqVzJ9bGCRyLQtObSOh7hnV7Wu
z1dNQbifsnjCuVIG2/IPrE6SkWUUjH96/jBhrqoz6mzHPVh7VrIhjp4SGwnkrhTCr6Q5DqLmjCY8
+LRkpXq1bf8y1fKlEWM9uwgXBydh5r4nBYzodfKU2ybZ2YTpCDOzC63EX8NbD9l+Q3tj1pDllgDS
iEw6c13dOP47ADt9ErMIwL6n5HguBFQcLfNV/NvaItfp9++/KoHftqwHw/+hvK6fn4Gwbcd5bd2J
McOlqVxt75YCcitPobvJImaqcL9eEj1DzYcAHw8C0+djoL9GmbYMMGLhK8WaGohoaHOPQo8ud7HO
FO4eAfar1zvyo6Dmz09YiecsjawpALQsB74sbHk9hmINuwud0e+9b8FdZHCxm5TgA8NirD1ls+dD
SwTEnWCOrYoYmGQUQ1ej07ooTT/aigY70WFG75G5DevXDxqfCr1ZbPLhp/2583F4ByvesH+2XvAe
Kf5d4etXtEeGtgdTPhvehHRDFs2TpkOtD6DI2b+Mpy2ubjzE2UPGlkl8YX1A6YqE1XTBQp1lqpCz
XCmrhXNeCjvCo6/AXG++4ulwvh3RiT/YYPNl+NEJuBLqmaPKxwTFX7/RK47DGZFg6Dj6BMDHYuCh
pSM1UmTYwc42lHAclv2W4DWDA8/MVMOh9+RR6w7pgTl6vn734ofMRW+lryWzXonj5YT6iwpw3X6a
tIr0grhbwDdNfXGQnfND7sSnD+vu3jV0M98OJvWGe+B/7Lj5GY3HpT0TiHXuUIY7DpuePZgxLDdW
Nv0x61gAdHbHbuRYgnBufFTs59+VCzdD7LvhTDkaEBPQuyJvimwIclJdait5OsP7/LU96tba72+J
ris5xrNFy9aM0WSOg8zeF1U5apOpN3MvrKRIUOOeidiJ8HPSCT+AnfWDe2pPaCgmsrthlXvoX5Ab
PCnXl6QDJQhBdioerXGNYZsXWBBpvvE3dY2Gh8B5AVrERag2Sk5Yck9PgFhMbdcPwse86ZSKi+7U
B2q2x1fbKVKQT8tkqhcShCboKbYJ2Zrlc0oZNu4NyUAgsw9CPIWc7lqhoRtAo+LHNkc0BGpThIEQ
bjGQfCBdQuSZDCTBK6P8GvtLjlxlT+E8FaqFHGiccQVB9cbQI9/q7/0NalgRbZ8VQdXEpithxUYP
og1VwhAGA4n26S2ztiCZkclc6P3llyHxvgzN3utpnAAEsBWkeRLfwdSU25deaQSS/fE6mrGi0WOZ
YoPWyPbmqhXOEDwm1cCNw/YCHeIrdaZMpqVcg3/yvjqU7nNc4+B4ZW8DGr5yKm+GLRwiFZyw4kku
xarzsiqx4Fk+NyXPg2KyVYYs/roOwNqhbWFQ5hDa2tj0Sr7vshaUBvRvObHPo9dCYw3IklGkfXg9
b+dZDrpwcOTO7cHkK05xgSALrF/pb5T0nwmr4Bl/qTZwXUt2m2+1OIoIFmRUNCPIexeNZRxOYZSV
U+SGnp0eeCNKoyPqYqb67YoppLYYLGQ6nmb6FgnhTnHwuQ4HV1z9I+1KUI5j1gqy7+0OISbGbDqs
oV+6O5IKy0WZ8Q7vw0diDN7qeZq0FRdmpi5uB/GRKI3+QYZun5BjtW7NlG9ss22YZT4i4DvNf/1T
BJnqn8e23IiF5RYnOL6FH6fdVh2SnrIQf9b3hIHSy/DNUOKSpatiaIVFxB3mPdwEaS1k10VoF0YW
rkFQExAuywnOsq96zL9LtJ9DoKehwElFbBEPFIRbCid/LLjGcQhhYLRpUcJWehC4ZqqC3qDId/1m
vbqvHIY3DMWaapIRs4QHZAW42Hb6gsx7QeyjX+U2KqEMDyOLAETqWCal+nMPEcR/9w3jnA0C1Yop
cqedp+cNIC29Z1BNEd9sC8yyYsSrebDtdRFUuvtYVAIQi7JsxtiXcK+HokGbdIs/R6+tqF34C3ty
uBT75h5leMiY07mbSsjPa16v/mFSnk+iMP90MDXdZx/8WBEj6VZKNqdTd9XwPcSMhEzoKhTGxlzM
JqUm/XwmREy6qJKGnNOPrNvos9Wa34ZTuj25I9c0ucAEgcU5TzNE4oK8gy9FYtE+/C57XAj2W+b7
ht6lPhtT5QXRa+0xH6t+4fc+j/Q2BURH6JM/EmwaWdI/tfKiSI4/V6MfBAQ2BJ5x237VyXTX6gpR
Zv5LuzYgwpFsXoWTpfXcRANnXErtBOYIvfX2JbZSi4mfO5jBFavLnPUVTgRyChyJH5NbDxwuik57
qsW0B1LCEvd3MU6rbQnFV/G1k7pLbx+lB3bXoS+otzzwfmMLhGBu7TBCUPQSUAggzENz1ABacj3D
z+Ht2TH/DgN23QmOk//0yOrKeqjBwNn2CkFSuVX1SjOul1qkomEVuV6DOYum7c/Rr6hJBo2dDP/u
5go0I/IVDa8W9X2KrROHOW1WnQh/RZ4k6ci2xHUyn4xsykIgfHQs5ZW0QteB3h5klalYeq6W6Uqc
eM9UvXt9NzIDzIR7md6IvQe2Men8QFy/gff7cRomYqpcE/wgTc5U56+WxaQJDR6b1RmXh6dDONQZ
tiMYwczHDbYqRNbMdnQKCuhM/23ltXvOhApnHY3N2L6T5amdyMXxNDcBkvmskeGhEJO3SfTHVV/s
/gYYRS8SASTRoK/IL1NMxexNxsk+454Kb3WqlivLqw1Hbn0eXherpNO94Tn1ofbR0o6jF3BoLcrx
6+F5VfMMfRytkXX9j+qp24B/uL8rsFBjF+lIEe7I64yuWe+Huwmc0r3LK9Le1YR6gbWpdpj+FHNN
JP/V57Z3HXREcAy1+IEUYw3yQ3OrY2TtTFq3Xufz6OqhuO+pPU3t+dH4v1G2AOjr+zqShicfgkft
L4pCciBtVdlCod9UhqT8wW6ghJbU+qq+lAFiZZWyVynb7iUAGMIb9rJc0Y/KVbMLONMiHO4jGa1h
r+mFm9UNIw/gYU3pgHpd/vr+vY2MKd8C7ZYY9ietW4meTm9igcecC0IEpsZ32TaCy40RtxnpHqyL
WwaMHefQ0Pcp9QKul6vZyIlP97yFWQMr0D/aq5rMq2KRvwgYn2GIxYjVbIexdTl9X+HC/h/u/x4s
R3L8+GjRJlKsy8lq87/70aErge2XWKEfSqX/qw6MkniPbcAXDaPjttiuAfhwFx1j012tedcDjISN
hZYNl1FUBIQcXeiDRZ66CKbtH9zJIizRYtYf71GQLPYC1CJFQd2vG3tIQY+Bara+AkPb4OdjtYhm
mU0/7yqGvlwqJV80yvmPUR3V1c5uxLVEpDFdmOriztw6EO33JQK6eflDkxhroxD6CjH4732o6Trj
eYmzpBeFvJ4SAFTHZS0TvEhe94gzL9Otdz6+yCZaI9j0e8Mj+gU48axjh0THdP6c+fbmTth/9vkY
T2Eml3B9Ssq9otxtm03mVaJW3HGna6vc6mMKUe5j8i2Hu15oRvuFa2gmLRyzLkrsrz4O5sPiij/C
4IRfrY81wat8JSrzLcCO9nqBBA1x8y+1RdC3avtDKh6z2f1F4xa7vyOG8kU3V+Ogrj1nDU/1IW37
9Na+wErEq9gwGza6qtarxcxDw4vM2Odjfo+isidQf+5+YVG5vQEmze6Fvgb6M5/nGq2XYadcHMGl
oA1HUpT2VSXOS9+DwD5LDdkiE3oHGRldObNDCWX2kp+1fsqzxknDT0Zqp/F/BGBqNLFeIUPjXZB4
SfioXW3T4JczOr1d65FHadbuaggF2bZdzH9XD7KMXyrLAP/oLrJ4IG9p7DQ9iy1HSyxUg4myUvDD
YzUXBxbEUiFYlnHEN8V6WK+hgw+Pwz7GPQvzKEEsoezCXpN2EW22vBTihkB+a8YAm4iCZsUG9zKc
s6DcBWtXYpoMKRpwT+tzmmgOrNgkJwUJ3vdUIn9hcBLhi6qIlR2NsNMibDmyJ2Vuok7lHgHQQFSx
3c44qmbtlt/VbD5KycQTNSZtvbugqJ+uVaOWABLPWti/+c9FJ++kQQgUC5jddCf2vRcrXQ7FX/m/
7xPIgycPMJ2YgYzCPZ7JQlgGWAUDFULIrXVFn3Fbn4eBS43YJKKolNHx7zKazxL4ZS7k3Gcz4D2l
6evcI3C2TY7igC4ZpUyR+ca6rKeGQxHWYSIXmv8xXG2pG+soEkMSO3MRLC1rvbQHRbtxK4JEmvW6
5n+G1uSgIGFaf+iFHFX0uet7a7kW/3/+nA5ci4qSCyg4micl+GvLuyAAbcJSOmx2CCSc8XDFhGo4
AS9oLdKB0/nSaDV86nRPnvJ+hAUJ2ZJw2++R5ZNgS2VJYsTB/CIrtwoe8jmLNqQelV9VklyR5xEG
nSNmrx/4OEeJcb/GKJUy6iCsT/4bmOQE9p8AF17SQY9mKEy8XNQBuLG5dsRHoggQPmGVrInMagn4
GOheoM1DEtAQKMRVXiizY5O+HMgKh844PObmoU2CyMN6zcFQ1cFfBodFclwlx16saeeDVnLoJyG9
zAfpmmU0w6IjIsO3+db6JXr7oQTABcAPr4Suh8SEstJyqA1jsbNr+OOxygy+lmPza3C3nBRSOnCa
nd/yplimBrA5SVW9OP0EQ/tIY3ulw26x1F1Rb6zlWxEF9WO+8uEIQJs0sVBuCTAWF9U3IHUPcRMb
s3Z452gPKXA+7e4EKBS6PrY74P3Me+cxHszrKdCmP3eQ6Wmnvk+hjlNV8QMIh091005iCABat9Lh
De0NYlZb4L27bWxZkhwHtOdX/1+lwxcxOxw+FHHTDRVnmhlKq0JM4eNQBmIATxYXm8U6qzQfkwbZ
Qtrkb3e5gJer5Q2qggKadKcJvSpNnT8x/KPWqDnWNTupM0uC2PDkJwlYeaREfrVs0yycMjjxX/x1
Plp0RFHRIgiNAtop8zd/aOsjt+1c4qkDzW35Liy7BKnnbn/fOE9JhoB3DMp28JTU8LJDQH4XwmVE
2S8gHyv0QU0q/obdmi/+be+f5BfSm5vViUvlFEX4BMcbZXzNGUhw5ApuhiUEsciWblkC2gbqpVrK
QwYvzI60ep5cs0OJAr6jgagG0M/imMg0E+zvaX8WlfxdFUwtzN4Rkd7S3WrkY+WudJ5rrkB5xWoS
nBwLOQCgtrAgsQQOco+bhRJgK1m+86Z5h0+Q7NzDzzphdIzQgZA+v5QQDqK5rORmbv47pMjboJpe
KifQG++CZ1js8Yaj00fumrdIZAjbc9AWtTPHFj8QZO5JEJq8Lv+pGuBVQauL36RnqfQ0KhEdwkgb
24YEnxA/BQrd32kZxuT+JrOXmD5OcOEciy264/WzKUqkq4P1a8A0z/RygAL2M95QCHhpW2IdOVcm
xaFsaPY5eNnDBPx2cx/uzKqR4779NEZhZv80fFUpLDxK1kxbx2Tg9VDyAjz8+YtdV87Pe1EvTNcv
1XxqAFx+/ZiEm7GmpD5BMB6vjOqNAs2/R1zzzbcUlLCLMj9gjvKgt93RCbDOjRfmtR5KWQLRnd1o
YsMN5z0JbgsVGH53zvqH/BIQtkPTcAHjevF/9e61DivOVpStLVGaQVuexjsmrpHJ0of6ITgT8DyK
xvRm747F2nGnGJjmxRgrN5jb5ohrZB7lQgvs4rYxDq600W5cPRkl2ZxoQM8UZf7kHmlFOACse+Qi
KhKX0+xJtgUqXWS7lyaDqerOEBnmZGj2YUEpUZnXMHXkaqC0gI7avdxHZmuvbQCDFvV08BgMm6Tu
84psH9ocBMvdj2Fza4NTuyf9IASwuijw68G37LxWaON9rAD90DUHKkua2Fc1n5CyEmYI27ONCT5h
ieckVRdxkSWP1yZ6ycbNAAv/+xDGEpXZU5+ooOBiCk+WohpzaZTDplgpAgKmaKbVtDRUrhs9KKpM
ikhMBW4vIHoXV7iOYc8f3gzgfMJSyMKAfuBRLC+n2zRH3AiaDrPLpxfq8kGUAExuRN1ymXpgWdmr
i9VPlDMO3nPFaOIXoflOM18yHJ53Whxro1MzSU6t50Gxna7JpkQU5JdSbRH9H4ksxuwVhbY7LYzE
KupKseruda0nwUJPknuR8QeCiIrJQQNC/RyxqSvo0vhG4LU6YDURXgskwV+EIGYQuJsm8KcEJmx1
n11z1Pyou943UiE4Xi/EmALIwivLdnIXXoHsRaROY/coCVqx0oppG0PgD0vw4E2a3II3YhyHC4NB
ev4fksXysnjbZbg/FJKAsVpJZA4EUD/HjAuyRW4KDlOdji5jLbcinQThK7+yiR++Ew6sdW95VZdm
vXLyGbKRqOpSP2XkNMIXPv6tMPjzmMae1L4rQGdGSEV6LHE/f7j2nbnguo15Mmaa1iTTAYoU4zGn
RdtgqmKsWYGo6ZGaMAGHB3wn/hAAekn/GQk+nno3fLggMursA+Il0SgFS5dWIGWRBPruMTrDmjnR
iIKqYqpj/H4Kg0nCsMJXZyAPmKP06qWIcpZaqxQ9tWh/dzNR+8vUoWe8nT7J+0secEun5+twrdQL
CQjrJ9+qVmB63mLh/fWf1z/1FPOePqJ9SFY/5NpMTNAztXo3tDp0tADVsmeqQlUDbz/dREC4+oRn
1Hz3wL776zEtFsezoGRz4IufLhGa0MPOxPhBGwaiuhW5/BPhoUclEx0i8gKnPG+sI1wuY0/DPy2J
OeL+RR6zhtKKKTxN/xCsUEY31p15dViqLcMcArkJPgGDdGc6KaRrV9eERk2hiWR7TlOsj136+OH6
wy1KS08a8rGZ04AHucXhpDrGmvncn7raXUfhA2cJ+siZgKc233PJeZkcn7uaSmlGsSWG4VFR1lMu
apO8pZvOGS+iRbwMmtyWM9ihXMeBpoFLNpenwGD5/Hfd5oBkBwiZ2RUJ8J43TikvIvTjomT5dZFF
aZcOUPbjDWB9RiqYlL1ZItvNOTtDxyF55HrARwK1da84rEpjHLn0o9jCSfgbgTCqc7xB0oNurgNl
+qY/Kdt0B3gUECmETt4B2bjh27uZ4RVoEcjoLEe1GtpvrG2LgHH+cMGL0ThnXTp4MwCVnQ3153hT
fsY0cZ7vjHh5bEks7g44B3BDhg/aPDSr/Sd8NaTrv0HOGDM4dYL7UBGhKH/t9E5Hu+X8QDBQh0tI
HUGrpKvZrVUJtLc6mhsVhzP5h2Gv4XHCz+wil+M+ZGTins8ooftiax5kQ++QMfeFZzAf8Iom2Wlm
XTxY1w1Y9J0+QUFA5O/Vt0n84727hmpO+7QFG4UL/Q0R218uBk38Ka6s7GzThQXpDFMIbJDR5RqE
PE6wAKBOIOWRWO7sbJcauzOp5VfS+GvIhyWlOhsz7fqYbWPsxcuaIK1IYwC4gzpyPDmJY/BA5HmZ
HYjJGmjcFQw/wHMA7vREi2MNJYlwYgf+FSkMo4rNNxgQGSFeqCI8kdp6TmhTIkMUTHamFy7uSa6Z
c1Z14dJutG2qPXkGUM9+1bMkmG2x/rkiJqI1+aa8B0G1sv+ISmxdzeNxpaELPRpIr/8ys++Egjbz
gOBkdsK2UDnJxtjEXPf6+aox14wn8GLgmbbrOxRxgLyOB++5PqZBwCbC8RFHyj4G5H81H2QEQ+01
3cTH3gcOIf91Dg/ba4dtX8OlKZ2EWYOUxlGnm94I9TirZwPIJrrprSky6h1CAmqDAc7I6geI0B2s
tTa5MZv3w2V6BgFvVdJcupif+A+lZgdrx2NpE6vtfjBV2I/Pe16D6CeQeR0/qXrNSQ7ZG4GE0mzu
sGWDj17c66+i8yvneEIggN+7v8dspILrTmPK2WXk3KgEkQNsYFlWFFsXfry7UOtPDttQrn8Ln8mv
kgL4xvmR/i0nKCzmVBA9BQKYKzxJps9GzRkcyVsMBPXnbvFrede7t3kIeqRPilzuaNTy/T4MEj4F
WoWlDBplB0dp913MsqceWX+no5w8lFj1feM+7kRaaTDyg+B15UExctS2sx9C/NcXOlJR1Utx27nc
mwshM9LoUncwLDe+OXD+xXrPSl4Yehp+Fmx8KzcCZ7YAkgeC3EEXbqJ/53cYehCmxwlUZunLtSpq
nPpZdQpYUgSxrwaifaYfyBl9K5a6SikkIbH5JPAKebV0sllvyIYG3HVSg7iRQPqk1UNRDovf3IWz
JlPj57OIw1Iz6TKvxjb7Sx5buFaRGVkGUCoDNjujHRPrikT0O7qnjfeM7QghtFR4fEhRbCIyyc7S
6yfzwub+kdkMBbMWsF8a9eFv3jVerVkGcLKlEXpiaaf54RiQb2o828uVLnM+zqr/G1gvH4lPwbHW
oa2cVX4CYSrA9lAZsuj42ynnROKNVfjAbb8pswqRJ5hZpHFFRLh+7Qlw9b0Q6K4Ro25pDAlCWbyY
kbVKC4wBC3hgh2OZQ28lucA0zXp9+h5xaMCpD0OlXRzfWEdBB8DQJXZ2efQoOqTYLJcUDBANZYr8
icmg/X3dug0pI1XGUBQ0RWXU+X5L4ov4A3uU/WbCKTI2u6j7d9XoFkzBqvGKiI8/eAg1r01Ehks5
NRTNlNK1Y07v183RMC+JZpbaGwxjq7qYn9EvOg96VxN6lLTM6vf6YmElfxfE6MSr9HA3quNrRO+C
TJZ0YoboNaVi8Q+X59G82lTOmuosxNgnKefHnjzTdXFhF7+sJxZOX4SmmVH6MrhNRQL86wswZMs/
6OHN3rAmbbNwgDzauHicPglrWUX5XOi2xHCCmFsX/eDIRTNCxtCEnkTVdTg5hIPR1pFXikMg1yWn
sfqRaQESDU05TyStLRVikNERmF0RlVN7+7KMWy3RT6jqg5sRGDbDShuydujbnf6CZFCxvkXM1Fsa
1tZyeguVsjl8Wz7PQmbm84qGiTtuYXx5TLmGMevJcJlrNZi4wkYY37jdZzKkJhr9shBAz0WlguGg
ea6qkMs5j5q4dBzOUGaf6HDGrR30/2N5n6Bmr8vtxIFzxIZzTIdF6gGznDE0CbybkxTdcWH42ksz
mhZg6Rvtv911gjv+LkEyXBuPoXhRV3LeYwiIjr6tq5AXJjGBF7BAAie3oy7Dmd8lx9/EAACMOFiu
fBgWrF0leORFc9WPml+nR9NeBbdVsILTsC+i4/Y2Q7hiF0RUWW/0ZqdCEeRaOtB9ZoyHdPZR5Iq4
ZLJ1oXwNMO5YZo5aH4s8eVxqtvxWeOgGhdSZTAbbWy3fSnuUzgnuz5Lysm5BBgj3FlhwUIao6Hi+
9dC5lNDKRczzp5oWvbSCeVZUCG2GkLcG6GSPnta3P2agfUf87gzBmE3TDLyEfreCfLzx3SBChJC5
tTzTdNzBE7CWiyUj8r7HfMDVu18SuAFYbLUREuhxrwrVvC25mFXpO2BbaE9kVtqZkbI1kVAdncwJ
fzXDXgDk9cgM5+Zdq3XYHukb5aKoY4S0x2Q1O3y3EyZYr8jOs8DC6u2sSyrzc9293d/QPGUc148Q
/JS06JwPE2TyO5VTFMqyKmmbt8Qh4ygvUeThW9WPcdxS89ZEm30urclG235NRVAN84FKqrbbznYy
kh/9cGKsdIDWhqJ7MAHgBAA3JRWKDv+7GlqxWx0HuU0LFVLr8f/hlBxCQMCrzc6PiUtvoey4Qbo2
7wDy/eT6IGqKMyDkAUVmZmR8QfXa2DqSBfFqUKsiqkQDx0GQOWdL/qMTB5NOQQzRRGAvSCxX9M4R
hfwXoChxUu5IqZfLm73ur1GegIphRBbcs31yN1V4b4xGVtuL6zUYm68JJlYU3XtmXlem0t6qcJ3D
ivnMd6hxgcAdymifpHo9BRIgS58GPJKLuq+7pypIZd689+KBO9gw8bEIWuJieepTTFSfTnZAGHGn
JK9G74xHb7sGi9fQ4uyS7jcFTWMCg4Wwx2N3dANurjke50PLnvsLDWYFhR21PmPSulMZ/raN6j40
xJcoyK4nlk+gd6HYmW0UYO/f67ebG71tChVrDQQtY0avYVoqD8B+L21umkRICk1R9C7MITkpn22D
rcKfxEIPqH48tI/sRHfAW4VP2mg6LM1vE9B0AMpBm/NZgDwD5Tus+9GhEJ6owfWnNqsq2Rof6B5U
ie2Sdu+p91Wg12FoPNN5sgNmF9lRS+t4U8CVWFvKejOg7GdB787eLUFT6ZX65a2TJJq63Igampkh
uBS7MvkGrrhmKBK5sAtmDiJUO8TPmpC0ZvMp311mcQsmg612UN1CWdiIBfFB/o/o7iPc25R/f+nP
kSbRim1d/AfzrFlpYGH5hmbdXXSjnMACUlo335rVsg4Rj6AV6VFTR7kuFQe3uW5j8oO91wukc2SR
8YYZgpLxnQVKiZ/+Y1lDOjdzxS0vmDaYxKQP6dm1ZgxL+21kyNguHcvApfB7WQBLGbPXG/g9ooTg
iHS/Wjer05gxd/vUJDW8/c6C5OuO/QGt8cm5UbLkJrNj/6ek26g/XwB9lUmWfHHYeiWztK5Sj9Nf
sk55L0wZZwsiO8wMEFp7NQDBVAfcCJMuJI8+gpH2antXSJA4+IwP/rX8xRWu4JoRfO6xfGB4l78X
hnGcr/Dqi+gsSPmSmB4to5n1VuYmpCoRfi9xh/2DdrYTFJ4yoNGspY2RInfR45MhLK0Qr0Kapzi/
J79q1X8cIeFE76NL8/Sj8wTgG7K2b1QY3sb7GasZC1qw8ko0YAf/BJvuLJpHrCxDiYhhbfVFoVzW
pCXA0bvrnraTip4eGJwP3mhsZnvBj4aq+I5yBUACw6QsCSnVVL06elj5PnGMotax391gFWcFIS1V
Fd6WEKEjK11byO5VqqejGIN8WbpbZlqIGZ7u1NJdztQrVn1noG+lkYO9mzu+yOjRoc8PVDeCSGpC
PbKBiTV7BsOxw4P2wr8uEZe88M1BZ0aqPtdYcBQnVJ7XPUSxNfMK8Dc6kiwN8uZnjNIAY89fIyXZ
BLZcQQ39O0A8vrgi8/q368OF0X5KEHVDQ8pgX0gNu2tilCicMPkPAQGP+GU7xJ/si1EzJ5WNME67
jH0Ut4rWaR0BNz27KLk1MZXnw1F+dYnnEp79PSj0knKgVErAEGkZiSlA8IvNEfICVhVA+aMx3MkB
BguanziiCdhv29e/V4TJeuGwRb6dKx4qs+VEgWIRFXuziptcFpTuHbrSFGLiTfmUAMbwYGZiNRvY
D31CCkmcElU7f2Tm7TQzVTz73zwCpOi//2kjeVBzXdrbtOHFGSlYBChE09zSWBEY6KmyueEnD7+J
gdThfU37DyDwSmHpEZ7sRQ36xvbzT1702jdW8I+GZVd+RMJEG/G65twVpwyBukKhuQusaQTqjcuQ
Oib7DJV7gb34Q292Auz7d2s8pXVhF+r476AzKh+9b0c++hJrFWHE0WjiLAUZ2sT1tMYPSCiGqZUU
H00e8bq/WRilog8gJpxXCIlXKUUKRd7Jd0+6DNUhfoz410ZKEUZLXBfaW1Qco5FP2jqb/bNBjGqz
0DXOzt6BHSizAR5ZqXyubA/04zjceMQJ1V5UbINIiOlkgkQQnoTUM2WBBAuyQbOf+iWLypvY0mni
CqB0kS2HZGNSiMzNrDdACiSBdJdR86adtqJwojObUIEAMk3JmOuXhjaQOVZufkobyO1loZkCOUse
82IiCdSZSOI09aDet1XgsAMZ3+wa43z78d85osOhocUhy96k3BIRW4hRsu0A5ZGbWFPP1TXiEg3R
gVnxBsUZ6UrBqF9xQyj3PradPhXHXxCTx+9zAHVGxmKRB4khCCpixMQs6H0q4csTzZvpFKulhtZK
sCtJkoitiqsA5A/BNGmzwPX2vFkfveCfpnnI1v4cNlNvY1DtPVzeRXE0mmlmmwMS0KgMjVbirB2z
oNBoALZOjs+/RFZWOwzslSpTBuJoNcC2NtoCeq8by+kCZK9OemIcGzR4SMKpWhFdXkT12eQ7/kpJ
pD3aig+4V7o9AfBnUINfQqVzADdHNIQYx5Fot7d/vXxEHadRXWhnJOVYWNDJOD4qciEL6bLEWcAJ
p7ZAM1P/btTFoTIFyQdyiWkgnWNoS3M7z+r5+uwVLYcV01KxmRzLCJ/ZYoe0GG+GB9vvIUQ5WGXR
YE7hoQwMm4mjbTuk6krQ/y+G8D9bvfJ+8jxwvQUXXKhTqCZKYPKpDfUr8HL8jQoFP76+jB/Hd+/E
1Y+QXywMcYuoMzbnQPwfqJ6OuWnxoMOxgOEfqGNmOjHbaS2dsbriy045h6q23w9b2ze1GQENsuuu
lg71GMVEhn3ZtQpmFZDT/btwE4wxOX7lSAiEoZ7+aH9Oh8MUyEnri5OrPIRROZ+Vbp3XXWdfGhc8
43gntDHWMCMJ9EMYqSwm/NcdiCwUpwkfjCdGfpqZ8AIPxG2a1Fa32hVKzKWNVkU5clpcqnVVgP3l
ScZ7qWQtVqSC6yQyjxf0cZI1P84Mm+UujUQ2sbkKwRRtpIot9H8+Ggd/RjyL1N3GWNxA/RcdBVda
UVvEHrNRXnyQcqEv7wMoY586ij7T6WxwV0fDIe5yycYQ54Xz4/rbeOPPxCpum/qiP4X3uNPx5fh8
GTOYWxTgZKSWTIn7s2A9E/H8cfmY+xIudqunZulOANdsi8NYaRptJGKqcayueVdZJApDf+7xs7hr
jte5yFyoUOL6iJA/kHsecECYMBTlvTIO8/5haqyXj/U071TqT+pJe+qTbaqbpGxhXEHVjb3TL7wy
WI1J4lxUMsehjFeAuKHfLwVNNO5Ix6Qe+DxgzgRaEs0NEw5KrfzoqfjSMuO3JmbeNz76vwaeg7PE
HlZAjQUXfjPCu6P5jjR1Lm8+Lsa/hEdrhi9d8CsFI/Ge82tfWsOrdBC2MLe7v8WMLpZ/j+/TRwNY
xmWqpqToNhJItDfUazOvt5P58/3ZiuOfPm8IV6l++PYTiC66VVia1w2+774X2CgJE8g7SG3ozo2m
qoZbA0UeZ/IG3EIdCOZ8fhhDLEXy9eCrvGRThSO8B3GTxVotXhixW0EF6GEbxay0SXwRlt+TviJi
hMyHv+4HZ9n5x/HJ7WDYVj+jAjPty1N/lDAVeXpoMS19RvxndwjvCv2gVXpf4iWnUo8CR7mBSSYN
1ft/SzmvO+fUNm+bvd0T1l4RFvD9F0INZhAIrmWxHb4G5SZtBuXYOVK7euyjrIRAAvJLlMtXTYuz
z9QMqG77XgNMjlUU4ch/jgP/RgKxI/SDlef/TL7wkSoHa4nsLxsJSH/BgznYV1VrAUj/T/0ZjQUa
YtdWs/5mmAh0+mN1yVAl4fCK+m01AHrfX2/2ed0Lb/op1VJXkTK8oq1N7SZI/2PsK41HG+Mh11Bx
pyXI4McTD8VqXmIj+s9lQFUNpcbXtjbvX9hIEZ1H3LcgjtOw7joZ7TKN0b2d2YyTdsLgCKY0ZO+o
i/9MAxiKYXm5w+W7wFshI34naHpKU4P4fItGjVAdxK5hNSnxwAvCoVpNM7xtcPZ17y4XVunIkFSL
z8pteuXiBUpG/r1tMBhFj+WGBrgHXixrmW2A7Ikpbj8wgutDInmwenJbbyNw47+Vb9Gpjywt7Nlf
2/qMzC99fOIDioTsjYTXsjXRWnpQ7UqZ6dETz9ZjZSJkLaqfZsdxb1Z9FEL4lsw/F0CSjepo9V0O
rFVfbe/50V9F3LheyxCHpq+MCVluxWzKyQ8wu2LGFDcplCnaP46jj+07dKZF+RQvy7igt6tfhuTt
wFo7uVWtCVJRv2nd1M450mgA4uBp/cLyH5Tmd0TvCA4qfnyL3inaBJiZk/IJ5jzAtTXi1BtdEmWi
/X50Gxf4rKsJSP+8ToLU7SNAisZYLb7W4fdfyDvJ2pnbu1zhwez8MRNEPsyDBdhxcXUoMsKmWIQO
tMOaEhaAndYcltUjMPDbrrbE6Ko8PvlYXw9jHo3kH0HgBHe6oJQSoUwg5TJXkao1xLYmMPJxmOPN
5zrYGB41Q3Bv8ERdQe5gtzmFO7viv2sYize7iJsFM9yt6QDnDbjxI7mzmrT3BqvQmpw1vUgnK3p3
1mWsTKvx92ta+34E65xX3GYqsVsN3eqbqDKmbuocGHzAj4SH5NVyqwaj/JKEz1xnOXUT344XsiWu
Xngm+JK/UxUt0hLbY6smbIYRW0JT79gRpCrFaUfs3CKCBqqUuoCj+o0BVktkt4VzZ++lANCN4abs
mFJ2UppfzbDhGbploGg37eRp+bTdfPb6pwLeU2VVTr20e1bAdVVK2RcqJAh7L3YfhfiwXBJWMaAY
pZe2vgC50MEgy5qeumiZIvpJngrqN0rJNkgfLuAywZOehtczlXG+oY4Lg+7rVuJ8gQZ0wSgvfWc9
iJMJ4oy2fnmWM/eN28fr2xJCB/XLLavM9+pyKaxf+11IFx7e38vQqdxeZVtnuC+HqVkjCShWomW2
mjPX9jZAHhsDD7iiFtcQ88MQUPMXbH45OtBt7KAwmdkfmqytuy8ahOGCPD8t0srhaRscULWMR9lF
qVLHHd6bmI24B0FKIQ/fmxyTMfAzaQVRBYgsB/XLTUC5WB7UiDeD2AhamdqTlAUSjta2Bm1PbEL+
HF5quRvZ/DTzyOw0GLWN7/QazAD+mtnjQsnlc2oEaJUu2T8oQeInVmO9Pt/o8jWCODUWDsqYeNhZ
cZwdjhVtW5rEumT7V+EjARW/UiuRD03DXxCEHBsDkIrQGhurSLeKCG1xEv/CeoilMoTIiGu8kiWR
i2A9rcSUFI7wr0XzdLMTSbcJCbtc54gdKVQ7ewwFTOazHGoft6QRqggiBPUAHMgvISi5B972gT80
Az7ZPW3JM07O2wp/jsE/lZqjNuCxaxCtqQgnZBKeLbMDvu/5ktWnvkZZvE0DL/3kEJ/Lvbqw6OCh
kdgJg9ME2KO3wnYu00dOcqF93hl3REgESc5mBwi+xGnHsnDD96OFKm9vcKux3tssFyG1NQrLDOky
o4IjRGkF3dJb+yqtxK1kgmaaQL5UXWdtl7A4bcTyxzA4dKUlJrptHydFB2k6bgFpD/Ld8PKg0Amr
sBNvhMeXmM/EwY2UZs+vv9XE8gigyNlaUFDccICR6PPxiWzebo8srFwEWq3cZoO++EBWPBLbuH8L
kMlsKw0tWWovUV1f0LpqVU3CS3zJBE0PX1aebQaBif7hqW9T6wxrMfzh4bf3GXyZ6UPktuCFnj40
pnpI2ywx8UPnBFT5kfDGmUVHZJ8QmOvgtGslco5XRpHB8wx3XMoOULsKFUjicQyGJfg7B3a6UFOL
uyvTSMkGD84loQtIWszX6WHORl1HUcX6CP6RYExHj0jbRXMXcuMXTvuTQ8AvXJvYiDI9qT9aODXg
3xmhENrwspnLVjpw66BYnWqM5XAesYKS4D7ABKcVuzTLteuFfGhBJnSYA6Ii9FVJQUL6t4suDjQu
YxUqW/EJeTI+eNeCFo6+x2VOEMN0Jo2fzv+KTQ/TDjINIvnFErjMLtJjdDY34KjoClafl9eiSe3h
r2JPq7TnLU7VSKeVtWf3l+QFNQXv0wtEc9Qirv8qv7LguHLiPQzKATJwmIyUOwNaJlUZRok5J1kf
4nKu7/JEHsfH83cW0sdpLltsOjG4GmxqcEtb9Ib8qCQKNy7sC8vGrWY/tZ5Kviydx/uEMU9qdaNF
lEKMSUbtPoGY0ncamNZEUlBR+QMlrYnLWKtWo0oqXteylw0x3j167UO3we1toQsr9p+AuROgFJEN
iB3pMFxp7AbsElA1pwIHj5rBDReinhPh4Z9qlw9/Z3B2jREQfRfJOP5dXw1vf9DG73HnjTDX8IOZ
t6gFH9MxIQCF9S8RzSpp3zdRkCJwt1kDrABWnpoPiyVroxa+DFRzb2Ag+nS9oYCWq+2vLs27P2TR
gOKeXbZY1SRCNq3cSmu9hU2bj3/6N7cKkQTBQt9MAu56RpfX9OHVi6s41sXkB0bl/QAavw/wjV3a
B2p4zt1lZoHQ7XhGMGDeWuTu+qGrz4jeCohATE49Aa4yPbYLadvhauX2EB/wshN/3yT7bsUUqiIa
P++lW94bDDnvbI3ES0FZ4UrflIw1rOe7N3lxvT+OXzIGMQOFOWlriR8khRhv7x60m0HMvajO0bAX
GQ94QucHn0MnOx+lIQhek7GGzPDoRorSdCRwPRIFcIynvyJgx+DJ2fTNtnE5UP/E0ShAEcQFkhVx
JhgrE/n9/LPyhi5WTr5LtkrmZF12587nJ9sF9u3aEB1fkTTKxFVIK3T9QtP3abn/oAhUFgIeu4OU
tUEr1uQ9Qvi1l96f0RQjBtn/eNrc2OFtHEvpECNiyEXfnsT7Cop2C/+K0PNDZw31JGPa48Q0dsZb
/Gk4SAqZ8epeyDzvhv0t90B43NjYW8KHPmfmNzQcoPb9s7ifyBH1XtUVhQnFsfjWKA/J8gLqG9vZ
hZh3WaP3Nle6mzXMJLeBsPF2qr97lt/2gE55kCWTlmEcAsXHiLmvFema8jrFyITF5vYI6OJWj41F
os8L2vp8QB4GNBsY4CXXVV2omiMkzVS8B6gY+Uf03jOjnc4s6R2zBldb63eF4a54v69wMO/MV2Xv
fud/RNViynLllPLH3Gsv0f5tVQgN4cthnB2ALY9q+P9tajW68VqzIHiYmbnGyKZRAIk8OOyAKnzi
ZqgdjgDgIbHrX/wljlO1jvjS6+h+/Ik7TU0aicoQ65XP8hYnW14TzvqjQmzm4Sg3QaKmASGypSLU
hIqBZIg7B/XxkUrm5uCrprlQFHKSJ/WYb/jw2erWRIjy0ULmeBw8n9dxRPIDNwvnH9sbhObM1ONY
bPHXGEabDNoE3b9jH3tw+dXWM/fSEnuYn87IFgkfgqjaW1od7gsTEL+oLaA+c3CGDZuAImj0xt2O
hCkDpApFEHXiX89pARfWjUBw51LdaQ63ynO/F/gBUBIcJH+Vyx3TR0TwU1AgIJLl4E7EBesLkonP
OLuXSk6xQz9YgnSURFx8ai6LGUgFCzvg/NhqQVLBPxrfwkFimCskPcM07WElobv792m9SiEdEJ69
daGAzRvFNlmVyBvBSlWfPhkAoMpTXAgLOgtcevDrDEnsCtB6EzFSyhbZr//o1VkVAHtTQfC6dykF
DtKpR1Igq4NffWuyrfJ2XN27wtaRmdAooINyd4y5PCCo6eqLvNLO1OZdNheVHg/AkL6xIc/Jkqd0
7+G2QJzrXcJ77R9MbRSec+3qtDjOck5vbFUhChSvi5dAg+v5Yr5kuf+AUgMQHnY0zDg5JlsfGHKa
XDsCVHDUP3DD804A7qkgys2QROWD2BIerK2iilClwj5ICHO/jfrSB/xQw152NiX94Xy/pZ7UG7T4
WMstqUjgiy4+zRC0FAS87PiVwf1lqzwR6GrWLsIOgsIp97qPYFyDp6WeOUUG4EwbuhehaLppchbi
bwB/4Fd9RngJW4BMdOwrDp72nx5HGuY1uE8kT3lGZZadeh/AyGQRbGlYdOq6EhJ+VTwxA+m+fWD5
82RLcrwni2Pg8MwG25U12Kql308rChxkLcctguD1KZXDb4UYawqCv+sdCTXRL1eKmSD95M9ObPPA
aJrcWttehZIsOYDJ/E9zRaScLwQ9aRJRQUrNyVdcsXB5ed6g6ZMBlbmsz1L42YmP79vycRt9W4ln
LGJtDEG/5yjjDUbPZU4wwtXbKD6/gwNntl/ft2HvZKrEUM4LVTOzaiRp2WpvNm8k+5s1Fknw862h
zk6NaZV8tBzfynRZWWE7SiFQsQUI8dMwQpsRaRbchP3j2O2FhLCKMa95azVlN4rtTVZqibuK/Tb8
DlD0QKdMRBIXQX36ddICrv3vMsZaKgSZk67bnm3kQbY6xp3XwKUv7Y0ScyesmyTrbS5ciYqKCOM2
aMib7KKTXbs3Sb2RtOoYQSajdNBSE4Y209ycSlUCLLwJkLqtiOSssLoPGMXme2/g/Eg7M87e5u3k
EHwsEY2atQ8lEZm7z4RjGVKLbVxsK+dDSvwt9MlPHGGfjXYrItuYJ/7sw1IfuzgllyoONqbx7/iX
y1fE16l6QF5FkenfFREzcsgWXo0AIMrzkIULd1Wup/DX+XM0SfBpAiidMfsb5wo5KOMlqfjvXFuc
AicEmees74DMRp15+mV+/xW9m97MbOTvOafV5fNLesfPf5PmizNhlIPjYb8LWtmwtY3FUAcprGfW
Y0lST4lI5QX2IGjUkSGTVpELK8JMpyvLveKL0tzIWE2oNPR2R11h5lV7B3c0hDwCqlMcCFUzJhG5
uEConN5+utxBSklAN4z+3KTg2BG+QDNsuLdGm/S6/4jELSRPzKYq5KHSrd+0LnSl5M1fRaRKoA6P
NibGRM41ArcfRt3Nf7XwozGC4iMjHHlg8b+l053CF+v9B7svB5SJKuzPZx0PyRl2+2TOFL4g6wRM
aFDMuk+xq9kLoTYtvTo8nXTu/ruzioMow6pFSS9NRolnqNhKnarf3trZRCyZI7bSg75TvULHeQnp
yyZ3wUXkTgr9/9Rks5hncjGnvIPC0ATaistxiu+6+8OUWrqHys8GXK2RNYjhAfdnpBi3k9jb8jmi
rkwjRKAOBFjlgWUm15op8tsOG/Bi6vFxt2Qghoz5HdnOh/MRTEVsmncv9wto3dEB7F1fJZfUM2vj
eawDNy817i8WyAunc3kqsABLl4Y6THmgqOCERqgEHAOoth1Zb+tmuP2hJYb5jqElYe9m7+FUJORX
6gIg7F2KEVdEU1cKj9Vkn2qZR+3dvJQBXIvhsbMrBXEg508n9astrZMWs99W++Pia6S6CdEgvGNd
v3nFAbXV6/vfY39nlNaIzB8NCgDbF47jmLfGCulCAh0tgBhKkj5x4yOqYEW5J99LrdJrKBkzZKTm
1KDLLXZ+QNcvtsXHyv2Ya67pkNEQS1cRZbUHivKQZDl8s4gnVAXMHkZsQpnjbbg2S92x3lIRMEFQ
nD5rtTmzqVJPdZOoc8+hITmNglCZza8SBTUqMbnZEQ3hJ1XYlerX9+ukCM2dQidWZu5XhmJFZzmk
9qNEqnSGBhmaZKMjT+LvMtgvWBO4JOAFdw9uyhUeZq60mif5p575MCM5egEyGA99mO8kOBiu80Id
TTn19hi4gRWua1qvoqCknUJb3f/t+0zc4Xa50pX99fZHmOa+pNNra1E0nVqtvjNvoNVip9Gfl1yG
qjeqOQ5jtBR/fUXrB9RstFLYvN0IpSUqEanqQuZXesCTANdQDqfATHpdQuv5YDSaiTem+sQ+0iVL
vohZf9hnX/QMNLRmzj5JpKRn9ksz7Hv97yEVNRBttop1HEv4l7U80GeP8sH0/gKMQlZNqLqs25u/
PJ7Ny2uFB3Cq56+zbkIqLTu2BhH3IKLPRIzRzQySeUuO6J30OcyCtVTJMjXuFddv7/jXhaY9h64Z
bwti+akBQneZKifiiJXpBhxsE0fUd770BVAnNWvvHsjLZzUO73IrcyaudWNjqCW4iO3PGnBaeKe9
MdUj2BZI/dlQowNlD0yg8x3FJ3eCKzo+zC9odU7GuA6yvqVAYMWKjLGNKCoBEZYjOYy1cAiHO1RU
tBWGRYZjXZWfPjRWbHcP+5vaDqlpaurq14Bgpd3mAxbX8fqJb9rkKBUZkpv8qGvzWqMA7xBQ9Od/
lnJsMefGkEn+DalI76hYbAb31LoBd2MMgTAqwbUbN/x6s+RjvR889X/SecHbAFkGjypVIOCG5+MG
MG/KVDjzuHUB+CQ4lWGI/N5RxGIUhUMinMrq+IRTgGgtciHtvQgRgnHGGUHM5fDcycjkTgmeIwD4
4eGqjG4Qr1hAi2jfq4rXYRkZtmULXWs4kTI7UlBY0e1STRtwjaDQMLqQtvpmWmKq97qIoD8Kd0WX
80x0SQGEy0SCuvlTERBaePSpGRSzXaLARHVLxANDldWaHL+HnNRkEDQbhJjDetdtEMXU1yQDXDGv
caDdc3Ea4ek6JAed6huOvHyHNvzAF3DF/X+4WsZKk//G0HMfheIqW2uxDX43ybUPFUQ+VyrYcal5
ZgGvpixgvMxR8UGMw9GjJItgCI8gPAZp63frHIjmJSS4QyMKVc+Vx40Am+dHtS4PIPpn9Xi6e4at
+lRerYSUygZEBUPgsuzm35z5cMs7oB6TJ3k4n4NdUhy9yPa4wIcdXIre17vGISN3HOvV1ykvZiAP
kzeHiAi1qPNU8VRedbcHfhMZMXzqjuAFEhmwZ+IZ5HHgg4dp3Q9BqPsrBne9u1mm71p0gWF5fQJN
KQYsihcEJ0oPgDBSmi7pM3fDyY55oLJnCXm/KJ8aZusAQVwb/Ftm9GGbjtyVgCTjBSKc7LR97QJ0
Kuq1YNxzEn4+/AKD/Wj1vKh06/Rm7+i5pX6hFHCl4Q5YxSDtq85FXsjVuQRCwC2t/YZ4Uf8OOr3W
S5QC4EXxe3q4QM+GG0Ts8zP7od3jqzTchlfyTuroywf6Ac45j2hPsaybMdAKL7JBmFNZ1h75+zWd
7LUgqa9X7QWWouO3UXAh9itILm+/uOwsGDNQW+V11mW50BYecyME4lsvincr9p2SwH34UkpLYEz8
RD5CC1Ti+/7OIpAmzPi0vtq2BfEgVulETPECq61i0Ee8pbbFf4YhWBtX0tsC+mjwe64F3Zq5ZgQr
wHx+TNFzYZzSHoIcHbdgHdcws+SY4lAsY7dE5OZQ7QTGWASgmhRk+LYBMOwe97yUT4iZi3iDfX2r
myBTA1gH3nq0Pafwt3J4dPYHAGVSofkr51lOjkLZpynoQgZW0c2vuKjhbY+ByDKlCfameWSXqJ3r
V5W8YVEtwftJV8HLB2vZCW/p5Y8g2StYhsQLYTyRbfNLc8lP1x5kGlqvEeLJLKHCJlsVt8oyiLQa
ViUDdjyIORrnDccIeArNxvZYX3bG89wUE25sLG9FNQk1jdwRxElJp8wdhqZvpjbPvlVY1euV2iM6
YWPEYhCaVxh07NfM3VLsBhos7q4Rx9MTirEVGpz5d6zxa92luJkgGasDiFQ2zG5vZO50c4ciHfwc
noz/Wcapu72/ysdrtUEuPmF14wkuBrElcExIQ1x9jhAN0OYkFaeDTxsrjP2gv0aFLi0qW9oGVeqa
lfzngKkOwX0X7OXiiYhKgcjcers+4T0rvUkEud7ds+wXxopiNK/eYZYaCsLNkhzsszG0eaziNpXO
29mEOUC9lvjWVQcXeU3pUZ2RWiJacN81GDmLvkFi/nhaQkKc54CozEMLTebBRVytZnLVX+a/JRuS
e5pN1ypUiHi0Hl54EP6UvY8j/b1LwN+ZYv2QYhr8hEwXFm7/flRNnLyxo4OHkeGxejd17Lr7P319
3gHQdMPF91hOD9oTFzpcYRn+ADH0fQkmkMZjHHgp8LGxlYhVd/0taA7DKV4NkAoWHYAjGYeqBm04
jLUGNbrrkOJfvZJ8QJyoptJKWoS3BElJ8oeqqAo2T7ZdoeTxFaPqgLh2LwF3GGanwBFVoaNuPWKk
dIz7FJeegxatHAxtiM9psSW6DwCJocNCKA9HGaHBbokmGTrk/+gVe6UkrL0qEMZ8BAD56aTSvItO
Z3phg9aMQ3Ey009rIDVer4cItfeusBxCxNt3P2NquGkjS8TlBbFM/3eKtDdDYEblSpfdkyyOtQkZ
cOOcj6OLWqlEO40cKWjGLMZIDn8//E2usbHyVK67Jxfu4ndWMaSP61Tto3qbnoFeKxCzX1yisswy
hH19VWUmwtBKTyAQkr2RH+/Go5XqH9RaN5CfNDW7a5saZOM2XL0VuYTbht8XkvOpRTFTb00QDSoA
jrW35WZ33KTb9O4q4TIFVTo9sUOYGt4hdULbjb6q22DFqvNR+fX42u5FQQM0lW7ekJXXZ4M4E2Kj
5gKAwhM95/fQaNWdHGqCq6RQqounmmNIKqNS1dWgWFHW6AcCEUmXhIil55Czd0JJIxuUxMbXsMtm
nu/nY0g2Rc3Tdqi+3145Jlkq9yTtTQDfsemNOHA/23y7hboZuSF4ZijEE7J80NymJ3/HdxfjIIK0
f//dSKgkPBcqLfVbZZE189M2YMo5npvFiDo64cbeIPGM8TBW9KwbGsW3ooVU8IHn6cYKWEIXd1Qn
bpa8aLoayiVZAaE8VH6XFdpHls2Ap0mG5U5H9cpi0flz7/mNKrZvDjowQbbtbF+vcTy+66Qqo3Iv
/osCr1ngYRkbYVjDWCnyl25pvcyIJFUT+lkWwrfwpMrXFzONPoL6f9/KzO+3Xl9VX0AUJoxPHmMV
HgO+52qJQA5rgukP8jbNevyNi0Gi7aytrTisuXxms8UtP6c1sZsD4uc9JCxrbxWEh3p8u1gqEwWN
gVCzYj9j1ozYqFyVuFl1N5pl5QPQb5Qe2krq+lQLPVCY+ol4wNdpRqA/6U8cYl8z2G44nMQocAhP
zKYPUXg+sj4X4ro7Mg9CO1jDQJeTNDH/BVPffpubrv8VYZRzX4sLrbofI8o0BcB/OTJBbuffb0Lp
TMWthdz+0mxNSm6/pfyKZeQDN9GgBjNHGWWBc/Vvd1Q47bB04PFXDh1+jgX8XFWXBdA2FuB7p1VM
pxTAOtEKGkLGYFgOkzja11JWHHR/yKaT1mhzIJzQW2YEUoXdjKunvXwApQbmPuy+MuWUTD5LbqVA
+cAUg0hoGrXY0RHo2639YVIqZPrX3lipDcaviFVFBFLmpEcqfPHkuJVkJXni3zHInWQjrG0Ei2Yo
NOa+w5EnYJtgH9Fe/HpfewIR26XJ1ioAdwkLQr407WOuKN6oWxnl+BteT5K56ph/6jsOBUf0zzIZ
xSkW9mPh1iik1NHwBVJ+lmowtrQqG1t6JcpG/7ojOt0baRrdtk0SDohazwcFM4F19j8xVF8ZBODO
6Tc6O5WacGiYrw3GA0XG7KnlurY1JOK8PBP24ffa/RVqNrEk1gjik1HcRQ8KybA2ZneA8E0xUiX+
i1ek/KneSrtE5gqqB5IhLNBh7uQW8+yOtprd8MVRC/tfgtjfKALkTlKq+WOZ+1GBj0iECWArmDiC
IENuQKcSGXDl9V1k/m1lAtSt045VDmxQHPZAkgmMxgJWmUsaZfI+9TdLPqml+xJfgmXU0sl2MbDF
eGDVe2gimuzADxNG42ChYpW9uj+VgMM5CVzSPhYExjvilZH6FpT/HYCsGsgobH3ORvGw+B5tEvsx
kzFVDQkt39R7iRm2F8guJq0Vch6D5hRFa7ZuUQOmrwmHMvPgRCUsXv+ZdIqOvZgPCy9gIz+8XIwb
V2d80qd52dNsiMspLJgwm8DZ35RX7h+wHNAfcz9Y3c0eUJaT1kchTW2xhS0zD+ywrHw6DkcyL0TU
8shuYMKT7NnCUGt2nRz7YYgflN6Eq7tYlGRnUDKgl9osWPai/8VxCTSk3rENoRXaPQowImWWG+cU
vnYI8JU8XxjlSm673gWVpWCvulYL+LCv4T9B2/KsqmYEw7xXWDAWDFGOF9m9RJd6LWwLjhTSfmBJ
AMOU48loNhg6pvN8sIRgrYaTSfEN0stDvyrEJjPqAl2xARkK3wQFLwWIsRkUg3pMlq6bt5hU8fkX
WQFe9tmZTxbwbtv/NPNR4XCKWLyYHTd+t5BdPWLG3BVA2Oy09TKFXUGeiA0BCdLvM2Eea7g8Um9X
usglGkyJIFZng57EUBypph4WRL05U4j7f5M9MvKKtvsC5h0o0O1SKEnBYbdr3A5WEPps0uP6xKoR
p5NGQhFFmO3rRNY6DILebpNQfo31t4VfhGhIi1w2XIkzByrsq6rdHg0nuaseqBEyKg6bPFeJ+7A1
uRavoZ09qZ6wVkDKI+ksW5EQuy6FOwwZ88nR+9e/w9wGm0TYrHmcCRuyRpLEgVPWSpHw6iERwl5X
d5eAwfwFpn7LsVF8k8XFu4tnLn9cD9EJhsJh6WvBHdDrct2sdZLxAopz50dAUMENCwcrmE7ujmRb
IdbFidDXG5N2N1QEnF96BWE0MKcb3w9ad7/huiKEv5eJh+tQJKE72g4iiE0z1K4//IyY4Y5GkdNn
OOxX6idg8Zu2elW5s8fqkkKMIYZwotnuYR2UxsyadLnVrOGUYjCpLxhxzQ6ZhLpCrZWcRE190ke0
XaoznfoL1oMtb0MY2yHU0WzeVZlkklK/VcNxhUcQxOt/CySXndtrSYC4O6HAF1wNrFU4POyaSVE/
bWQZl4srsAoxCOBxMYeX2BoVQebFYqne1YKQo76vdiNImJc3UYPx13syU7qdxweni3m3aO75aCAZ
rnxgy8Ny3CbZ/9i+fnuN+jS4kGMAFuxbT62XtGrCOBKQgRGN+mphVO6BtwGmWkKx2jml4jeTQhEC
eQjGZcrsp5MGJ48KA1VSIdQv0Ve8QpCUzbGAWhL3HrFDZ/3bptiRPgmBjojKRcXZha2lVq5tiUeM
Xzxr5x54ehyXzW/QjP7rSwoiN/4Id0Ge8qEIomKayWErfUAyomzJ2xeuOEnDLy9vCnU6xZrZ1qQ1
ZsK5N8sBjaP2WnuDgvq//kPnebLfC+3kG287LJ36jZjE5c9s17XAFg+w/ONjy4ZItJ98+IyWQOQs
HU03J34Ecg9NCRE78yTaQLshIsBUxZivn6WlLhVBiO2BTpU4mf8B5v+kfPR6UWXwBoXocy+ZdAkA
Ihlcsq3o9rPEoKbNvN2QyzAK5wXlG9s4rox1on++TIfsttwhuDLE+grd1nmBpqgre2JanLazMFtX
RZahqwkJiYUBVLqSvjtN1/BhWTD8jXXEKJaL89mkmyxwkwcs2h7d0KhUO6m+MEoYp9ET3KqFfeJ5
OI1JfYXjjvAdOzMiuQWGr08n3luTHuEdOZN6pRiq+qCCuSZCkX4hHpuxqm30dND+vG+FEldlRuTh
iy/E6XBfIM1at/JPXkyuNQGkaQ0SdVC0aEaMwaFssUoNaVK4LbCJ+YuMXVbjRmtj1XawKDjFaVF/
KVIhmtzOnMWeKS67x3l+FBmU7yaq33QrY9dkMkBQZjz+pcugtJm2Sk+u5/P78h4gPzhNY9sUtt8i
ihlINQjSiWoCN+VkCvn40NpNg7JcsL8jeX5/QCDnUbGY+SjeN1LlrVrSUnPR2evA+z/ZS/7yQVDk
Nlljf409l7PxOqnPG9uD52VIqL8fnrvwxZDeM4N3PVu8XN5Y07TsuZ+HsaprE3mSdnv1TsDf9yTp
1zfcsD0uMvChRs2ZcswvSEXeBJhWPLYQkk0RoFBmMkbwdqXjvkZWD9y5sCCYU2Ajz4yjr20u5Wxj
HxT67JsuUcFHFMtHdWNCQUVgsQmf5C8IVVLNKw7GHldgl14/C28ynECchxWeqtmHlw8ux6EGc/GD
fAPMswYpwJsvCP51gmt0Aria9oT/WT6deMgow6hxpBzLXw0Nk3UYXXIExBnk1XXCWeXGljQeHW/1
sMvYPXEvpri9RySnKnqvON3GBqkrS+G6pobTfaigPrHwOOZS5mePIpFQAUvEhLX/j5t+3SwkZcjK
Jz+UpbatCuIuq6CH9t+tmqrl847fljPewQkD5VTURDcy09VWC/C+Tkz82vp04Zt/iNckpTRzpPz7
ny+NWCNZ4m+FtafJj/gqi6RLo0LJFQ/lovx9jZxmJBi3y9ZR/WC6oeN2h8Z+Xwni6v6XFi8u3SK1
J4xEKkbB9SaLS1nFeW8E8N4h4bkTclD8AZuKB7aHJyjSIy+L5tBY210uonPxCVFauBE2DjqCvs7C
RZmhgMqGqyaFJD+2NEgQ/qFptm38gQRVmKw4f0P3Gi6O5+iInQT5UGGoH7xYP5AV487Lmu5ShEby
syC9xOyC4UBNuHzvTgRbvRKBUFAUDDeKEJcs+9JnC8cH6elHZQc/Yw76cxFK73ci3Oe2xeN+Scnx
wS0wNxPHKJY/Tnx88arW/GffTXvFRkiOziznT16INztXJSLPjkHBtNoAoLW5I704iGyRy/jW7dji
dGAdWeHaS2BeJ8q+5SMF4MKjXFZDb8t+XnLt5e4522uWD56Qsc/aC0+yeesGTh3OD5PewRewT6wR
Dc+I1gVIxAoMSVQPDgRTl6RlOhf4sAvuk5Vc4I+yCyK2DmYRVuSaj/BnqYmrbhEpYeJrh97m4V7+
S6sxYikY+Jv4BXL9afG/GueZjubJtWvb+32gLsdYJoWS/GxH4aWN/3ldz/cIK2yxqRzF/fZfu8rO
0JTf9z8HQo5wDUZzIj/ZJG9Xi081glig0E8sBiOX+dul9iz1i0v6si0Jy5CnSwIR8SjRsDvNswRP
GVuXKxgq1mqje2OtOU2+xgQrhKTDg2u7ybX0d1Y/E6eb/W3gYx06YxKLVNJJA+ibg7YpyJpxJ9Hd
P428/5tdP5BN2Zzv++HQI+yFlwWG4c6RR9sKO4mI1WMhd1Mzz+SYL40Y0SSFHJzHKSEQRAcylunK
l2vwmI9T3g8HgYdjkDYAXRkzE+kDQ4h8i5Nt32b6F0nrt9FfZ3ySZ6IQDeMQb4FaxX8S1xR64sH8
rwZGvLBbI2BDnj/N6Y8A1D9RNWWnar5thlpbKqbW+Kx6y/Xve8c5JLO0/41l7ICK3Bo7eXFjdB3p
KCyAWCRNyQstdaXkhUhtVeEmqtWNthLtnNTx30fYtiCPt1BLzj6IIW987J/T+utd6IYv+m64lsmN
HyuZHCiFYT5xx1HvrbHDxWOYDgOWM6pZIizI2TOzDpvpIGZI+rh3P0ASVeOhqWMGDKpuB/667rNK
k+3PExEaJfOkopl4XMW9IrwFzjIKW480mXAzMtHIZgOurQ3BG50kIgLGFNwAP++guO3pZKiKtuul
X0dyxLuvORl1gyWEZEmCS5MDKSIWP/OubJ5qmbEYPmeA7ucxuO0Aj9rdvLDnhWC9rrcGoX0zPKcA
PfEHLPJDFPA/NbfG5OiV2vnl5fJhiC8Oj/m0mgCFNQF0zmMfaRuGSquZCPIxDZeo6Y0/+h2j6OHR
MQhgOEE2tAngbH6UAq6EolUVUuiw3E7WqLVaROJgBQjRbjcDc3uA2vr/M4eQi6stzFZFIlvJTsRT
dgbiwOTtmhMbNvb7s0kQ29UQar4EEVNrmTCQWxKHBhsjq4dqjQwjvSQ9V7WR1Z8JRlDq993ngZeD
VDNjdrgdv40DhbBjXMK2Sd+unF5Mg8F8Isfhzg2MXseu35FkaRlWuwSOr33OzjP95RN4ZQ+mztjj
5BEY4YWYT59naL+lxbCLCJrP+9V6pp4XT9+xafxFSHKSsZzcRdjcDw9eYTWg859Z6Yl5BZO2FxyR
glnfas+1KYBb4WUmTPJKAbElqBoJVnjPVcdOw0yODDbLbAcecqjWYTVG9Lh+DcJAA1/MIYUsNKSw
i43WNxSbVQX5XmJ2eeVYs9kBeFfP1gzUCnQUS9v1mNP3u2ue95whYqIWGdWQ/rzgLQujPqfBCByF
TaaEStK5eqsUQOg4F8+DsHbONbspiO4rRmFpiHrW8USqNOTLFvwsxzpVrrDOWlqg4jb8frXGSPgK
9fdRpKYYeu7ZgnBUo/ew+h4mAqzPIAskE6pNpO9wEnt61w7vVwQTZDXxsdLCF65DVCIP5oMimK6g
TXOc5sHw4spp5TJfowd4R20V0hnhhiUjso3tmg0tnnubDGwJxESLQMBMURFSGO9L2qWRK4vRdLPq
CABQEgHLEWsHDKTjBrlgB+Ih59+TZbXc2uxJ7HfhijMKzZ+XYLkJ4mnGuwJI+i5gd+IA+GHTvCP1
FzuNKKgqFd77Verl6pkwfOLeSm6G6eoHP3MnkwTgr9xIEoZRbBGPPF23UzK+h7ZtnA2Gym/0SgJX
srZ9XYwIzkCZ3/jc9G1BIfKRxA9DrQ5s84u2wevo3lHtw7/xwkjMmEo2A1xsVATs12X+f2nRwGLC
eiTt/9r/I/SXjByKm5zfoCKqaODqC17VpHjgn5sf7o9zN64c1HjiKb6KRbzgpZ6rOI1Ei+MUTWh4
bHAbMVuLdUKPcKsy8l43VGXYlqBGsWRUvdXhd9hKWm9Nb1R88hVn382F2UMJhsI53a3IKWHIfMDJ
jUhII5lFxr1qAehoCXmh4wJFl87My4pn+0I1ZpfGshAuLJL2QOlvtil2srvYQtk3WwcVl9e5Lfco
mTD4Yhh6bL3/hs231pRKhQy9j9N+jFJZ1DrNzzoh4upqDMPexlKHHHIphIlGcWdc9eBSYtoarpOb
4wrzznnB+c5zfaiGbrJeZrlTGGittXHteL31ShWnNSCU/ubrwvkTF++ptue9JYCk2u+shbqHsUOc
l5ZMsx2PDaqWbRvE4CfNuyz7YOMDm7iwcyUk79y3hwqZktWvBS+oZXbHpWnBcslnTY+q6N924C+y
F6O3bkkXVZpAzmWE5ayf3hNSxzQspOfj1k8h5BwpJky7QqUCa6CjeE0hs7lN4kNyzrGenMudpOa6
bP9FRbH7wuShqL6RZIlbRC3z+32f0+McCiU/OOk+DMBxGjD+0ULY8V1QFuEWW08mx60z/daY7hIj
IHvuf7VEOhyaLctlSruSieqIn++ki3lAWfG1lUP4nlogmnlBfvOoft+Kh4L2rdO8+UAubNead23x
G0jH69g58X2n+a5pBPKbeTJMhAo6KUElmYicZZb0qbu31VvbrmgD8mkpPj1g9/N19+op3FS8xoqA
kL2Uw46b7cMDkcZGDeFM5ZpvBbM4tpKBTgneLYLvZjYRkt6kkibAEr6IGRkFR9xDAmwXzxW9UU5V
c7s8BjRsuFF4UrPhnDaW4PN8kxWBZTwkX8Ey8MGQ5p4k07mO1l9BZI6pTcdiJGGSGk2J1EG1P8rb
7a3WqlebCBcj91MRISdZv2fDcPsaCkJfD6V191XeS/nkMsnhYxzSZzFkgaozkyCJuozK6PQkxLTz
tNQWFTfmR9+YDkWPhBEZ1rdkIDiFu51I6dmqAik8TUQ4VtyxPl2etPjtZPm1dRL1DNXtqNfwI4tn
oO3K9ClQIuj+w37tFJSKGmt7zFC5u3QVp6AjHtqkP4NBBB/4depHamjGjTg1Q0o4iCMF81Nh47mN
XD8w7dV2lZV8S7689xZvnVZiJVikoy9mE9VDqFm5EdWav6rFyFoS2wYnaYhX0TRPOdqHvYgn8F9D
Y0DlbwQFgD51JT5njSOX/9tIBE5FZcaE2AZWqmP1wGx4lHn714JJYzHZpW6rO+8ygRn8IhHS9r1F
oy1Ud2xMKmYnQ3+/jtXPwMJI9EF1FMLDmdPzP+jouMQ6uj1Ac00/pGXNFXFXamrZH+g1ACYMItz/
aOzzJk3SWc+R+npZ3rMmx1mhVo+rjtcItv85TfaL0ZM+A2O/EhvibGZ/DAttG4DiQIquTnLbTxij
OygsCF1PNZjEnr+ycyafQKF8A71uQnjzmDSL7drBnw4wsdEbbH7K7D4CW2T30q+yNKlGuAf2uGcH
LklXHGZK2LNMAxbMZiAu/lOXIP/6Sxn511v8mYcz0ozFZGUNzjrW4zwuYHLJL1UFOanevYNZJ1eh
X+IOTj6yBKKosaKhbAXyZkpMgeBp69NLWv3+ShrHy1HvUZJYaXtPMVx7HLZaMhMfNm/HqNCfVJE7
f3Y4YJMc14D682zjKhCmns8osfs81Tr+na9B6M2ERlYAjTcOFRyPNemmU5F8B6amTFi+X1N3kbBR
q1r/bGOnhJxpwZbMgtRn9jjn8j/iYhJYw5Ji6WMMJGMlgfEQaKZWZaPrZDcD1ZNbmQIskgMTK8Oe
iabcsrrV1e1e+YhAbR/HZygGePrMuSmUWHA/+V1TuMe/G0ITVT6eOmKIAeTO+vXaxgmPVTk3t2AB
VCEyDmyFkWYKMeSim9dp2cX8qcIHVU0h8eLvCi/8hPyRHI0gfNHNov3ULYF7e9v+zzsh88x827Iw
gvnZowVL70IYNt6nS/rpj6rb3lo9JCR8OHIcDRh3WioP27YjyGftojU0ZpQeVROX2kRPs3K+JRvz
fXVHfkAqvxXpN0YgQ+9ImFTXUJiAx+H4XgK4lYOfRC0SgkSHJzo/KaGpmHPhhm2V+D+a0fxrq/i/
oq8v+5dNT+1b1OnN4WNxmD3fdgE3h/LzDXBGjdWY+EkILdGhcNXE2Fz0QXsRbOixpsT1Fla99GVo
MhSr+nQOMq8iQT66Z9f8KsYQO6oOeboyw1qQGDfWWWQbLjc48Ny8hpS8PvoURRCVDTc0EpYL+zHu
Yz604uSXp74deT09E4n1K20xC1G1wsgb205khiu/MvYxdTXYuTRplDVprvP8Q1gBopo8DdATuX+q
Mc/Ax0Uqkwm1F1Lxznl3hfMBhNhQITFhvVJe0w/zWYvm3Qb8D5+zicG8YrEnnWJLmsstpvo0mYv/
Ki7BI0MyLKQc1IQ7CLTnTkCztpuRHriprwTofRTAD9W9CqKDQDfSFtgGZf+C8ZkpjY9XVhB6auOm
1SFpwhoRlr0KBrM5zBbx9Aq1AT8YPKoMtTmTKgbJw/WjoV3tFBUBAXMHH3qvSr2zdbDHGrWOqrbH
TkGw8/dKq4137Bo/o+0TxzgCcu4UFbCzNwhuxWIxtb9m6cM+ToDrgDVXuXaCoBwkvDNidVCJQMmg
CCHInei8Il/upESL3qy1zUGhDRAFoXUsncwn6sahUQjiHaP3e4lMgDnghtcx/1pj1B2ttRUvCRgt
4lOw6NOwBhnyWH1+A+BaswjEHh+N5pMo1tSaqz/wAbFnwkQJUcBVMcdUJVmuK4bBczEkW4P6aDe5
dBxQ/nz4aVVfi/WkxQxLodiv8iTo68LBE+XNUFTPeJKMLgHJJrt3xXUGnLKAqe4WYYzwTiSxGl5v
/gy3XQk+jjd7NwBapd/uDQ8hDN3As3tLlJDdNtWaU4rrpMGHhQzX9o+KSETdttzENnWZPsw/fF3I
I5lmOS4Zvz/TELx3GetfcfPsfIJ+xZZb2xJYZS4YZNSzuVF95xQezHIIVIRTE1R6CDAmObOhb2XX
m/hd5zjmpxKOIAw85VmKtOCbKMTepGIGi29XuvlCAMFSpp33yapTG7yf5tJkg53Ir7jM+nho6zMH
+ZUBS22IgyZz1orPk7GBv2bNi8WLBMyIS3rst0m3LOdVOF75Vo97OBehIdnXt7BKHaYDnpbmJw1p
SlE0sw4DluYyiEMjvjW8xyqwJKcGpiSODWyOuq4r25hRcMZa8MIWwqDlHtJ6JoYR7RXjb8O7UFUv
DOz5h1UJCwjpF8KMRdtwH5WSRAAyaJXQL7r5f2qGjfJVCgNoqxSQeu/oFb/WCBADfDKDG7V6Na57
5AR7rI2HHTnMnC8JMr/S6CBnvpKA2yn8M0le2c2f+1lrhxoTsDUNMJJqpGzhNgRF0a4rK7Tzcbvc
WFhfqKz7FT7AOUpmZjLCIYpJXgiWvO5aRB6bVICeODSXcU/FlK3L54NVqQZ7J8L/x0S/KACYO1x5
K1Q7b8D9/W9PPi5H5Lbg2w1A4RgnXsEsFKpIm6k3yBJrvC6Y+BAZMzQw4YaPN9B9ZmQpRIPxWcKn
+JdYpA3RVSKniIQLWswHOiBx9VAVXtdKdb2ucLqPxFDk/9SbAv2lE+lgSxz5QRzvP6QRdgtHsroz
Vvbe+nRF+if2L3Of+OiCx+6rnbiak6Da5RRCSx3o9644xi8xSoUAbu3RV1iMGdJNUR1lwIxgxiKX
3DO3zNDhh4BTlsc1QGYGVU4HhIJDJ0OTSQjp3p9wUFyk3KrhpuRTmzdaK/4tfLU0zrOW2+KvupTT
CvPjdlLY7lpDGw1w4ujaTFwQFgyvU7tfmPnVFMmL4SYhQiF3qwodSyWp/hwGKZLhPbyHuhG6twvN
L03Z/SEQ0H/iZAWJXlLU2bcGMkkasioe4BfN75pav0JX0LU7Zm+BU7TMYo2K/q1brPWB7KjQ6wyq
WgFHxvqLtJc+ZaoFuFP18ioHuKqtp47TrfoDZJ61+aBQ3/lEFf1gEPDTgS9Xviqz+/VeMXeJwqos
lbtYq2SstaGbhsnaeogpSwx5af0FZoEq6vAjPUz9BwtD0RN4YhgaFpuWDfpOO9ipLq5qbcekn1cM
qo1JVNkWriT3e4UACD1rkbf0G9MN2u3Ft06hQ/BuGIRcB3PaKUtkwyIT6FjkUhpeAt3ZHXNcEXbi
LR5xkIOpRWiVK7oH4rRY47h89Y0+CXVU8vmJYMbWFLIJoagLWQjw5bk4ffEJkg7DNkE39BAzGvas
OI+DqiUlF8XC5NKJgEMRYdHJE+3lbQfzJLpcMZfpdEavKzpjxvriGeN932LHDs3vDoEHVc8SiQY3
DIWi2liTgOw1O5Rk+9vF9NQoJIpssjs10MusVKbsJ3TDou4kdmhvsORrlsnW19yudozOBX72oLdS
OckIRGHz8XT5ziD3MwE6Z69Oiuuwm94FojzPoc5Jnnj/emXhVKJqKqQkurGS2fI5hbkSesPczmLo
B6j3Mv+rI7T44yAeMvOa6WyPMYfXE+Cuvz2xl1WLa40xBmBs7+rA5xGJ4SyB2HR40zhJoEaUGvDW
OTzBaQAe/0sIRfaVc3WKY4cIWtYQTZVXpwBs+IZeEsOkw/uquaNpxFV2/ccFRCiM9VuFpZqyFmHY
YXxw68svw2HGrnDaPnDKN3F0WGL5UvqF0e7XDwL3DhffmC7XdFrrGoJW/tRxphiBaQzL4GAyNjzX
R7Kym0PX/1WnOOQpdXp4f/r8DpoVLv+mzUJrHD67oxvIFoWEUXJJG0fieV3Qxj93Bch8xO63nzRl
QDb4aoS4/j82Fhci9qzqPOjEx99uaIV8LTpndTe0YylQWDBwbg08jrqJF79WevWfRp+53kutY8oF
4PDBPIUaFsFlbaQpKS1ou/QtwZitOJ2yqH1QgwWMpBV5lg4b4pYPPdADMln6OoJZ2sn/1tUIU/CQ
0mMEAuWCMBZtw2YWVMBWczLMj+qDB5C4thIZSPxnCB8dFMJeVQTEfst16DanFpgz3Hm8+T8k/mqY
fC3sfHFBSHgmIxpI0eS6+RJ4bdk9H/rQ8+Gu3BWfgKuUnBGFZAe9dIyJsI3rD7XAi7+J15ARztSr
6bXc37r7utFpThckE/ya+ozN0smLKjvSx/BUAi+2ff2AMg+pS/S+uzn8Hf47fRDvUNrKy8z2F/+W
KRnrIz6XSwfFOWtex2FSxSxWvGBjBiqqcneizEvuMJCTQWPUlOISQKK+H+HjeMgjgCjzK+UWlt+D
59yQtPUmaYSc60rbje2uGHDKCWIgIuHjyxLqzRzmW2rsq+2IXdigLAQwJDcIByz4Ts7wy3wwxR1H
3NJYrA3By5L7Vo00HVKYd32Za9VwtbME3nGaIXe9DpBxqxMdLGs22BkYgMIERA0i995Gb/zRKtCq
KZgPpPw1u/niykcjLSwDjVhckDd/XohNEbTnIv6Wfwrjg2t6kDo/uaHWa9eL1RvgoCCW21sIo+BR
DPvtJMO+zD/AbudR2YLcsNxsPpoBTyc+dw6HDxPoGsP0ydj1ln7Dm7VI50ufh703g5p5MG+xkEX/
+vwkxkZGHFdLcrQPf+vA4aGroVh7u1kM53TN9QS671EGkBzJfPgj1F5YSE4leaagd7n+PgQ5X/bC
aj9Ffum2bKgn27o20Dxon82nHVhxTbwtC9slTKOCGZpItJyzunRlz5pgiK+VNMQoQpeHmRkwkzpg
jM51DlF/4VWkwirxNRScMjkcIJ7d5Fc4R0EulFHTB3SWEhnPF2QAECv9NZFS/NoE9O5hQRzGcrn3
V3WWbFBO+lCsGeeKnKAliaInSL4BgU+DxjhsfWC8E7N2h4zGewWWSaFeOlny3TyVJ+BF2LwHr+N5
hcrkU+64gQ9n50IqtPJD0bNIMyugUCDN7FeUP4AUyfvEsxbHvdAdqK5p9NETTP4vYzRQbbF44plc
nknwc4wFsocdqZGA+Om4UILcZB09IPg0cEF686w9h+r+6qXeyNRmt2oxGBFnbO1/9BuKNsIYJpVv
P3NggLwB+tUR5EINkQikxKeBPiKv5nTpA+kuhDR/mipSvj4fEFb0O707i/IiEN0NE9JySnlrrTa7
w5/xGfIrPx/+Nq3fOs6zxUtPCTWqqxyyecjdCvtc3SdM0u9DtCWyo038DpSxBurzPMsUa9Ae97Zg
ztuIW/wdacL7AuhUmJJcYSlcitlYTJI6SF86UjTDbcSS3alF1BUPVqydwqOAAN6E+X50oS0D8eJx
hgVoti3HkVfP4sYWUWmGm3v4xwNtKVKMT40CEYgvcxTPgmk7+KTbrNzYnoomZxPBtmOL1HWypFxo
MuxoluG2cVOLKBHW4WSR9o0OFpUolBxanZ8kB391/Bt9dJbsTOUAYeus7HUwPbcGFaQVVVHv59Qv
DrLoVUZ/O4ZzoPi9Gg4ye9kjOLnzBM29mQ55oMcTfZZLgCWeDyi7X+JA5bwQUDGSVgqqkAJitD1y
g6tu3ORVAYdk3Uebv5RyRt8SBGJfzjSUnfGGSyum0JzuqVOxh91zKfWHiC0M88EBtAdyGBL7Nho7
A5Kr8JWp9i673z8ir8EM1xOWefxdfNYnFIGqLIr9CxxPJdxcE0/QMPToz5Abg2hiJB1zpDzYbiBi
yVTjUdoGVPO19jxmsjS0hNYPFuzC2V9Ef78bngHiPsgIEvHOBIegJz1Ne3nPY8GB+7yXYR1VUWFB
coWmCBmhgmB1IArF/5/YjIQ3aPgru52v+SLPbmq0piYHIMGmdNMhPuTwXVSbNNcob+xoJeCAcRWI
5LEj7UrrHXy39BCajBznfcNqQab+D68ulJ82C68WyZqzYjS6CagAn4RNC7qQntGImFdQCPhtGOoa
JUQzIW9aXDq7iksyD3qqbSvnKe+gyu7cMRD0fNALcGb+aJLuNe8QYMGnEIDtuc27Yx8NoBf/sB92
KbJiL3edIZ1gY1ea01FmjznQ5+wz/Ycu6zrAcaWFL4UMIaJ7+lf4RFPxGT/mPSpB6+Fn3gTkD9ji
PC/Qiw7clXXnTCulmxK+YuIzPdb4mnRnMcxn6ii5PTjnKV7QQCEhqjjWWdPFwEON1TM/TtLHuigY
6l0zeJYdXFh2ghzFnNuVJdmLbGFmb7GgnYFrb3c1lROx4DxW8sWGoZgbaaQUxfkeo18ftAG4pDze
V2cChEulU1Pw+CIvgi4ZtAAZ5eb0XBcs8cRrepOUTv5ZXfSGWd8wZ/bmS0vq+4ptwgW0FHqS4C27
UlSLzLTssd40gOeG6ULtq32omaA9PVrYjrv4BOFdC85785y/wnXFae3NJzIiSDEOvkXbkQf36zxb
9Kc34DziRvj5r07ddmg1NE1dQ/k+oke0USh1WjFnle7M5El4Qe0jKcCIUt792f5TGaHeE/HEsr/c
Ces5GJtoifg03Zc6wDp697ge3zXZMsEh5sFUYWLJm2KAHE9DUGEkNUf7rQxJCrcpQ58mW1oB4gl/
Fc6/QtM7GRrQTVJEP/SvtfLgZ6mRANbKqkBZYA7h0p5INqrfE8v4pWHLQx7eYn21IAbYJGKhpWtO
7FF+eUy0dQimpmLgxCMwWwCRvfwFI4QsAJCnAGxNrRR6JB60SfLtExePmwALO6TbIIXf150oXr0X
2OidVmOo7cu4CXbSYyh9oaUl+75855Gj6k4up2icMUrfERj3i1dGXzwdT8ioRIfOGJ/JWqmccDo6
ohy45KLKQNV78HcxaH3wf43i9TWm9fBjB4KmEB4mJ4tX/7lojtivDk6eF8dAjTs3MQgDiR8QhcrV
YdCm7uNRoHf+91QW760FpYM6jTSjfEraqa/gNOw3bt4CCPtcm1DAnFVOQgirOoDEjYIjSHN3RZMe
Icz1ynhx3ncQLpltlse7Gih3jXROC2Q0YqnWWeQZzWJFsu8fKsOPb1N7ifHpw9Xf2XwEQLOz5nw6
1ZhoIIBCuCzFv0ux3dPdHq9QTQNVmX8yOhKAVVeolhxqcyRoKgUSt/ULlHFKsvkkVPuPAPbYcvar
GK+hBS5Xhi6bboMCwL2LoRLUdR2KDvyIIwd0flUrDC07tjgRC5c/YR6gJ7JlURq4zOtJEyf9/ARv
9wcJoYXj3zVL+yIcOo9Ddi057eeKZVw9s2pK5VfY9fbaMvLJB55lrmAwaslsDw6hiY3OM6+smYgW
YvvRspO0wpEu5ctd6FyqxHV6YvxQ6lTAtyOtg0j9a6EfJukOe5831LUfWXnfMkMcw1kRN445ovDG
NxXEQAWiMmGRkje7poSIGQkX2ryyoVlDSkgVCg4m+ZsHNXLXITofn6pLux8/d5fOJEMkcyGNOa42
lGfnE9akv1M+eqS2zHtXkqJTDMKRgkMpWnv8IETAOYJ4QkZwqvxRNZuObPiQ8GXgcIisRxn1qyYn
gQ3vuEP8qKDnh9Q/zibDOWN10chR+9PfACMlDoUcwctcncjhd/k67LNAXMKltCaZXfqaAmBeeRtA
PmA/QpIX3We+RfcDDNvhai7Y/cJWiiWhcyaXuyJCLNgdloV8l3D0wKx32Zlr+ecdxsewTwK6EC98
21oZX2nggnGmgNO9Zxa2iY5e75bzIZKHcZqUO/cZbzZEl7eIaYovSpafViiC7e7ANtQG5rKKU5l6
RzAJAnt8U3Rvgt9ehEywYDynTwU4mNJdHA/JGkJiVHZdXWTByzhD1JKq/N5vkeZqyuUSh+lD92c5
uqoWGlbicRrOTPaeBoDR0Rv8iuhmCjiSn6pkXykyyTpKKsCN9W6WMG2KJCfhKSuAGmjSj23PJ38M
xI1q0VW0k6Ge7eCaJZZvpBC4re9NLSEfyuumJJKVf0V0B0FnEhbj1Zqs3rytzaqOPsqNY2N9VN/2
+wnmyzjs+y4DwON/IxZe/DDfLsn2BqMxH1TAMH52JUp4jxo7qX0+l1ZYjl8cE9T/p/HommkDg4GV
JocfrugZqfail0tKxiRYn9EithhhC0C12AKDFP/glqzJHOVW5CSf7kzKjDgGXR6WOu8AeTA4gyQs
kF2cREXMBwsPX0h6zZkydk+lAwrgIH0pNXu9RMhBnIS6bAwcZbpj0deiELuH0XcPyGHtQ0uAtDaT
2/tjkM3Nnn8X8GjWrKbuii2VKjcrLPTiys7CpBikqyCzASIyHnDztL66sKcPiFaLPxOsb7W+DLcH
2CGtbsxbrq9ec9w6+cncdHUuzledxpmb7nbjirSyqiei+XPYcJ8vHuhFg0ME+fl28gFh6VO2ijst
A6LYMI5KolEAFEAlEXDcrR/g9ZamjArOC9LsSEIJ2yNPsKZNvFPrqMCYhWLuz/YswpfSBDquy/N2
7CbcgVa012qzQ8c9ATPqqwf7SSgUqCM4M2gbuG/9AjoeAF5qR+vDz6xCDQp2nEzixNFeAxJNls5n
5vec8WGOsxlGaPBV+chY0W01HwGPNNZyKz0Ng9nhh2QX6lBZdAnB/B+fUho0QbXNIQvoEtqJjvI/
GKK5lVx3U6LxeW7CPqsciMId7mQcMi0DExjcKNJZDrI7aTN/S3Dp3vXgrBqlSqsO4yH25TYR3Xqj
qLlgo3y+Ah/Ml7IK2qsF1tFFvmhHgXcft0cekz3izuhnX312EdK4LXISyjh8D86dWbjjnCqXRsnw
BZWJuNyfHfRN8Pe0snbBqqJB4GX5BMbYIdB2Sb/F3YjBXlhhTZ6BQSI9LUUp25HEuVj2VvtZa/Zo
FrvokqS8OYpRrr5WLxbLBfJ0ttmDhaI3ZpBSoVhlNxBUitzSuYGICxdD4zIuN4CPxfHHe1SeT2eH
b8tnfoWiYxkFxTyrz1QWDEhMhDcRY5sHzbSyD/NJG/J3Zqmc7Une2FARhCyk4Dvv8f0o/YB9PRoG
82HjaE7fdjr61IIVlvE3Smz7SKkm41mF3snosn4Zyz5gsrTNE+jAcHiC72kxY4b2DC3xNd0xmc/i
dJGeREsi9lZOl4b5VyYmTFkN2HjVUuC+VWtU1lHni0vFEWnPx9yQSo+EGcY00tYLimPyJC7potlQ
x/Gu42blr4viyG5PCx4URxqvJ3/7NJtkXChYid/bE9MrJ4fNKuRPDQTQN9GvOqp/jyKk9/Hgf/0g
J+1HFmo7+9vTrm+1U9AYgAYd6C9oc1+lopllKAB2rGHTLM0BMlbY1VUZ/dP1fBItp9DB3jx7cxCh
vj+8pwWdxGjnKPOkcc5EWGn0pkMxhmeoSaMY/C7DMT8Tusb2CeZnDNIejbsGQFo+8nvD7qfN99xi
wk0PM4z38Htg+iddK/+7YlWtaPUqPuoQ+h0uXVbK74PEn8dx7vGzTO0qOPtUuhS4t26+FN4wweqB
g2bLucSvG7JcRH/p+vcJcSEQry7dnKg2eVJf0rT17lIL1RoQg2vdlDrwtLWrm308U+xRKf9kuSY9
wfzXfGBMV12bG7kwFnnnSWePcpqaTww3t+v4iVtzkOOL8HzAIY53AguldZydZbu19+CDNFB1m0H9
RtEipbXAWp2DF5i/hl5Itz0OF3Sga5cuLvCXvCDOot0RPI/cmUc3X2ZYhL3M8tJav+7idFBrIf7k
iKyfMueMNJSKzfjJotUKRgIkIVHtnT7cQd6eAuWswtgATtkEHjWRJadoQdiEmj+myehhJhl3SPhp
RMBjyYQhGEAFED8cM4TvQpAK51GljbrX9WCiqv5S6Epnnr6Lf78NKXmV1nM5ZHDDh9OyJHXcW9rZ
5K7sBQo0eaLgWxW22Sr5V3w1p/BEqPHgj6+ieRWJuHOAZyP1oJTXj028JI2rpFA0oqF9RoLvyTHd
AhiRIjdNuqHLn2kOsAxMTeVfI3Sj/ryvIbRLeqfVPJIGDjHn5uQEK4y17IPzeVmKsaQ51QvYAJeO
1p/MTsnw4v8neLFYs1YSBdb0dkPqK0GD3DU3sEJCl8ZDOfsNnydkwjZzkT6hAKKr9bUrGI7fTela
kiB+XLPoVFOwSjD7y7VxUn6fLEyEZhb1sExLHOUP4FAs4UpkJVHmAvivrb8fJmbaCeFFgzKblw/v
KSeaR1pgw8NP4UTNLDNVs0ACcxT0yXiBEA1tbfNlHwW2+qykyne4a2i9T6sOhTnKe+n70hhirnvK
y/KMGPVPxVneONc1BsBqjBiMSYz0SV6D+WJwCveuz4yhR4bwz7VHREpWWGhRH6MSAu41z8xnhj0Y
4C6YcPO5EePQdALfpaOg7gWk6SNb/MiIK9mFwapZZlKscfOY7sFbXu27Nx4RFsFOPjuSpfFLrW0b
9scwVymZciBFQIuvWxBfHlET7nt4FMpJZCwl3D9kTP2Nx3MV5iuGyoQO/1v+XWHb2VcjHYRjKBVr
8hMXXD0vIRt/NSmG2OHSURcdnSWo2iFhBdIkEeP/bxj9LFBjK5ukd8Kiq41y//aX+8N6QgwmLE3a
Ltx5sDdoRTo2Ihi5txlxTsCjFCcCqW3d2cLmvILC1fg+hzF5PAoKv/eJzz6uHQOv6mt+Mfqvp3Pu
JBaBL92I+OZURRDRn59cZeJ3QWW2abgd8EMur8Aeo6G/ocUmqH96WuYxXtiI8McVx7XNo6DC3A+y
5ERkt/rAvcvobYOFWDWTyJzd/uiRM/wXyVzJ3gvyqhMBVxj7GT2yD9KmB2gI94MKPKbrX/zPoqdu
0jmXWFPpqyfFEM59n2tzqJTemaiFPdNsbU60uhnrE2kkO4LS6VyKPsvnmmwNJ0a4KPByCSPse5tI
hRt2KbmBPn5L5FAG4awbQdKkSS1DIhpeIPjXxS5ZlUtoysKcB7hWhJujala4wLEmC52J1kdHHOyf
TQquubdvHBNqDTXRd6x8894EHlXqBg6M3ByEw905AT2naAeMnPhbucWH1ZpsXxdw2VDeT3+1DnNl
v7WH3j1gQtlsSTq0gKdmA0fO4ODTlaEsDbNlFQouDRqaCT4dA2ntyD9eGbhwHjNekpXyxE5JP2Zn
vftxhLICnetE6KG3ET7/pl/mxyS4qNKxJ8SfUehDoA4kz/heefWbx02HbNQ9FjWEGhUxR4Ax9Tdb
uSg9hnSduI6aCnEhfsIfDeQ2Ssmcr4Xvt8viy/CWxlNbGua6yJFKMMw4Fr+SbDMgia4dDi3BLEva
StwpuUsel8+krrkkaikFs6JMjltAINXjLlPqtno/Rr7OocD8kwFpBQcj63OoK5pT7y+46t+E8GLN
k0C8+xMgvlODe2PXao/YbOqqLzQx0MFvj4Am/qOU6BWP3flmIs0FOQnioTxUkVYIzOUZdsTkOEHv
CoPjDQqKCwYy4wuxVvOhAn0skYsvnh2eqeYOLSTpr37gl7jvz4qoR1Ii5vfDWNbHr6GkfiQBELS/
2eVd3xvJ9jT7shGjDWWOe5V3+3okvfEAPIBFURnxVZbj6mDqH6UKzVy3iZBX7y8kDwJHDiDU+KO5
SGqvOs8ca8ne/UNhWakmdg+L3gd9sOS0j3ZZDyN0n8GsjKleQGF6HRi1ejEWJ9e6iExaPpfpaCYG
9i93b5QIixSi8XCGOAtPSpypS6sIk9bQalfVv3Refvh7hdRrUvt5zGkhqGKymipNwbNAy5Ll2goj
YOJRcq0fIzhOSd7FVgZpXDEDMna3fz5TZuIj92+sz9x/6x+sCHLnUtjivElZvRX+yEmPCNzCJ3wZ
J01WsYmSsqxUS5Qip74PLLndrc131n8VHfT/e214/MVD0KVcr2lYf7sVUdAPqry4YWrp7BOfnpeA
U7roCHZyF0Y4AkwKHqptrQKA1ScTAcyn2g3d1d2NwteuMFmOJE9ebJEQFn6wx8z8yBPux1Hxo7KS
VEqaAshujeTdKPkq9FAGzy9GEqlb28NzBZ1kfbjrmjhjzTPkUlBSdu5toYI/DA68rtLHbJ77egve
kux1IqhrXzvKKeQF/N/zjKmzcHg5IGlQC9Q0MDI6aMIbyxtv0wX3PR1FMnOCloi20cM2xzxOe7nu
iu9Qtdkd2IyLDFaDQcJNWxdL0BNRwayiaKv1XUaHtHox+Y1ahw1nmhnWKOV13HzTYYOJ0vJMHrbM
SdBGqSZVIrZvdi0YJ2rwuglE0eTS4VdGWY5haoTxFjEwbvJdpFEAi32NEvIXSHn50pXqsCftG/y2
G438qxVv4M+qZhMaCRTUAFrwu+zjIudkKJxvROeFWqbh2Xvlt2FyzyIc1X9MzQ9x5wG6AIKvnsHv
Ggpy/WO3oiTTDSNqyGgTQRwPvYiYj9+Bu1avVqQSTGdN7mJxZ+asN3cD3pJZ2T1CWUoltOS0IbHl
440P3pe7olc5vMlHY+dw2TmGN2hZ9Vc+NGDj72PQH9gGZV45Fu7en5UvGa0CIb1FCTlOlctzvuib
49SMrx8stnRPL+69/dS9dN9NHBW1SCdRoXzMDFb15w5iy+HEkdhFPYoWiRbhozXe85fo2Rn81Fl1
QJbnY38M853tP0b1EPyqfTg/XrfritE+hzXWsip9RjEpiyTyRoTg2nyiQDqwklCAf8QczQ4UHelf
BV5dAy0qSkdnA09Z3cGZaKsSO6uL1ajrNdz3QxKag5jvQRLqysTIvWSBMsmxsB8qouG1VbHy5EiV
NrJEQ4WT3hh8t+YQE2oLnRnowVka9iA9tiXmNHHnosvrN1XnNLn6s70diJ3X+CF29+0UTou8lEMI
bt9+KchQj4nn+8o1gktQprYMF0U1TYXPHevq/lQw09JAtqsU2uch0Pvi/+9RnwrbL0MwL/ocS7T8
xzRhd9sdm+C8964hCOSDekawBO3nSLBTblB1E7Zbm01OOg92pNCQFUiUDKijzi2M5Uji6yrIhRsm
i5iHRJ9QiPsqbPdTHpEipqE6eUdbh7rlyZS0geLmnj2pQCZHClElwKUvWc3FMTpC1D9AiySMNwvA
LmZCXny2RBSCLEP1hC6oL6G5auKja/ta3wzkLeZz7F/GwusPnuWcFvRuGTqPpqk+lNtJgbK24bxf
VfAJxDU2Vl7Cw14Hy2Crtw/7DaO9y3n4buHy1lp0W52swUczad1BjDXDDUMdzkbRugUuacU/f8vP
IWSWk3yMUyO+H+RH15n1VukP7OqBUE24NJ6HlsQ/P9bNh8yqLGjC5+yVHmxf6rc+BDa1L2CG6HMq
NKFRHOUKYmev3hAUYoOXUpSRbKnHPwPw2qQ10S3yqKqH5qhWjWYvFb1h+pabrkG7/sqB78shiTmB
Jn4hwtILSmFokA7tlZzp2R6UEZcVmjFuaYMTrg2eOgCcvuqCK9JCz6MxOQ2kQiPOEZZyW7H5pAsy
hjdShRgPiq8Tc0BnXevqD2LSp5xAbfyefMf1D6lLfIIovVTaQttVQ82nrRK2YkncHmBY03q+bT+6
1oSMLKktn6QRluSj4aSz717So48AroyhLS2TmRTDErbBLTIKn1YPCNs+Jpt3TWo58krBIq9FcgKd
uJjhUWJyxkHCbHLrd90If8wtolhSu7VC6UDrx2Vu4gWNFeYK4jVmGh+Iu9Yf7A+5Dzkn0em5pU6B
xSmm2VFOQH/AMqztjqf2Q+6I2RXL+RutAi6dAi8FImTc7Wi5a4F9ArTnJ0/xxwBV283LjA4ZQ/Wn
tTCsD3Cqgsd9Rrei3KdtZiiCVpF59wt79CtQqErUVJJnzrxFc+tizaj6b+ZBOe8L5I7Tx7Yt3Xti
gqrLvW9CEMnhcCHOoBvjVF2UJ8AOYElJM+UCyEPzD2RgGoX8ckkVh+XtNqktFPeTqMDn5PEmY5e0
posY8lKBo3LruwNzTb8WeEGVNFVvIFNZ9iu65FvQHSNrg+y4uA4mjXmddAB+1vZKfFMX2wyRY5J/
fn+iWiqQndx7k8ZGz/de2p1u2lPbLR0UrvHZKGYCm+ben28VjuG2qtH3f1bReIr4E4g1RjNqODfW
cvdoR+/rkJtywgshflPzIXIxHlejtynoI4Qm1x4LemezcqXVnh5g69vhFg8QNtRFwwC2n2yLYgIm
09fceBzZGN3tbKiz2h214XebOEnJ1aQUup6V5IvUucvVe+3OdcSjgVGjoB19rlS3oE9gvLJY1ytk
LaUykeNXc1sg+HC4xXREGHciPDlSfMdKJXnlDvTMn9jYizrd7dvhJP7pSmS6bHdN3cAOInXXEiox
dIdpXvA9IPFMqz+HaE7Z6ER4nnJaaeyyljPo3ENEkjJOHuGAwEqsBWVA91wPCrfZDprjutTGjo2s
pJM/RIEWA0XK7jmg7fFbtq/O5MC0LXthtHKzLyxzIvAfnCesmjWQz94tSy/wBBamhNfIyTBkddk4
U1AD2/zs9jHdoR8m5YKjuyPOHE+PqcHaqABZeqEBgbl6vketIfbaxelTJOtEiSw/Z3hvAwKNZtI0
nYn/W/2z47f6bp7Th476iihU7aUCebowPC5QLJHPx42nQWryxhTYEmLhje17jwBhzvCKzrrJFAxf
XdhNFniImyLGMrnd8CKE2E/Gj2JzFoQ3TPJlf52iaGvRuHe9hdmPO6eGHZANgzQRHrVPwdTj0kKE
XNmatecO/tR1qqv3A4s9V3N38fYXnh3Ao0Uby8ro4cyuILBbDDczg6tPG//MmHLaWHTe1CqDcTmX
3BRywm0QKynHnbFKVU4nqXFIC9fmBenvpasuJFJQvo/b/nq/YgGUO7kv/pvHw2taxO8iiulbuTI2
hy05BS0kVCKVFxS1/oqQQH+fWmHdhy40meJE7mgjUIKo/stQ9JHmPeTIEN6tHqphq5AV/26X+SNN
fBCtjLOxFG+wubNFCcGJGejZ26c5rFZjDqLweXUTrGmnznFQxmJPE0TiEigznf1ue+z5LX3Mvp2h
T/ke37CftjSdFTIUMej9odBhOVe6Ptti0uQEzj1XvZThyZnsDhvBQPPb/oip6WhZYR3Q6BSs9O+h
Hr1xw7R7r6GEjWMgNgKzKPh+A8TtMu+WUptk8pR2Q9ceRAy1q45odMC1a3j6gSzMadQjnormd8fB
2Z499sYA5Uu1H40r8T5g9fR1bS8iuQQnkJ7+oypIThmEu+kPYth2wI/DsuIMZkvHNRh8v07OATy1
//dEKLa80p8crtIO68g0YknsjoiNN9Rf7tJXTUsm7Fl6kLlJc1TElYma5RxwXxg4GjGoqv3MIrdp
IinUN1ZmdtMZjt5dS+SYuh9EN5xVre/jT5GaTRs4R8X4/HtB8Z+AK54bluYKMYOwwpNkVxAXboYH
6ynPrK2C6x0yiVTJpNhzBowkfuDv9Nq4XXb6LGgam2JBsMQY+Ee3plxrgtLqV688gYOjGPt30LuY
mk52CsJ9wskzGpqbcedt4P2yKmcMKtIdw7/CEQyFcmks9j3EezlxSYrVD1nqH3K7la3JrPyovl8z
uHx58vDN7FSPa9ERvypX/UWZSOhc8KjdL+C6aCDKwHC2n6amTNAEBlEPIhYD059anFAxz71BBTZ1
mk5Of7cVQKQ5Dv8a8orHVu79I69jBLdt2cfv5HwbAJMxTbLg4haQXZXT7uIALc3cFAZoKNlThvfM
uptwV8CIQh2VRiI2r/DtIrGX3NswOnKJt9KRDL81OMKCv/aTqIDqQ1ZZkurf8wzBqag+ZAeOs+VG
FRPvD5ijTMSdaBuGCQpvC3tA350B2ZljJTxsbb0kJYiLxArEVlIc3EvVlzwntvqGns46hL3CG+Be
Igq2m4pi8/bVwtTHmXpSJGFdlt/8aQKZW/R0HzhlicHCNHtKCLJLzn6/T9SV1BBQelLt2fBk1ylZ
+KrQIRLwMHDREhtKUeCASVZwmtoknF9DNffpR5SQzuc3sjlpDl3VWOXDZom0j/xGiTs4gy9s2RUY
+FT64RoFbMdX7nvP3wVrRI9ndng9TfyqBnIDmy/E7RVzb0U7k8jwJeEsANaBstZGBKMzMnLwnEWD
tI04Ck7VQ47LHR2mNDU6LJ/QR4IKF/ukPzPlBhAvbwvkKOfOGZqrRQa5MSPnB3kDN9KVuP3/0Ajq
vRMTxvDB4lHwO6IzqXrDIrXi+6YDRWJMKFWqJLVLZZW38N8oPj+UHxyHkpk0dc6GCOHozVL0Fja/
QzUDKscAAfjTuGpyZtx0kyQeybFZhXCGgSE7bxLoW1+tq7GOCY3nhdohyPAccZI/K2WpBj8aqQKH
WY+Ldk7Zk1xS2Fy4HSX1X2NqpqivqHT2FQxic6ViQH1SYzXz+/Y40+k4vJfPu8tlWnc3S6ra+Dy6
twRcFfWjhXUid3vNBm6bTjG5jwUQGrIctxDtXC8XL8XAJY9scpLGTFBPihuULN/OQqbQGx9VIb2V
O/yFMUhZDb7c5V08YsJh0lhD8VXDqYoSKQ2929+AFhf7AbQa9u/WQuMMRX9HRtrN+2LuFG+bchLX
pxwnz2xInWoiZJQZ12ushe5m3bQEJuY9usxu5xXulwWPEGAAmFnUNghpOvIqH298QW1zWiItv5KB
i3CsTY14A+V08bm1ugfb0t4//vGc0jJvcY2O89zcCHUE8qAkrNgP+X9LfAM/EtpmfEbmShQwq35j
Q6TG4idYzIsbFLhzg+Ldlk4qgKN16QXkw2JcwbfCS7aPGlLK4LNQemY2Dp1P/OlKot7cfFfS/MyO
4v51MDUblHHjDqLpfnIH2yPW/sqHwV2bExiUUX+HLLIpF+6YmIZIX3kat/6pGVvgddGGIvY0L75f
vdFbFX1Ryr0j6MGdeCDVbFY2s7WlYDFTavMh5/5zim1D5nCL4IcVTyD+Av5Ahf+5/NdXiV/t1COv
02s07GV82tjDhfU21AXedRB0SiJJIzlCSO0fQ6N+qL9tYS9aGm0L4gCljvRkYq4hnujfTMZFvwKL
6y9ijXHHBTwPIKHQISd/tzZoHIFF4mDvGxSCX5pD3sJQVlZFNQvNXc1/Q835+VOVcMIVJ5s2gjgh
5BcsQXb25g0tgS9tCEkI641GBYAA3g+Dmh8U9AJBwWNLzIIvm3fRjaH51t4ve+FSknYPB4ODvd/s
jijRMDjULh+p1EXee4giqDgQkL1vxRNBpThF6OZkSzy3tZCVetyGcC6OW3bIQLPUxj9sMzWUNjeF
wFiSgelUsD7T0H1ampOxlRuYIGy/Xyb9GZhDYcm/cZIQJgKwLgATphqt5SqQQxARjvrnHg0u045N
go/EGsk7mzORBtMDTgUIGa9rdxVBx9m6QtGqe54YIp2+d/CqtRx+oJng3PTCgedRE+ekhXzOxw9S
rzqo89Vy+2cbB/AC9IoLBXNZfoi6+FyIsJItaPA5JozDUQitdPjHa+2oRZAtn292UYEpQmmigKcs
97ecjTGZv7/dpwWrohtuxrm1ROeCxQNQol1MUtlHAQoqZKV3TTz2stc9kqO9zwH2xzkwOVSh8z01
mfCM9W87zlj/JQwkd86MdIcUWHzakNB4PWk8k2aeLbnYIugjfR0mWJHlQQduej6KZk9N5hl3IvKC
RMsKmdMkP5oAXud7ePQr5mMjIWZq5lcv44JrOX0OtNqhmWLcXK9oCBVBGdMEmHZGlP3oFqVtvBqn
b7iSBSXfuWKpdnFhHcc7r/9aW0pNcjBDz9Vu+Z7dffzVrA6eYfrYWhm0hEkyR3GAtDtYBxsEYZ0E
Gnkjpl/dlEbgUZPtLtCX4mRixF1sdqqb+Ulc4vXhDLmDvqNSf+6bFW4rNyJwlh0mShuh1xGAycy+
OBnlIC3gebj1zSa83oHBe06YF6pcjzvZv1PtuyBwwgPv9kZtCa1IvUQ+Gj1CWRkPXxeKny/zZacm
76iMS40raAI/c9QMS9fuq5sAyVbljuHvvCcGzBAjpLCYae72+kn9WhgKIUI6JzZ98JVhGbYRbX1i
e06qw5GVU4cWVbftxF1zPAXK5WkTwDKf1sIdassCgQ76cmobyOBOYsCwa1j3baecM7vUg8tJr77n
3SM7oNJzhIlaaOykVwKr0g25YxJUjnY8Y7F1hsacSJLP06dgA6CAtCIk2sc6uXdobdT8w2RoMTvG
YWO7fvByjmaWp5IyHxfUbNk/8UfWPks4iILyGl0RarKOJ2izm7BnFFfY82cX1YlZLV4U2HVb4Hv5
jw5I7H/qiiQZmFs9jtCtWOI9NIjc1hKDNKPgsN7zUNcH7+kVaFRV9vZGSNxCEAn6l+LnfS+8tT4F
Es/J/TZ8E/LRmB8ERRGc05+gElGKOyEFHLBHiAFGvvQF9BaZJC4Bue0hG5dPv0PR43kfCtXLVDxM
b4cIjGItKLWlYwKVFe44ygmzi/nzCyYng7dA4sg4djXQNb3RK0e7cdY77QSF80c27c2svzCMb2Pj
FNJQICYvgs4BMt/6GEvkhBZEGTllRetZq13PRxgDq96YSO4XePyDQNEWf/zOHd4xQy9lMfN82VJp
VUyyEp2K83SgriNbXQw4DR6DBo8W5oW+WvEHCqJESQy7/CQ3tfOYvPDmtAFiv3pd7FLcL/ycD/dL
tfsX81thQNy2sjm7difWETgcv3VwWu5Wc/FmDQW9e3WpNQET8q5Zmc+IBnLm5XAM1v81MK+awgYK
ywjSS5zl8Wf6FQT7DU490vkPXG4AckTanQRaBbha2dK7igQ5GXRcywqnQuSUP+ASzOHZ8lCqRZ3c
kuy7xX/T+bz04IYilrQpMOnGp2mBlBNrxzpWTFpzcVriplYmBPSVDo/YQBuWLB0IfDPPV1rSexk6
/z6zoXYFpLC0uXgNvFbz9w0/nsRtk1hF5zjkHyJxlK7xcrZBUWRrbvmT/l9hyjkhVXzMs2WMCNPa
7P6yRMGKQgbjVUFpt8Nag0Xpt04PapjlRM9jKNkFGqhnNoVeuQE588fAhqCicpoLp5DIEj12zbzs
MykUx9JA9YSKJgq0jmMgrhpr8T0xVmk9CYAdAYEuORx6a9sf2OrT6hUUFtuQTaPxlzMuF/eKLuKk
axYJ5ommqdP2t9Gr6jpuYpnsmUXP8PdDZDUzZzuVfEj+8AuCYSyOn0ONuTsgcH3acsIrx0nEOslC
eh9Cv7qfsV2Ypy9s8imUzWlYlP+RlYI1kkjSwWIygdm5zjbXIrR9w0B6ls+VV/m/YgCl1+QMCbGG
DuQbdj1B7tL1yiaHXRbEdn4bCsJRs836mOUHn4MYpjr4QjO7gZlsiKvFlr/RQ/ggyzSZFsF6UZS9
sQyH2uLzKLIZgKK1cVLMPgfxJ6KAVkZZ3TutkhE2vqNdRoRLYfIFy8jT9wL4c77bvECw8MRDtF8q
OaKf2d7mMjlGFCJDeZMI6HVyahicL72bnVyXdjbvR9qpzafMT54gOIj1FDNCXuhoX/UDwsrEPq+c
Wi5S2M4x+WMB2XkZS6uPIBL23OxWTaEgm7JMUu5rOEMLaGH7bmzFyMGcPm/mF7o9ppucasNlf3ib
p2aqCPjlkFt+lJEE7u1cW6kh1otZdx9EPIQ95oItd3dAgJ/kSPx/EaTcucADqdlU5I2rPbmTDLU6
ik/0KEeftgPZIxU5jWzN4E1zDOshmM6NfnfCQdPPEGVcjLoFMYR4goR7DB15MbG+Ap9pl/2j/bxs
tEUoKVW2DDAYHTb7bCrnlxTLurLof0WTcHRH3bRKdr2R8+RZ05/fHtzJbefDfxehhTyMj9mEtXMm
fbR/dkUGKvrhf2KWRCxWdmvs7H/QNa6rkCe9+jCmMuLVV5luYpTo3e6JU/eVkxZKRHGKW234jR76
eTBP99En+N3CgUXtMet/hr0dHj5j9Bw3vTm+uF1aWoBAzwdDG/B0npspfuvfGBMv2Hql6LgWgSYg
ukiW/t4AEPyHmtnigFgWuajKFZQdEjRq+psoQEl/gXTj7hVvoVzMNSwHkbzAwIp0YAADREtnyCiQ
uQ4D6JXINXtl9UCYUPn7+hQb/Qa+565XLpyBwP/crWgpklKrzKl68XTJ1fzIv631JX0HWmgGFINi
oF66oMNl5CQBV064dF5Hj+pYiMGiwI1OrtZNOmfpi1HWJTgNRzhwCEIKA96dqFaaXkNkGCNzWzAR
W9eMls2B8Ug1P9j912d2ZyvDXtOJkMG9HYVvj1BacAh3yj7uYRxa2hMbsZOq/tlJDKWdzFRGMMXz
CGUn0BzxqJGlf8yc72YbhataqGhRQU4cdMZVUihTdmLqUzqKm5XcNk3g7DvyxvFiDS9TACAbb36n
NTk6MlUux87b7gRgu1PTKdWyEGO6HaLETP0cYjo95iHhU9wCzFQEn0x3Rd7Ij4IKfW8mMr/p6m9B
m47BKs0lSfMe+lRIq6EVHqhkDUq9muGKR9tEuQtVGoxytIcbLnhFN5+S+CkSQzZSxJ0DzIi+krYS
G3S1PQGoCPehAQ7BN1WlHlWM02BILfNIl58+Gd63viKigheEHiZ3xDTJpJymhibCSB/lS1BkB4HY
/039KT+DJWttzjBQebBOJ2777ohCjdFo9hiIu+qssK375CtDqDfuV36rnMTurBTBEG3eU1JjAEVK
jehXFb7DMvNNPMjNM0ZCaZgqK2tVrgim9doGv9av7FxvrL8HbQRm/h3hszKtwNkxwo6/pdeO98C0
vT3bRkKNkAdb1p+rx19X7UdD9boUbNSkiNAaTOOOxTNqcxzWLwEhYqgde3JCUmvWx614zTpH3Ifs
p8JySpggkyo9oFIo2kWtkPxyWtFa1NbHB8bQuEAR9LbKzPK3dWpI0twhTjFRFSiTOp8p9JjHGXyA
nlhsRK2mfGUdQPlqS3wOq7GA4HMLwMO+PdIO+VDsM26Jqll0WmgJObfI5yVQivWpCHf7EHt4Je3N
oL9l+F/y+DoIusl3TMdPsVAT4ZbZ4hA+LD1RwvaY3xcz7x/Y7sKD1c9UzdcnD4OdKcHN1xoeFX45
8BCj+yzB0Fpg5fRw3n7btLwvEZ380AZwB5mDuUvx9nTx/7Z990p0LbWytDR8EnaoVLh/lAULvXva
gumJbiNF7WgVwVNUC4McbFRmxFqGyt1he9zCSpUQ+Omb1KM0UAjOZX9GmO9PTGrpcwsecEd0PJza
iR2Y5qVGdSL5jmSXCf6ZoWd3KgwWI3NXqEBn8V7BdW92S84B0K/ksk1e0svQWApmL1v2TTEpy2rB
ZkkYUxMj3JCq9/AF0uLCID8RC7MunLjBkb5TyIk9xGE3bEMFFoNPloTDRSZmqDNW1VYV3D55wIPO
IKHUV/ZMa+d5PM82S+3nwkRvR3s2cH4541KxaUUUN1cpLwB6jof4w2GGaX3klKCMO7OXadCSW+5i
wYDmLGGKoCcVjgS/YAhjeJ/6Veg7LUWEDiJV+96yQdbXpmcfQm86aqWo1ehNn/hp7/pJctcJ85IU
WbLrH1araL8XiRgfomWuXcu2tHJCD6mx2hkdXAzWpqR2XPBuJJlW/He2UdJx3v8wfgLB4Vuayaxq
iqPNabJboKOOEpTS76hlopLQcCEfIlS5ZqW/gxrCKaFanRquMRBd0LTPd12VP7UCOaNbDlx9rFJT
0p5bGb31XiDrhIME7zu071y/3IdrDugqtBrCo/bg54z8jSrOQxUs83CIQsjNRJ6VCrRUYmC2/6xf
bMXwnUKnpa72egotrl03Vd0dJRd1smcP1ql5vEeG+k879lH6NkQ3ZqGNFNPyXOwUMS5dAfJl4IAe
JV0smY6kAp60etiaxJOmeYJjPzMmxdq7V2A8Ux3SY9SUJvvuxGmfX1hH9pzPdYB4F0BQXRA3kjAG
I8JaJ5WFuRdHdpNS8XU1AX3annEqnv7y73Cxo9bTYOWaZpSkQQfRYrhH9Y1cuPzxCv8+jtp6m8wq
UwwABE/x0gC3ieSh9ae2yuWGu/Zefyb0ScuaO8BLRyJMpN5v6y0k3NBUC+bvCEifcE4oIXf1o+MO
UYOwXOgjAdmNodnDBqsVwBIYDt1RLpf1iw7s+dUIygdxvL/bBYBHaGlBICs28MelvQNx+EFgIbUx
DVmocvZnMOf5nm4LVOQkz2/zIs94dBYnuZypTp9gopBdBKXO/77XQQ6S1aq+CpjtgpyD+P0VPS5/
H5OoKdC8r2rEdfoKt7HdkL0lviWCJce1j2EBYBMuhnAGY3gLg/rA33EMEab8piZ5vD6COkvbratT
DIgwhvLWVzNEVC2gm8/jX+U58d6I54xyDYwfZxQmieY3r83wRjyFNVuHHDLZuJpb7huDw2COvoVU
ADbxfNmiheSBj7r18nrdcZ38OQdLpeHZKCZrlGeUb27PufEoZiUw5jw2VVRG284ogA/mm+afLkoj
P7NCvpvZafnm7ffPtngVITP9m6+uD85AYoxZmopaknlpFBJ5KhpaF5r2vdULjimVE9XvwHP5hWLc
AdBMjCwSwubsfOsulA0SncNw5uauMmnZAuD+T/he9kmL8ffsAMLzGVvb1hNAaMRiXhJNsL/zVxA1
9b2/CGTJ7M2ivQAEi77/4moug5mS8laIHkLL83loz7Lim+nPZBdn0ZA06/3rIdj3ou46Z3BQeaWD
stmONBzJq9V9a/WHxJwEJzVoWzi/MyQ8+Wknwml0zypRB+gYTI476sdyY3aLflTjaXMUEKq5EbTs
kbPIJNKmiPz//dPxVv/HtPDMKEze2YEKpjImZG1MswRkGXcLMUYKJ91Vnd0hBFyMb5WwMRoL2Mgv
bj06BJaH1nONLgDYg9sqYQ69DvgppePa2M0bmbZrn38k+MJV60dvj059kKT8kabqIiCt4wg1VrXI
gq91s7+dwEA62+9kwrl37ZFAJPn2WKIps+w7cCqMPrzQLMTSIUt1EgPwZmDGKYYdZk7y7Qnc6s3s
FiBUNymE8LajyaU5VZq8KHjNNvJajalSFv88jVj3P6NiRKjpMzRjNoJn+tvkoZAbca+L7UbrgwHK
ybD9vHEonxlky/vkekGIu1KPlQCzlB+h7lYBTtAZbryQwKYyErhR7j2US6vBjxzGfsFjeheGsdVH
Es89ZHAk9JITU99/HcXmA5mZv6mlMeAD0rXrja/Qc9QEIFpTdEzam2ZSlKB4SCdkAI0g3kUxcU+R
NP2wGvgLMqtMb0HMSptbCDbsIgtstYc/JjoaqETm/DtQaILJ+r5946yvmBzJLWxnc7O07Sn5+61a
v1Jr53m9EZDZGu2XLSSm5Tr6A0YbaSZsYsHYHDZp10B4z6acl+WKhdz+OWctcdauqm1zZF5URf86
/Q/BKdC5u+1Nr6i9sOdXqYAm5mF+1rtWtWS6tHMRS6sDEkDQEVtdIrnzHsZrSpfJVBX4j8l5G0Mh
CNfwUasWUj93jX+eO5HeeEfEeZbvIG0h/z8YPMVKBwNNtMI0ZzhZW9IOMB2ftjXwou/Fui2lLufa
x4k5sw6BnGJvQS8//QYrfPswZdUrCPGDAhnl8ynEun6oWWLAYLqoDAeSw4yKL4vS5z8zhU8wGX5s
BXHbwp0RmqYoew4N7ZIKrfOfKNin8/imwHsVlsTSxOsaMgoohlgtwYlstWoD/TklaVQPxa149F4X
BlYF3D8AVcw6zoASKRhqTHkVzCwyOMq0glVWUrkaFH/haJVhAdebnrICzGeHYccxpy294y7H+LZU
LcU7GDihfvQghJ9iOoxN1JIwDEC6JTBplZfNu/aAPpnScYrBYMSFOICKVvpPt6IioDt5EFzsJ+Kz
f+8Ap0YQN/IFNiX7J8Dd0h6xVOynM3HtjQVPt/7SPungvvSYYT5EMwy7c49EuEu0KerIFiXJBNaM
OwpmecYBPoe8azyvQxnzGrvcCcv2U2dInj26z1FMI6uoMTDZNgYQs/BCS4BlDzSI/tvigGcclIAQ
FSYTqvMyb8Q239foSppATK0My4JD+fS31JW5T86lUrZ2yUIe+IzG0ke5VXLrLNYkjOH4Krk+fPGb
9sNlsej84JVqk8u1HEO5FyOeUPgLxZpZdZQ2UD3DiFOfa3LxUywNSnDnZ8pBiM+NmnzD5YF3/7E0
VW5sqMO74f0yi9wZLWej0U/jbMdv1MytySxuAzPeJ9I9IKRFQZgWafPoKaUyJvmx7aLbYySUaAHg
Xs2rO1pX/SjYHK2yZVd/ZwheacMJtwgzVHJlTYtclNyS62pLrU+8wEsv7Bdhpyo8ZuFLDQ5zrDqZ
WWrdaPYD8Va0501Ngr+mdU6Oe06+6BsOzgP8QMWdyLbL46dRk/OqiKsyNSCZTFVkCUV74y3F7On3
PJlNjgeITYYVhk3yP6xNDy8ErUL+dIm1IJbebkV+NIg3gVyDJOX7Dd5JVKYfPMzucdLcZZLNqjXo
IJ4+0u/OnNePxfCdi0Wl/evwJMCAN55MdWPbpkwTzrSqoiwdogmTsA0+Ctr2zFMoAVDHM8nl0r9L
IRpZ5/PCs1iY3oCODmxnyH0uKt+2HmlB3McqfEPoa0uZzmdFZDMn/XWnMbttrUZ0Dbg6UeYqC2lQ
xZ3qw4Qg2mgfj1VjjUQbUEdwBfevMy4h+N+U50eQjw0EYqWHIz2ASOhFadCaDPlD/ubJe9a+2P/E
0iRLxbeQfoLP98k5IKz/tTsSHZzBxNNUa0w4wlurbi6OY0/TNQVRudw9ZdsAdHWWoEaqbdjrgUUf
7Xo5LXz2SgoMGIbubWmQ8YoWDZKTSmhR3pRHybSc8e9J18yae3BC4An4EEvjVep8n9SjMgb7xEr1
cQhe5G4iOm1vaDyvFU6RrBc7gq3TdAsLub/gmMaKQgxdMRb8NbcjbE19G9PEk0k69lwrE/L5cBGn
UNXCXh7jJJv3e+pLWbfU08eQcdLwdDHLDr+cdqzf0onmdlOJNhQDBZKGzThC8mQmju+gLGGoHWvj
XdYBkulkznfSRo+HakLFfjc0H4aPXIZnOOnUh68LsLXnQ2EwAfX0/qPkTq+efw6G1WjFlYNXxYUG
zI+RPzT8folgwxwDpEsjroJnZR6oRESBFJqThGTmmm/N3kWknGCHvHEQlcK4rYUG39Za9coZSIXy
Y6GIx9Q1bUvOuDamRg82CFUQb9hfKKPrkMKzKUvJ7u26sioR4LLxt2jFdP0HD4C6GpLIwR6LPdpH
ZUc/QhnNidK5FhKUFXDfTViN9Zl6RTINBjDpkr0k6UOmGWbllLKpcyfUCpZj4eCbd/yHIc+Bv5px
ynKjJZ0bxfGyG008jveX8gNX5DApyEEO5p74bjnHw/E4bIdYItzWyYldihOQOnotUZzlv5rg+y6W
OKPQwtHCTpbDlrLIhvC5RwKW16otzZiCulQZu2eVawTFvQFstTN3p+6vMolwQPOfRWNtDMFdxHkZ
8J1N0njTjWSLKQtjt8wswCHGbc6xJh4BaKNYa3sr0usXFQLxvlGa+EYjUddxurLjouw9vyraaDym
GYUaUjTVLzxnI9y4+Q3HQui87S0oMpTi/D/6RWKVEIKoo0cDzU7cnCwbS24vMaxn2Eis8ThoaKg/
ALj23NATqvIcIpwCMZykE7K0cwUon5OK19d0acn0uVWdJ5SbO+7iCfoASiOYuUPtiHFZIQCisMXF
OkqBfDnGOZnIGkYA+nl5l9PpT/+afw0rDikT4aWJ2pKwYTgHBGD5fJLSRlz9ISTGqVI95ebMkDS/
UkTUKZt+iR5XfDsc7xMzGVZ2aNlQswM6itqlE7yogBNklSGuR0ydDZfpAXW+Uk/XaX6HnCU/hZpZ
NDq0tvjR9rO8zSE8Y7J1/+rSzBbXkPmpIKsaGmOb4rJTb586A0YhQqOKuYp2nl+Aht6JdwFoj+sl
OZ+M9j2wwGywE+Nk1V09GZcDOc4cfBi9pHBJrjAXWTpfnhCd+vPzuWUOm1qSvqYmdQDWH0aT0Sb5
+5KTs/3K10BeSShdRQj92Wz451ntHodZv7Te1usZBL75mA215Q4c+cPuUwFhv0fBdlm2NviUPQX+
AiwYHtNOku9CtO9IW0qXguGRPjDhvdu1rDBqm/Zf3wBLWRnwTv4hKf1wZ96gegvxds9zOLwsjbtC
zEgrbxVKQwhvTf/LTrZSR0PSZlNhuMPsM0Qdh3wKkQDcT1uDEdAOIMPrXDT17J9JZ1upCB5WvbfQ
E+qUYDSydJLZJVurNFzrytYzuvSdRmltgaEdfliIE1udCUO+NL9JArLl5V232jtg2DXjY3ZxMNg5
M8x+1/zKxgHhVikZjiZx7Kn+haT4Ov/eAij5JBNfiSv4rX0678rz48Oy52ih+7CK92y3lT9mcPVy
HNwhmWV3lG9NqRlA0Fkag177S6cv4B3j4wKlgjtzea6Ft8fBTif0qIPq1nLegmAAIipDnZ6PNacw
kNKtTwvJmB4JmquN4A57LlkbfvZV9uO/0C2206Zh/4RiennSmITxL20rSLGK+Ajt92t3oe7Zdlab
kckgg6/4t9MqFEoCkI3g3hepG4ocVozX2h3q5ggne87TgdvogF+1D50kenbzxariuHPjUW/Q3wE6
vk5HDf7uGdrajf+xxCFDFz2I4X9zrezJhqEIe2FUV8YX+/Ky/aUDTeVWeGV79chTXPU81ClyLza0
NGYjb342qtkY+I62sevQkBQJtaZNiM3JZa01OY+mVghaBARbyQPpzHVf5s/cIkwJjpoUqmh5ZIMo
QnF0oWuhUShdam2vf1Ati0UdcqEYEHU6I2JOROYd1GXPmKCr9CHkh2LBbX8nzyP9j01f1VRwbXiT
DTCR0I6X2iILztcQdVO4WaZD3l1n4S+yX9eiPlP8pECpgZCgslIFyGOlldGy858B0uQ4CLgGHH2j
sfMSiEbseul85Mpuc8fVIbiVEhQEMjnUiK9Y3JGrZBHx6Lay+98lfCi0vpScxdV0coTz3aENU2WS
2lp3q1vzSYjkN4zblqTEU6xHbPiRHZU9BusVykIe/kFRHhVIg/bvu+nJIWu+lun66HuUHXP7xgme
jHSGRr2z5tAWI71UUyeFG1MadvALOQ9K0vNQb+4zHdGtt+M8HuVTBJ02w6DVZsMjW4KNe8I5OPXn
050DcI7AJwOzeg9rSopkJCDwVCvW0l4tetdt7agOL55ZZETznhv4D4lG4Ie7SQTSUkBo+SggO3Pp
0Pur/QlxI1w+UR8/Czc1ywH365Aq86/G8os/NCWLAAhNS4lUJuLjsiuCxLBJj9iCvs/94MJPEN6/
QI87frpevhApH4IveXiKKVbn12SiJcoYjNb6Ulig36ZaNnAVQLnGr8TmiAJeT2IjcnH09oZzODaf
18gkFk1Avg3Y3yqAyRqaljTrc9vpi46PrxdIV55FZ34QUl3A1LW+2zE0LJSXp22BcHwkIn0PcsB8
JM2DW34Fmr2ckLhHhV/kJM4xAimGLbEtyFVcwgjDfGvVpxCAwqGx6mKsxM0F8QCb3tn9m7HD4hmw
pc6ACDkVL33Am/U+c3o4LpZ/Zi64JJ5+/gN9shVNliaB0PQmh0RcswjbaSLjFfMR+7+hqecN6E2R
85bGAhLF4pmhkcy3jVMWs9QWXzxSddd4ajayg3jxjouICIWKCGFD/ttJfXr16Y9o4mwLVSc+4fHb
st6J/oDTI/YMpKFweLR33WHvjc10WiA2aAQC1aunhF6uyqGpoP+fgQfBoEs6UjV2tSEtjMAfiaXo
T3T0rnTA8M4/vnZ3/iIazE1/ZjuKNZ2qRAKuDUFK3Rd77sxpfk3X01KK87ZuhLhyR9sBQv5e+C4i
iGGUn/8C94+o1vp4TdnyZ/HMVBy8z2R1/o9SG5yzctwFqPubyBtKSlrNXimJTwJKPDxkDPgCjt+2
3NXU4kl62ULUuHFRcjIntkITlhVbMnld8geexQU1R0qs9Z/4/6mXurzXKc0Tm+RZrK6i4edsuh+w
k2f6rvIDy6RZpnNd0or3rvobLsgjLV4ygARzsF0P75nQqxugv9rRI90MQPS6wYRzqAqwrz8gXBPt
ukrrJ3ADFrDW7FWndZUAxLkxPCkYgKP50NYsRWzYGhlQ0cj4i0wUAsFOlO1HAptO7tBGLue76SIE
YFF++J0iZAU5iMR5JBEYPCXKGxDH0bgaFuujkAQbXrvGQo/pqlYJ47oc3HmeEo7w3nzTlPfkER4E
OCdfIgAJ9syQ4Ag4i+pFDopoZfc2ClVB4yEnYYrXmpvqSiJMQevoHuOpKJDPVFBkyJQ1yu1Q0O1L
EUMTcHB0E03skWYelgq6XFE2gfV9YnlLLDBjhK1hX+dp3zZJWG7fClqImMuJxaqmVMOeQrdnXPAs
3iWtMldY8egQoOmYNsT1lWiWoBjV+zoX6/Zj/gxxd2jHLmuiN6I0jAsyH5mgDOTIbsmpdBNQ8drF
MmkT6LdFNiKdFxcHPyK7791t9CaC201/1kHrZiY1Pp+3bj+fKSq6bKl9LTzXPLQbaWcMNC1N+QjF
u1FClp6Z1sVsPrMEZ3sDgFycZdRhCj1rN3Yb2Zs46mvmZlImCSryVcA2AUFvaOLqyH4IQ+ino6IK
jeM56cw6mtCjVROw5VZH4eDetELwadxG4+5sOUn0EZWJb6mgCFJ6+q5bcrNu7YB3WWnWftnGBeqc
mJOpAvohq+1TgpzgyQ/o/RtNOJFquvOAy0VqxKneUX0vZOyiWP1PY2iBFsm9mDxv+ItmmHK3EjGE
2gY8UUe+l7y4S8V1+x3rKKB1ICip5FsGK6T1V1oiPV8cNaOo6QJgkGUhRluDLOFukBBefTZ+kQrA
uYenrxi1osTqmY4qj9MoX9BLI9kKtUd97rEvkJY7k8nxicdMqLGca+AddnQTo0tqoGga7lBJ0J49
sr27wcEj5ETp3JvYMNuYNxJ/BKOFUruQzE6hl3DG+pKJQqlOcGY31tuAA4ei+q21E3WfvHHCEJmB
AuvET1nX2bTHA3YHTgcV5WrXE4CBA4cdjCbb+Jozduz4ayi8gEbdbkiFq76b6tnbUS1fs43KEIsk
YZwD1Za2aI9xUDw5BBj9QrkpriIwwZCS1qac9hqPfzh17ug1/L6nNT/MaMriMOts9YLWhQBFK6K6
xwSDbOzheiB7BWjvQcBIHyX2xISnTUGi9LPCFmPb/Xs/cZ7L1retT1lKKSqiwyHblYMSSdygj8le
WV+G/Zq9lkJ8tyqoFatDwQ4U3NN6vwrhSpUf598pfQSnm8X0vqmYCGgdHriKBav1LLF4J6mlIrYe
fI141QMu4rNhToYSzAcvKPBomRK0Me/LVV/91gU8IfDtIznXFpsRT6U7Wbu1l5IAfksl9bkTTISs
LSIUO04LZ+ZRhrUEQUllGLbYlHQcGXljVacGKrOcjj3Z/HT7jraa7+ViEepw7Us5t/xgSQLsorxc
rdgZVUkUJDxoNa3tInwKE1aWtQZleQ1SK4jpT8hhqI5V9he6BRHCHdGXxUuZVx/tFftXn2w56Q77
p9R0xeaFoFd6pdgJ7hV9v9JRuR4BbdiBKYzfbvDvp2PO5aqqfkh0AU3Em2awD7+DMCXBxxTp0GQU
BdysPIa5AOPwvaF45QJ42M6AUhlvAVmOFEFrd5c6gaHMQQLhYcrSW/LTKjm/FuzJ8s1WT6tAqbbn
ac6KF7tRPiLn0tOR+IqZmzVz7QivsI/VxmhmaaNH9DVROo05Dnmfjpy4/xFMM5ksOtSjOf4mu7N4
hcwXUPYyu2OG+LRoYhNGq8eQW9bJoHOe4sOkj0uAl23KohnaO6IyQcRt587FWTGy6YjsHY+4Rqal
ZOxyJH6fuivr1RolDjXdV6OticobVgtNoe+mjgWsc+F4SRtC25/Z0/6ePnJArYbLY48fSQYxwuzR
1zLbjwU/YE+D+hH5k8LHygW+UJ3s4RjD/w6HdGPkQlFOfd4UpWeyfW6NfoPLL4TLjRctWUb/vq9n
ZoOnbD9rbYb7xqwc2RZE+U9nX9nU5lbqfGklCDSf6qb3CTeDdbV4z3hb8A1U+JYACCa/HrgrzeIe
VmPdnnHYIbYD+GZjcwR9a0VR+wtQpqdp9EhY/frOihnkdE+GeM+WheYTKcPhJu6MPJ4LvRhXWw0Z
YEuC0YpBS+TfHq/kD2aHWv7z+02e6kL2eakc0cMAm2gZO4Jj15kKYFiBLIoY3RATSaeNaLqUmKcx
HzNJGtp9D8WgM8smCJIMaHi8+zEoli0EKm6Rd7hU6Cmcr9eykvtWmdoqMbTFertnEE+aF8MZj6r6
iLfrakNYns4Lv4aKX0nf/OpNLNWdGDxDwWvyvvgsynKjVEy/D63ZydTqkL4MY/MWkg4VWsuCysXI
M5tQWJZDOfchZBmjRjC/H3NFYvkOeFS/X+TBtO/Et1wCKvRcish/9/yTp+l+25sI2LCk6Ar1oEZq
VTAO2+AIcTRK0up4aEp0tNx5F70yl+X4Wkds+pcVn18SAK8rAa5zGon8mumXQH07/kQDcXN03szL
GsfqVThLyFK2Rerer5t3yhDXylSczfqhJiWk0XafzlJQ1906z9PgOATj6ZkwKZ8X3D10U2WmNe8D
wmlWHNJzn9Pbv8nduxUBN40cDhhKMyUsOlLERBnQFW/f5BtqafUIC+UDV2UB8UF77ksHaa53gy4o
iYm63+Ml4rjK188Jfx6ZF5EMRDclyn1RcTLxlzBDgtRILtoiW7k42yZrQt70aQmVPvrJVq6SAspC
fcjNNCyIJ0PJz59w/SONRgicgJu994A1OweDkCi4jg0PtHEGLfjuwtqhIt9h/BAgzJpoVFm4yWtO
Ssbmiz3AySTY4KvOFXxQrLhXSaRSzBJHH4/H0esklNuGBeVjWx5QnP7hafP3JeT2fyyYZZD+S3UZ
QP5o6s6E6GEShFWuoqNGLZxtMXJK1WzH38cnKfdLvkfATUQFAV1hKH1UxW1wZkxQTOFCyFavIGMG
WeC5kws00b+idS26UicxUKfce/jqJozns22vtZnGMWRGrgZYE3QXGbmJBk2E3u04YgINaB9NKoLy
FiyIYc4FJRjdja5iLbC/H3dnr6iykkUWqdn/He11VlFvyj7kB+02xT8DrsU4pFVrOSPrE7pYXVDV
qEQQMvf6C/Y4DMDIEUlrcAPYelnWtLNF0DvxuACQjn2y5b+xitI3mPMksuMf1hrN2zV94AM0WzOZ
hlQLVH03pP0HEP5OYiB57yuygMt1jeBmoARg4BcQQm8l2erkF3e0q6pU7K8tHxhd1CZA94GOMqQO
yc9u37xoU2Lq1jqh47sNskaDM5RaiZXPM70gtymok6LV8gYFj8MdCt0fucmLs5MMZHgs1FfgM40n
i68deipkh9yLhrWUZXvj8Czv+E+k/zGaDfW/0n/3U3j7XwShJdCfWtoXuNxNd5VNbPnsNFEUSjMz
MNdIJKKZMCXh2+P30CW6LOPMF+rxqFo/JPBsM4V5E9xSXuFeE+yndHQneR0M21eyK4V47/YGXxKC
aae6BWi1wstJqavgHlb0axdfH0pRvMzVWjRY5Sjlg0GpLUpo063qlmv0GoY0hqiiscumNYSNh3tu
awvGiXz1pkIGoTq9hwLcqryCuPQ0FJdNgNdYxgfy86OdocW8olW9MZJsg8Nw+YhYJSfODBDZ4T+f
Tx3/CQY99+QxS+yAI9Juku5/ky2TLQeWwCIdXgYdXlpH1Sjdtpd34BuFHG8UZRjT15wSR+s/jSTs
0FdOkpFFEwPpynFLFaJDqduvrmFiELwx/0lFzA+eTV2hiaXQNib77ZWM6UO1xoNf3lKhIMK+5TQS
GmhvYlErVwDF0V3OoAWr1PyHxTo/cIIJ53Gca21dAPIea1MBLzQVxTFy6jZYUzX1KtV0i9SbSv8m
dngHUAJBBo+shcxOcAwSjgV9vzrUiUCKRtmYXHkqwmov2yf8SFhcYl7rd7Few88Qsve8i1mnzphK
kC70tJJzOBoa1kxsM5D7X5L8VN4t33L33sfqFdIS8WyH9vmhy9cdGkL5ZDWwnybgFQlz4vJVFS8M
GCHFbdHjA2FM2dAk9yYpTJ3yW2XUX+XN1hxIohu6b2C83ImufAywHbMHpnma6/Z6ht/PcM9Z/Rbz
2M8oTsCQeaNGGCCxH1MSY9pkGpsR1Kf9ZFuRzFuSQVsvX4tR1XVSgGAx5Yh37YNN96yivEIo2gLk
wFqOIdQVcVH2mNiPbjaj1XSFPtXS6T2oqXfRbGqhGLKVGPjuk1Yd5iT/ydhCXiYuoFYswJYp+65i
R6Y2YOVFw64f5W6ed/oId/CiPbCIX90sJwJHGXLOgpUltPlVbIwR+Mhz9HhbeXXp6nE2lQnIGZWh
zh28fzoqVVXnycVBA7m4vCZOXxl9WB/CysNWbUEblsaQ9NcqspdWEcmZa/pXFeqHTmqZT56ueVQ6
2QLrINbwKnNWYYUr053uR7u0eOWVwXfBmCJ3kZzfqZBkP1UiKbBa8nW6fwHE0YI4R9xrGR67R8he
gDxe+brq7tbXXVmB4KBhcXkVvNo4GAbsf/pBZvX+15zWNvDMEGoWMbIlwe6FuDnvR1UdsxL1LF4p
X/dmtKigQ3t1tVjDk5C9Q2JA0k5l/HYeJjKt3mlk0diMGFOnF+Hp3c4SrQ2fq8+f2APr+cM53Kxr
iJrsluGHaBc9COrnm1CyjPE2F2MQ8sEic/k6TB9gKD73bNe2a9Y/laYp9YFFu/FFgRsaqfvKdJK3
OGIOVNChDxratxr8uAtGGgunC8yx1V1rM0smPRZl/W9UAg7j+qOilfZ5jqUZUno39M0uDM1Hc1t5
Ym733sJqlottOvjXBNnpqNaYicdjwR9oT7FPTnVHk3LWyVhzqv71PcruwME5rFWKgrqOKw5ZzgfN
nyl6IZecq6mXwxYRoaN9Dzv0krk5lVaFDcuvipFWc73ZfYkwfSntmkt+PtNsnefsOMpZKhogymqN
ZFu7r7D3KnnVS231x+Sr0Akv3W55X+fZsExrTdmVGZqqMpYoC/7gWEspF7h0O4hifAb89ePQOZvG
PWdmQsUcevgofdrS8h8c1oHMUqcHeiZA07AgWnY0z5My5GL0cA3WSnaT4+DZpWyh46lF7wgJxSKK
a2Oh5CnV1Nz/MAfISKU+wxuNg0zBpc+J1SD3nc02yTpq76Jxo5wDHsFpe4iVlBoGz+qqoruSIBcq
OcRbWkYHYMctS1HZdQm+4u0irIzLmwSxhTinik37jtrrbc4/4lQXXbjnvgQd2mwvxgXFIMKO9Y+q
JVT6uS7d7VTlXC2gTPIS1mGNVFDOfAuDUMJEJbhGmBUoDS4nsJlIB3kotbXEW5nKzzJxWq2VKS2e
31+BMKQHL8qxr/TOD4GB0tL4e7QeD/GOZ5Zdn1aVlTYw9iqMKkFsWHVrPo/Z2rLNqSGZ1vM3U6bA
mM4f7EqKLFz4SK0F+Hb40AAR7GVN0kD8Ye6sin9EPiB1P5ElfO4v6CWLccOfwtX+zRE56pvsCNYj
vu5Ag0IdtYgIm3txWAiVJT6r6K4p5ALRCmQgJ5dErgmC0LkU01CYgdMpkrsqgf3EF3f0GFuwg0MW
yE2QBPvJ/RaMqOGDDfp8RIttJny4p6xCvjoAsIeGSOFYW8BCCkWImmPHSu+zpCftFdgrbCtpGmmS
y7h3QVPyg7uSRaupe5w8ACWGwR1EHMUbDGWuvcBHw6AZ610qId/1rYyjKv7xqK62w84TeYPNZuAI
YFM7UN3WJny93RcCozIIAOFwsSV2u56Z1LvivsBzAumTP27qip6CgyJ5pZ0QsHvMNGYSz2OBCQzr
TgFsf8GJxvJNe2vWqLoI6YM36DBkvC+TEROocU/3XG9yadWG3zjV5Uh01sTBISoFOqVFuVrhFc57
Y2x+acrfFcT83N3ly1Y8E9CLY5QXxtnRVA/29duNFOuQA1/1IZJiJAYhYxyT5Ia1FtsKc21ss84/
0t1nZT/QbUizogfDYITWVw9ehy4VH93X3YHobCRX80A12LHjs0kcLSA4YwQZTcWbkxK793HJymX6
KcPwoBIllXfNmvLfMlZRr48X6jZdNDrgeF2Ot7wzSc5m0dEqnRi9x65TKqEfjhvuo7uFPMC4W/sa
GE2PdS4QDuWQGEl4GgDIkhufLG57bD9wjJmj+roRKSKp5/5XTH46SMhZT7bc+UTttwWB8QLlC13t
+sYqkMl/KbYWBUSnqQmye9gbOXmEe1aG1YezcXS9O2xx6/P9VMQOVHod8h2UFLoApNvMpCtXa+vx
izAyrRA/TgUVLLXaF+d9nD6JiiL9VDCFj3Udsty9oB6TiKndBB8qUkSHxym9n96ebXhReowg+Vjk
GWE07aljtZURcifAsSj4R1BV2ebPnQfEqjRwGol+/DsGVdlHXuFcsuIniPkinStq6poDMaqSzZVp
AgTJERhhKE/tw8T9CKBP+XZcAQD6oNSNFlNGsbkp7O7BVNy3jMUSxRt9fTgCOM3qBZXNErT/qnHn
bMaCPRvBa1mKQb3iJXrTKubjbh9ifiyIBsuLU9/IEppNMCH3pyTN/7A54gqAB3STjc2Kn3A9UKfi
SEhNh4BlDqOQOaYchYIFMguSGZJAo0EyAkvF3gTa9WbGRg5yM0iipQeUN0WwjijBI3R3nxRSQLSh
1QLKXf9HWyZ/Dsi0N5grs3hmPRoq/kp8QyHEgO6XHAykgncHN9gbQ6GvNAVtSsdAe48efVduwEJV
kkojvvMOtTvyP6hc5RECEGhk1vcZfpzrichaqxkv4h//yVEOwdLiY4JnaWej96AweYFB20eDsUah
ayhAQDLBJL8LRBk6yFZJ0tNNOJ61X6+E0jr9CXWORqxFAainifkeXzdhD+U8Do3JxTsOFhN7LiLD
w7Bymtsn5n9uSn5OkzPGQ5T2yZcrknTkYQ7tVcHskBH/OBQoQyfe2bPur6FNyIP4zroStmHNFEct
mhoUmk4HYZuMZDVW58hOvKx31Dxvj3xjmfhdZUzU4KOOYu1CW4d4yqUoc/mJX36DsTHuedjkKpZs
AExQ4GkucVxAvPUxNhkTU9zV/K00/L7vQOJRsN4IO/RnRvzTF9LfXYD7ndt6DK/ITBM2f/2mo3a2
vBqL/5n1LT7vP6ecrQ1PWxipfz4HVqe53qgWDDT3ItKidU39MoyljFSBt0bzzuxmKNyv47OTFtvD
WOcBdEi3lNjeMi9sJD3Rho+xCravV0lY4FLQQO1nbD3HojCjvakHYAae7iyVw7Z5fDcZ4AjaeQhN
OkGX83FBKVoVWFNjs1r7/Xl24dA82DMUHdCUokdSm1cJITPTU8Os2oNNSn0ZPkSNf2hs5ejE8vYE
yDS2u5ur2AyyDJUyR0a8aGMgWGDlDVeSgVPEF+4m1rwGVI/fsVLVqqnngFl9ckz9vHzn2tlZvxI3
KnQG4xthMsBaAm/UNkYhQAENmixubGgS2a495Y1fNZ59Bn1JMN2fRjY/jxPmVcxUvFXjmgwl6zjC
iaGoCe0JKbelgRDlU5mxyusY5ajWBk7JHl29FN42+Gb5dbT71HBJ023iVqmTrfAkUvlljKQHlhUR
hiRd2eT/+Vxv24GHlM/RX0zdZoPWkRtGfZK1R7f/NMGWzvMha7DGXFkiHrnHaIr2LvY5RCoLauU5
Oq293kMrvcNpj2ZyKKSl7AtqCY4lT/jI+o2EhQmJm0w3xBIdPEkGbdp023/03eIJefqCp4qx5aN5
i7PJubyDfFqp/Tlk5zG+bZG2Hv2Pmao460XxLKHIWhyku8rKc3hycuqoTP765434wnkmNkUj5lnJ
XVNN9Fh1MegmW+fL1pRj80RrwzT3oMwC3PQDAxBTSqKVdHFoeCIRSszwwqec3bPijX9WtllJbpH2
blKV3qcmOGp3JtFKbEo/tIcx+mH7OEgKtYGRO5BvIp06N+Q5UX32BZRs0l3/894HvKyA9o20hGrr
M28pqSRVLblvEEbxrcDp87QJAjbEvCtDnUYJg7qfckoYEmtrJ+8n++lFLXqL0A57NnhEFxCxQ1M2
ZQ88/VtfJpvCcyhj+DHXHjQo9kIHhL5MKo6b/Mh3DUzpOHzcRA7JF4Capaq495WKhVlt5OgRIlbc
c7tUklHICsK8dxlNhFq8OYPrQ7UGFrOu5//1JBrPa2ifoX3WFDCS/j3QsqrEOBewARRXZgfEW+ji
JbbGvj6cDjkKx1Q/Y0Ybcy4ELi6hWWh8s05TvnJQB40n9qADRAJLSc5ldNqF2/aexwnP13YHgsnV
Hxn/d2S7keneObOMj22teRZ8k9NdoqJkmgWnpuyrsJxK5w1PudaMvKb1Hpbp1Loxi77aIOS27cQq
fpMaPu0vnLYakSISsPotnf6Qx1/+UvuDi08tB+99NKZjdyeVnOJkbRb3BEF8XNJmK0vuSwVk+20L
30Drr3AC2pxevWBO96l3DpoxzXJJPdjAID540WTrqCkeBKKv6HY6INNTvpr8qSh79zLTNmF0ade8
0WbZP3JMbE3axSJLIdU7XxiBaE30G3dnSd800NsKeWl6/ePB/xWudNV9Dt0C8Nu1EhFol2pEF7C+
h3lnexMldXXIU6guEcogNSnRCRuKar+K2BvAPApTlqwoff7WNSHQgk2XabkVJltC1f5BGZ415djd
soAsqarPzaeZ7Gbui/Lcb9GHGIyr8eXVuUvJyQCBM1HiLhn87aT+leCFFeA8UYWJ1X7dYPGF8ajM
VBHP81QD3+VIBqhMKOwMN0VpZPjLWWRUmTfsEO78s4atscZs8xMqWkv9ih0FxnL4CMdwTODmOswG
R5g5uZl/7lChpIzEAb/zrDMg7/zge2hq4MKGyuG2vorEiau6P7HZPS4qIzYbCkVAG8XngJUdU41c
n+yFA75IKm0OTm13EFlTDzRNIk1hfu4EgM9hgpUs2lZ0kt7Y/CbQ5o21NoLhmh942RwDU41Gc0t/
BIHj1o+uHR5CPnqj+8J8GaAs7jkbbNE1RVV7zutO/MMeMcOtNu4XpRdYGmJceSAggBfbLPaBw/Y3
t4sySKofoyOY7I7I9Z6EALNrFFYYUfQr+Z3uiOz58i8/uKV1hzTtUbvWqlVtaUQBmkn79JWpoP+7
3k4mGnjro8pBoOFUvX7A0JA7rRkfOSZvePjMUOw5uLMgl3HQZV7KPSXUmdXS3qaFXc8nRrv5SFIh
kxArVGUilu20Zi+IZkVSj8zIORKGXbuH0CC+xS6bfbUTMLqk2FGI5t6GcLWFYNG46nK9h5+SncYR
q9mlQ5zk1Q9jzrNkKGD3xTXu93em0fZ2SNfypWux4/iXCzku8yYEBrlUA6qu0CeWisNuDyf/CtXr
50sY6iJ5izq4NXqvIyPSkWOJxbc0ymyjgJ9AF7p7PQe+2E8vYF9D4CAXeI2G2O3olAykkND3TqPo
Jt7OU2/X3gGZ+UZSTPgtXWf5J9Ya+KJ8sLRzHzZhGS0OgUyNa9baMe4UH7PDdzNdoYEzLheHfrG+
sXaFfjFOQhwMt/e8Q+x6HXLx+UHbCcSIfP35ydKn5xmOR2oAnVpHwShvnj5nuSqiZVPrTat68YIt
9O9RTKS+6GEha699122hDjTKvLCmbjJKfbc0lx2tyXMdaQmpzCFYadf/qyzsKl68ueva4deDQz6/
9FMIm0n52KMSYbWmIrEOZOkOBGBU7cjP9RfewQJwO6giF7Of9H7OQJ+2HU8JFQzuqk1gMCYQSKlG
jL53UUeLljdwT0S8KdkvkfFGzaqh5vqeTrsDLjxsk1ni5mGnB/zkN8PyxwNo9F5YGf/Y0YnUVQJu
BOU2cOf1oU4uvWRYfq1P7EzeyxaXZcjqiPl+tAz4GqEZbEwYdHjrQbsN+7MLZjlyPmwHu5EX3AW4
+vF2VVlXBJpwECh+r/97QKDSITtTR88XQah5rEpW8N2fPn/8OclaeOxHjLkLbwgv6QEpRvgSv9gT
CNG+Mtya1zW6JVv3vylY9JcehVMc9/UcFqe6CbBwWPI/1Q56GkPYp2q5qZLMVj3PMebzTrZnh2RR
ZrAlX82DD48HcxbjBcTI275EluOnWD+FY8ThoNIklQX4Op6uEWvpLnkON9a0V6IhmUQyEkE14NLv
uWC04jxnFXvVSPdNSgO7OVCE57sO0iSuwLfsQoawxi9jgTbdBBj2ZDpO7tcRDGCvn4+2uo43Jksm
GX54SRYbGgUepmPxOW9Yyz8SsmJwKXRJ+zgCe47qTBG1iEW+W82wMPDWLNrroxSa8/ocJM8y3+UO
T1Y6ZeJQlOe1M73nhp/yFg511LihJmzV7Nu98lT4xnyRhTrFW5InoW0YGDcAZfAARNnUkXYphnJt
yul4q4AN3DZ0W8JuM0mbnxR15xJNvADPPkX6PkVg3Wqlir3oXrhaRMlIMDJtaQ54AubKTZIOP8DU
4SZUGDglwOmpO8lKSOzFQVvuRWdYM8Yo/54+v6KsAlO+X6rzZS+e4V1AjrazbTOiAYfAfFqDkbTC
E/MGHX/m/9phlsg7ehTsxFntgyUnjt0q4yKNlRm6Zdiuv8d79YfqYLJg6h1k2U8AEghW4l008+cm
pt/JzPJ6pLRpYZpg4uZIsDj/b1BbaIrA0Ir2NJltcsYjZVqcqW73KDxx0yt4YHPXNorcpM1mMMEO
KpHa/fgpaL+W3d9ePRH4w3yPr7i+aoP5YRRhXRgKIO8iesyC45ERY/t8EXUmzlgxSOYB3U6a5g9C
GXKgeDXq/DGiCSSoBK2aINBowOtixb9WonL0i4qVIkHXbWbrRmXsMwMTckeUDAcKP/Phnzg+uLSZ
mP9x64cRFKHTb/AkfI/Euuyf5hDLeh3hghAdzW//fpNfIkcpTAKJABqINbiqBQsdkXwIfA68OW90
O1nQ2zDaywJ0Uvr8KXkOzCtuGjLoioy36iT9rCrrGfy+8oTzzmluR9ehS/nhDzroTsdo+NkysxLQ
ywjRjzrHKklKw2uZ1cwGEdGVjaOdRVWGyjnWu4hwXo+UEIZeOAcp7JAE0ppvOeC8CIrszYL770JH
M/UYW+j9Wx3IYOFNbTSNbVMwTPee32c/ztZziqtlJbzMDF1DR7oTd6AxuH3BpWTZZ16VrYAih5gW
+VPFYP7RS1VFKiH6uJkwCu322Oj1E6psDRcPrnVngL46H5CT96JSsUOAiAxEq2DvLkl4f38Ugzti
qmLy1V8srGg6tEMljLHqdLUbNhxeKwTATVbcDbJYQ7lXRVgvMysMidVv7HQfQzZ4CKrwuDre1M3e
NwrPn/ZXjr92wF2HBaiKCW2cNal9BEzSTwbEHIAel062MtY2016tSVuEiCde3tsppgHT0WqKkIT4
RfATYkGHIgBJJICM6sfDOIkokVwQ3bskNcywOtUB3EPNw8NlVhj5fqDK4awJVhWfbbkj3gsHw2Xn
WSkTlg6O5TT5C+5/1E3NgK7RwQxnkYbXZlR+W6Tj11kRz/ItESeQM4JhdkcrWp3+TokROqLGSWyB
FQJjYUZc+tBs3kE0K/M972CO+gz17/PAW752U+eqr6Qmtc2plL1AanvsYXko2aCgirhA09H4YCg+
iS+E+k/9dPg5drDwQhauo916k/0HzynYzVtMX3N0z7Ej5qS2s/dUVWjiB5rGaDoXobcAcMmQJFPW
UbsFORU2uS0soJHpMBCmXYQg05sYvy6tLOLK0QCGeeb7xfDpcuyLvmI0y7O8vYxbl34MjeVtLOb8
Q8Xl1obsiGcmW6yx1mOAxL/NGV0O/aghBlnIfXbLR1XEM6jtvgsPjL6G1+p2AzCDFsx4yITE8MpN
ZIaShSaykq0bJ0iTFfRgTtNNrjCP9wkTLtIp4Y4hSs9Kbkuiy0Wv8M016fmCh7Cd2MOhWf6CX7yE
wq/6LStSUVTy0oxwJomumU86GjQR1REFx+PTpXo/VzmHTWpIk7/73f6RwJ/ZY67bwJnl87AIwnZf
BBHV15sWTcpCUFVDI/qD2RgDIyZB3W1iokKvZcRSZAFN+al5ojPkSwwqG1ZL0atYc24CKlGqMrBp
B8+ezCqXw5jdX+2Ogu9Lzw1bQlOtnQLg5aJMXs6za6hG+fbM2nJfj7uplDXIityS7l/FJ8Ro4bfy
opA/8N2dE2InM8ZVTo4xHnBbFeCmU2/bPkRBIgfl8VVCcH+E/I6L2JbGadtDNOCTP/ybkJMr5Pno
E3CaxnQqu0CPKCb9YENhhYMJoXQznxto0lJKURdJ9qLsNnwXL+ynQlCKU3EBZoknOfihF8Xwzb5H
6wkkeqgEq7j8fuRWQoQqrpDMjn+Ia1Uqu/sgR6rxwLzvBglsweYQIE+xACFvoy9csZM8US3CYf8g
J1JQ/wwaMjjDj1Z8yTLmh1TwAX6QntfRvruC8kRe7BpwyBHqO80RiFrJEmY/CtYKn8rpmVRoLq/Y
/Q9eahlG/2OwxTr5MZ0Dpgi4aZZPfVwYh+k3kUJUbUQF/CxYl/0IB0NL7rTRmQrOnRljVCQTCh7L
TAkMgvIaZ5RS/PWFdNbcLIi8eI4XLAyXnqc/08lk2jBjyEIJx5qYgYel91EuffawakcxUsAIlCn5
+wvKdOSVT2aLwJQN7BQbzT7dbADu8NHouCG9bdkr0ZmtDS0ku081mILj/e+TRid8ZcFarrhbabmY
PBP2iCevBlhfssNW1pjKcJX0jtz+doGkjQFkXiu1txHhgY4aJVFsU/MMSA8sxGlGuFUCguIl5Fsw
BZ77YTTXhx2qOBvcTUvCDxeNG6eVoB7xztT0V/EYSJVcGEOo6/A2lwNFWuOJwd7uisY2IBAVfCs/
EuDEihiqVEVj6eLvbBKDEY/So1FvCOGNLEI30/wr1S439TY4EPCX4NDqhzU4Rc2mcYSj+on7EzbT
y6jMuoZPleVFZ0GGJN9oHU7RhVliWEXkKcju75qMAzf9Yz3ajgza9I4VaCxhlAHW35yYZRSyZd3G
kAUhVMDGCjzFrfj9/TZg7UJ0Bud857HRg56vUWhzCCnSk9NWiLTBHpdYN5Hx8hzT2PLYWIZZ4Gqe
mCor19Xt5F7Sj23DLqMwVeZ7gJ69cTgl/bnfkaKy6zOYX8Wx1tvST6czfW7UgannysCvjcUyW06M
jocWi+s3eosrDkR5Dk7e+maNRm0IJ8mxpFNtRiMtulxCPhyP8vwaNPmzxYrqKU9ZhecV0AbE1wey
P5ArD9y18C+UgcWGupW/pxAStKS1ocw32nAJXSwH5dIVZtplTFTISagZC3VmY0xVXwA+nUo6zSRH
a/zcE1rBod4HM8TPtsjjLwhhzPEQ7BYUiZ09tXClVcJNnCSTCDyHrnX2r6CBtnj2Aki9KFGDHGH0
9hcztUZqZWwM3ul9hi4cEMbUO+6qTaAufcLjRCVcXjltEnJ/ZQofvEkfESqlXJzmatxakG0KKa4Z
cwwztLlSlV+OohQpSMHhloDjYeryaSPWXY5nNiuF+ImeHmaVt5Rs+ZvwVXSMMZQy2RAzJADgmHAx
+O9i4YaLi5vBjZIumOglfsFhvEMlLWforNw+apjejsGdx6dCNONPwc8i+jsIk/lW8r0CaOZELmQe
U8tOd23iFRAhpVGNdcmkKmWwSbb/QGlDWfZau00wbctSuusZVW4iDOba+/4yFvNouCeNV9zo1zcZ
ySY/woCvfaGED3Lqgtmgh4JM2xzSmgax+1fSj4n37VELyCa71kJkH7UGbPnsRopGsXdrqywv/+Cm
Eux3hvbRsX3/VB9f85xW1ZG18Mv9R+8F70edpSy0p75n+ue7pSbsQ5araKzNI6a974khmDwkJWKG
eK+ZZVZh+9rSqUDMvKmIISOrBpevE/3BZQfsEZlvuxMu1WG7/XO74nom6bRvRFwJHu8arY2UjKmK
6rC+/pPOqFfbiN8eHtpS7avwFszqjMspvSphqSDCV4CTFmokpgWpPP5sFHiV4mClsefNPycZm7Q3
2u6zyKRuA6K86zaMZMfBBqQlJ5G/RgZpsCY4QuIZMTnL+ssORZriNSc7iDSjTm5NmmWneYzuVmNZ
b8SA4I4FFNvWi8WoDj6/yaXcEgMM0yD7L5uv1XnyljgzfITzQu+/0tVkoOYxMClNXCNvmkOdJwWk
fgUITbei5pj9TpKwrLZAmJsPBGIEkXAcYdtg70946MrYPBv5SQsZzlu0TVm/yOwdC/WB4IZWBRSe
OgwV9ZTUl4IOF/mIbFMM7udnvgvOq0bYUCUY4rCRVCKpyK7LHf/rfwiy+zZQPPwWD3rsRQdMRdWi
P1Tg+PQ4OKPgIcnKtda15MkZvRcbSS1vumpIeb9/8NkGnMYv4wvxmBQFOw6imYt57rcM7lq8S+a1
ZADxN3LkxH+PnVUb741Nx9OCa60C5VRIuKCpAUBXU75zLsj2AHJPJLVDmzZUcyb2F5UvJFBVPG6n
yYdo4DlBbOOKPwnnKCEiIVF1MEIHC4A5PVKxjQU4vxfzT5YBqDyAv+BL62Kf02xQEuY5idxXf6t7
jJfZGaPc/S1u6Ehh/4RT+cJZSCudHSRgrO4EJ34UKHmfWgu8ri3OmJ9mySQxkd5zxAEv2JAz/Qws
er3cL+VKdkMGuSNizTagC9U9h6Ki4lptsU8eSTdWUOZd29j9caMHCkTQtbOfoPAHR66t5zucbgok
EEFiLvV56biig1+FDDxASVY9D9Wsz4Qv33w5fmydyAkSZt4tOPRoNkEMQQOIElBOXAzclq+1AdrD
u156pqp5V6FlZnoA9++mlGwesjVqoFzxGEgBVfIENjUOtJiAIdeK5jjY/JUYYHDQzylSvYb8515z
+n8nFs0ky4Rv/0yBCLU3Y5MXU7xA/v9GJI+WSA+skdvddJj/D0WXIpWXofkyozWTqGezBPCTf1BI
DJYJijXql3oFTjApDxBUYHsyu8cQiPcIm7icUbXVgBKPvy5sgqVKrxp+xlVVbQDv2olJeuZeGb0D
+75poMIfi1srzd/3ZVTrPsGDy93VsatG6FERbwLtStTBnHUlIGiEa6aQaKyZulQDVVUQqBMiwhU+
JAMzVJf9YkivbrL9ApO4CDHM+JjfvSknM0lmNlmLszjH9r/m7Z5XGjdh9L8UFZPbuCSV/Q/Psj0F
W+1DnmJQqCz2RNiWZpIvamio06lYA9BHrtDH/8bLpW2GbuveDO/ojkBnS8pGbajHheDnZhmij0DD
R7ugdey948Ke8iYuVKAGBlT8cVevqUKGFVDFl3lieCUbQDLtg8qNRHNZ+JvkHlbq7VAXVWjdyahj
XKo6UGfyNlSgcgoNgPxUR7ZLMLD08sJlQSvHjYMrF2oXxAMSpN2PwM5jrU/EellwnACJI4rrDsS4
B/C13yeTmz3L30oevE6K2wInNJ/Kou/UGrKJlo3nSC7QOUnmSTyfXpvAcXU9iO5UV0yjNfidKEbP
g/Dr+WFEIa3IeVVIS8HNGoNSq4GdHCAV6HaYWiH9oUd932u8XaeoSvUob3xDSkSO/s4XF3qmHHGV
6bO+9QauDYvxXPflIaxHZZBkv9TRM9bx0iTWOPylQiMuLcazvhE9bI9oBILublpRRueXaMc8ir/g
n6HAtrnr2D3pW9NnfVlLsSq3wUcuyC1EwVz3nDehm8CJtMWgOjjNK8kGz/tkfKVkhILCB6+ORqt5
IlPOP6kkm3ION9UMdv8tY9mQbuh7l+HErn2JxLMiG4Nw0XRSrjv5xVwNVC29Kv29YX350isJiDVa
9lTKSffWsLUifm5ktWanJzS0loWlsvOBRMNE6+d1JxC5ly8xVx+Xd6I3RBUvT64fUSwI0jNhsYlW
loqSzvpVCbDoRKmWds1nV7AWBuhFLB3ue8kvUAlApUOsGmfJQi5Ph0lE+YL/T0J3gFp4wV8B8JdX
rqhPxmKRNDbqk9IeCe2Y9P2JIvHAY/hyegbEzhfG1sYpzw3cWcsFFpwmAD1Li4w6wojTavP2/Few
LNdPxXrQMlB/vFLVTILceHW2J44vponU6nJbvCReDtk5W7UBIOXfrMcOF5m9hOy3AgNECdI8xwUz
e+7lXijvP5M2DAk1yEAjB1LkplE7YpcMvaHWdoQssmMLmA+/HoNUDPW3QX24jgfLM84JKDOcO/A9
RCPLAG3Z72FdDrA/2qVSSf52txXd865gr95v+9amjk0wu8RDL24Kk1LPkekjINOnHGkMqM2ap6ct
pVXtie1i06qzAvL7gTjyLgjGLEwhyLMrtxQRacupn7/Eui+LqdiGgGm8KL1UEigG627UoMh671BB
XrnGD8Zcc7GnYOl0MYhQlvuPkWnBWmRYQ2l6P5UnEE0sU/DLk6yG1RIhOg4y+aUvkXtLMX4Oi8IS
YJE9W52APrk0mUPj87vq4CyaAczIqZGoBK4Wlmg0JpmifLuoWkWi5tgta23qQAhTs8Wv6tIv2OF8
/BPHMDtAyYxDBm5q/Y89AiTl/kCLuNaCKZvw4Vbs0hosHABteamNBXGjInih7ZbAeK5zdCDjjglh
hQUu4bR7IFdyEJJ09fHiCjzNl8AM6nisxnoHdolpJLnM4Mq+gYHJMx1wJfAs3atiCOaMPrtyymrY
54c0pbjnZyW6zvzJIjNGoYVBdpV9cigJQzJiCbiBrPijI3APfjBM1iuO91tb97RS7+XwY3AhgJcZ
PWVyDNgaCKatlxDiPE0rD16R27ZN8sTcVQ4qXtx+PJHz0DvfkDEzZ9b+uU0K4Fo31q3IcUcxQLyE
1udhJMVS2SaybkPJyiy6r5LfNrNesWqaaJENgS1id++ge4GAM/K1ElDq9NBoYCfXEdFPc4Cz4XUw
9I5XZBpyJhx9HI1xtBHEuxiws6aXww4eLT7BIsKrv9HM/ntSUsIMUi48hd4mhHvQ3Fw+zOxPqJaZ
tmFrtbOMl5A5yxzBgiBAFgg7K8OnNqS2lDgsmgF7XIdDqcJpWkSAD0jbjXWrRQTEJQwES4YHoOzP
IOhF/nKcaf1+CNIAMLLPklfXcWXLNpdX90WcpxHbdzeMkNREkoYfqdl3X7OIb1TUW38JhvfCRloH
x8n7o0NtWL9FQtveVy9XAoIYzzVSSMkoDpZ46I43NnBmKdqN4XluiLl94PPA5DhLx4qB4bxaW2Xx
DAwE+lM+42HK7XKVB6tqJiCQ8htbF4l3qFt9/w13UrBb2XMYZt3C7RWufamKMkbZgYhZQI6gTNAL
8I+JV5kBUwJaY4yXH50HFzlPCFWq4GHDifnUXGKeDktxuaY/3G7RiIxXNjvKnP2/NJXGXDqGSUmF
HWI72yd0Z0vgF1UZsBRsqbGRSDe2Zf5Z8h+KccZsUHie4sFuoECOlqtCReWzlxKI5Nl8wUrUqukw
tmrYup/Dy4Nr54RbXcwN3CrmDwaASkM61QMux7nYtc/JClqCziVgBguXS9S3k9hweqyQH2EIKU6L
cvmfNLi+BpYwZ+R6Myj9aGsWO1ixLJ14Blzh+5Gopb5CE/IjhVYVf5vrIJSgkX615NbXGBIlJiwu
tE1d7NfIQdaAghZ7rliCgFYm5j30hZtGmQcY61X4zSNZ2XXoW/UlmUrITr5l2eSBLl6/7UePS36S
u0YliY1FlkcQoLHIHBFQJP3moWhFJWsvOIHRCuTPY4ournnHpImSCtgX5RhRXnzZRAzn1bXwDU0V
w743tWCe2hSpV5lNCUq+ucMBHMRgcN4Uw5An1Qzb5Cg/OkwkCnzhhhVEQKzrKMb4W1STxXPTXmFt
5R8+ekd8fB723auqeTZPe98BS+qmV1Y7ysLfy6/EJXSemxHbb9Zi8HrLu6vKXGbiWUNVZZOOyvjO
c/MIa/XZlKEkfvMfMKdZ5OJPtM/AxIP0A+sjt1MYB0pjqnWs2RbijcfszpWj2n7oXohdLqryQuqe
7MBX+dYqbghilxBHsM+0RmGJzBJmFAUVGU3pc5iv0mvAd03OuB/g7B+fgiPNbLfWdSJlhWIAx8LI
veRK9FNvTK6BL+wLRFDXuH+EByNe4b5qZCerzc5CK4FMVe173gO+rlWHJQWgEMsUBw2riF1gWutJ
trxWw+bv8+kHdKpkYr0zlPGnQ7lJkjiZwTFo+ljfavMXbKiXiBHaN/La+dzoQVRBPz0WFXbpM0JO
R89ii+SpBb0O5/V6rZX1j1Z437ehNBBU9CvbXt1QdPvcBTPQt0M/cIxBNY6zlaSHn4Fr/hcyFTuE
xTHEZFsrplj4fZIna7eEjHA1WQTXg7jZHPObfExmtPB7mQFOlX/+eWrOK/gvQ8N/dltLl399OGPq
soRVaY7imVOiDcJquLJIN2wNujGND0BDwdq4HxFOUOPH5LswgCvlerSesk1tYk9IH2qYBu6EY3u2
UtHKva/3wwLd2CVQArRSrw/28eqbII5tYdduHqkbtgA+Xi/sDeFRq2kKhrDJhmW1ApxjeAT0JYMl
HX9EZKAZsSWBNbxi4phyTQYDGbXwkMc6wjHHnfB8szIvQ25w0OYy1mjrM6YiAQeKux3fR5r3Txc5
DKs90Wobc9HWhxmUnuxG42PsVrGZxVkOKVQGcxV9tioAIFPwNyIsDZ97MBuJExIggTv4GHsV21U/
ZdNlNwmMlHYYQIDeAKuPLLdnh9+ymXnZY+EtpkhfXdt3K9qVJyHDWtDiQvEF5dDztcId25nf5r3g
rMLQrAUPK4pr4XA7EM+0JaTqR0WD5zxKqqL5ZeYRxKuctXsPjbd+Y+UCIREEad118bEqe7jSMmcK
J+J+ocer8CXD4Ak8Uj9dptf/sDsz17H3GALFvfm05R0r13a3/3LlGyLVNIZL/1Lhwel5D8ZDoioM
C4E305AngyTfxfT3hTWimwdzXQTVH5Gj1hsMVkk6RpZqr482mGR6jPvvylHIrBqLKMpZoImNbbN+
AQ3sP9LjBT+FFhqIfZhnHnJjkrj3UcyPK8JGE5bffQ/7ZewUA5taEaW1ngKNvJGhCC5Yn6FWfXpk
20imGdxfQ1Baicp7gqhsPPshxbrQY1+H5u4QVH8tO64ZAAspIVIwBdMerakmtO5xpMTIlTa2RuVE
c9Z6ef39g37Cy44nCMLV3DuZ+hhUIIDsySlxk5PSesA205+bJMIDvYfK8M5F1+GNG2lynVwh2KHg
iXtEz4JHaaK9CHxhU+jU4o8etksWIYtUif956Cbv/j9OT/JsY76+73FOHkTW1lDKAQuVe5h7rgAM
jyn8NhFdXWPztNMT24lkC3JOePt0ej1bYJ6tUPCc5gTYos+9lVGFII1m4b5/71E/3myMNig2KzIX
dG5vWVDsS1c/BK4xReWutyAVmVNGnANY7OOwBDehlUg4LmltMlgkGjjb/KlnohNnbNowe4yCtGqm
+LL2C4JwSDjrYsDI784C843gDC3+qn6OutliW6XZEf+tz7f3QQp4W16CwRN7xilleW2fSg89xLJG
goBRGLwX/2ssafDNr83y+hxyu3Vgdf558PCJTclsZZ6IDFbkOEQbE8yJkmDBJL0Uc81hImqgmfsA
A0W7FmbP4bm0ay5EyF+zun+TgYRCXUSl2ogdL4ZHiWGmk5ae/XddpMflKenRkZaGC53fbYwCZsWu
vM8IiqfFg8fOMJq62QVDCoAle0trOEAkgVUiKn/TLdd1hzPnjIsj5PjWeYG3ZFmSj35fA+SPT7hu
2fZWyUwiJMbd3gILO0c8HKET/0gbBE9NK78QPZk+76GMmSUclrmNf+16CLLxGpM7yyvzGvEzXgeN
3YSXzMkGXmBogSsHbqOKb/fjGQE1ban8wvnlDIIOFbQbVPKSaC33TxwWgYyXeURw6y/vRA1IX7nt
nX9qo0nnYYxq57HM4R82GDNlG0COgfv050mSCl8zkbpfevAs8ctZoMuIFHkmtXLNQ4mr6+aGRCR4
C+DaE10ngXB2WRI6V/BdEjQ7EGgNnASJM3Z9Na870Ghn1xZL6uyveMBv2hRDlHSwOD2AfUAqZCQC
0O6/ZjVll/jnAOcSjFS0idanmIO4X+9dtLlKeumLv9knXI1pT5MatcKTyyN4p8GGsjVlKhcWwJ9f
fu2ZorlaElsr5LhTD7DluMiGiBLAjCMG2FZ9Q4Pl2oiInmvegeVdDEHbQU2Cy8z0DvbkzWoAFYok
wzOaFRXhvKGTT6Xtrg7rUEoanI5nBCiYn77uwVRDWJUVrpiCAkXFNgNUKN/CVNAeORskkGKWDmKw
AjQaGZy8RT8KLR3v9UKTQBsQVoTplsDSRbVpQfEulxLAqsVWy0vEhWfBOVr8J8S/1WgCTAbOksLa
+IkZquFUWAg4KHzXYdDgE04CR86jIP7S1UiGNx4MPmPKAumYTuBC9qSsC67QIZV/ZL+l9aSNCLxM
sXU0/VOTOrcrrxqkJkIswtJgtfdSO/McSpfOQZJc7ZvQqPH9Epwoq5LdP+JZR8dTw6zZn04PXuqW
iA0eNXoPExC2wpZanHR5yrnGN7f31jkjSrHMRpgpfHMX2zmcp8bGLvSW6Sejw2UF79lEk/laBi9t
Jjsj0fngZf7cZZzZVjRraeNlE4dZk1wQNHWTwASQnEP8rKzrxRarFOs6gAZWWHciimZfAtczJ8lq
CjYXFSgc22nmKT9jLF/uH+VFaaHFWHC0Z/4Jx08B+6GJQOokCmbX+ZhwycQMZXgzjx3pn0YcEGIr
umuUkwk5Gn48ada4KLSIlXmO9tH1zdTBGFcuOZ6SIihQLQvKd4CnX9fvbztf48e9VQi/010Tvs8Z
gElGoaWcMJB7SGQAMw7w+Ow9Uiq53PddadhJ1npLml7v4RQqjEBe5ewuOdqjBDFyHCdRb4w6BHLg
gIpuVvT9QfJNAKtVNBkexq8IL4EM9hVE032+Z/vqJL5kXEVpMCtqR6FLLOywotyMY6/kFxaPES9Y
r7+1i4A9SCcGg6wI4VPj8tESPdoMR4z/5BhpZwrB73LDsqt7tQRi/u55xYpd7EhhsW5x+CXOgEOi
LZQBeC0qvTJjAAZoDqvCohlDA2eYmwOgdQOAG2RyMtYgThrouI2nkKQOPdeV0ZgqYOw7P0FLvtcC
lQhimLlIc+OAy37hYOo6Gw+D5s+F7qXBo02xQia0fgrf/KYdWac0WlhALfbdhH+XWo8MBwwfpn58
TnWIXkb1d5yZ5UdM1KVu0lB/w4CN1c1Te/Ap6sycAqe+RMIB8NafRuteGi5tUzrpozFxm6d8GC+O
YEybMUiQJXrl/lTwEe8a0HIC1u6Up0S/lYoME0BUPOb+HefYGkmlNw4WPN3LQJPMZSLJTsLQPrwL
D9uJMAXyZqoFCVrHAmYxFpCRmccYLWQqmLqQvXMcvn9obmGhA2FdHvQ9W8UkTGrv7gKiOIGQtklu
x7eWaNVW5SXYeteowCNPGcf51JFRaLxaB3GZ/KtUPkCBVXDswvhOeWs1XHQ8QhcNpEk8pSbnerWo
zDbQmtbouqlhpG7RQnZUPx97ZQB8G4mS0RE+lNFOb1ydjmYTKAaGODk0ShK3koFulSDVnmsTelyq
Gq0WqXl/vMFqcztPH6FDu6JWDxLt9O4QDt6MVx/Y1rdfC6nzFgR7sADVNuXUMRyIbenBB4g59Uhw
pwzYahiM61DJxSGmHuYa6eudp4AoDTMxAzIf5oATKe1AOQ1cMVo4GLcPU6CDXv56NWXSaK4VQNFH
eRRGOB7OH1miKgaciWBDLzNaXjv8No1caf3Tq2SvqqcRDE5KS7DP7pziu6EZHJFR0giZmC7v/G0I
G+5jFDurAkTizY1pnV6NjnGA2xuhJJyerFuUx5sxEkVftZdQqEyQATnCz+vZ7YZFjhhEPbcrnF1k
c3xQC3JU5ogSYAn1CNsliHdAu8KMiZL+sTSX/7lreuWYrxFK0U4hxc0/u/XFXLR4NkNxfhHxe6JM
7gTzlpwNqdHkTdUnY6hZ4PBPlR5uuLXOvNrAk8H7/ICsThF4qD8x5MR+WSL8Z0NCNYTqi7msCmyj
A6n2n+T8wnSsdrQdII5dbXBk0AXdALo9B9v5qa1XiRdciYuNaB77ANIIXNVdlzLj9M4pthzJ1QoL
t/tnP7jZCYCmik9Nm+WnMav0kua4/62jcCsThb69Vm+5CVTLnvXvjrC8tKdH4F+K2eCPcH4azRRK
bHPs4gGnFW99oycGWk27RiVKwSxNkXvL/6Dl1UzCdte8lPFL6+RnPp6nqofz0MzMUYcdHnVZWwi8
uDjDMPTFtMLlW1+c2iaAZZS9lNntU3mbWSi4nU6voCT7zA4mWIBNSq36oixrHlFlJ7j3nOjubl8V
qkkn81aKop+0A89neVovWdHqp9XVOXVu/fsxhEoNMMrT5QZmq+gD+/rN0Jmh6oqjretRNIaRF54n
PEb8y9x/LYe+stmuxD+MuPls4ItENjMZZTUWxYxbleD30KpEkUXo6IbjQY/kg/Q28h15L15HP23P
N9LryqfrGMWU3A2QuzMouW7KgBAb/YyepvYbURQTwb+T5zKOOMhYawOh736bnNrX6LDuOrqtAcb+
FawkH10cXKgm2x9qwhiHYZOyqBZtVS9prYbJ1O51GYV1JNWdcfeR750VB4Sdwethxw6/nW8UR9C5
wkhnkuKgD5bjzfN6uqWbnEvjNfqce7G58+j5M3zkSWEzKR51iA81sbyALKOkjYoHgVTSNBvYyuMH
p/FW5Kkr37euRTgD11Rr9gs7byO9J+lIS9Es9pbIyUvw50wenciZt6fDe8BnabWCPq0ZYOXYJ+6f
t7/PA8GagVPU1n5Ji9lNs5oUs1CqhXTj75tT9fACrQiFVCN0AYR6RaCrIquFdzM/qA/f2kRsfIc4
3DMy2xAxVqLo9Yfl5osnOSLoZixIYHAAa8LxSwW1XMFNGR9+nDjpgw24NDWZoT3zosaZ+WUnEZVC
72exZ/vQo+sxMHvkaVJIss7Y1Po66TDMyYqTOfbfc89VE6LD83VoNyc7rvYnWFaYzrZTdCPOkuTK
DUhxB5L4a1/9QKN18yz4xdFyE+g4yBgpArOTQ7SnRUF/x3eBHsLKUAeMrGlIL+WzoxRm5X3w+N6y
LyuQNRi2vA7wcx+l+VgCSbDKkxcfMd2JUy7XZeHD57QAhQkUETZw75esAfVw/GaN30DcYkCvJ5Kj
F4C1VwkiKHbacERD0jsDfTfN4RM1g9g3pfmVCfpizRhUW2iGRN/ugtAo2Qs85DlvFc5U20ZFH2rL
B7WUtg9O6YezrV9dR34wwB950sh9+1BfQkW2hY6ViEMj4ya3BrfnjK4uZKDE5ibSMduawdP+Kd8L
RkEZzD00XWzxX6uqTuXjb7V33VX8XjX8xX8VccnbvAjWKt0XlQ9/uwfdep/EaT0TsHhreR9rGPiA
gcq1wZHzaL+1RAPF26/SaV5pNIc/K6IVSycOXopIG18UhDQ23Vzf7HzOQTMQmKh1oBZKHfGchtEZ
7wbBjdVUxmbY4iNUMPMHbzk0YzYdLA3qPIo7NR+Okd2mUHbN8GjrXDkO4cQJO5GXIT71/QvYmyF2
a9zlXiYAbn8ALc7a1lPGGLjEK3YKlDV3873gBFabU8WGRiEOp/hR9R96Wgx/SVFuWVbt3TyeWWHz
HvVzJJ16RB8E3P50B0BVUxDGMjwBWP2eU9oMgDNpSUl5cjYkS1OrAUHLDTMklRLvPnIBn0qk+Qbo
/QZ9tJ7ASjj1XWUiKUbDEETfcdamMY5gYCZVTvtj/LUtuDq7Uh0Bn5Ry9JOgUdUug7O+vBXnzKGT
+bvd7CWe8fuNvji8XPprxnZn8R4A6tCqfpKKIWl8UYdnrBovE++zfkvkXms+MVYVlPSdIkCfUjws
cDUtf/GXHCCm+cnq93iWact7CON0mdzB/cjQbPcqcyEgDQ3UeqIxeFmcUPrqWW5TLZ5QYfXwsAsY
VO5ioo9KWkqeOuVzZGSHHwMJgd9Iri9kedjZK1/13Goagho0DieKXQ+A6JyGLi5fZBN6Q+pZOHRj
qnsycPqCZ9YGsH0Ot2MjH9glEEwFeI7X4TY3VNDmYlCotxKwG689WACSbrDigBYH310vhf30u2WS
GJQvTg6YydumTsg9yuqgme4AMW/+J8uPKbXCC/gDtgq+KnOARNvX23Gu2odI/jzcfsLsqLn3LXxX
LPkyPGTUKHC50bxbEavz7J/8q3r+XvndQnNikuo9nSqSMJF2yBNCA2gaCoUMIhuT8oyUr0XVrd/q
wS/YKu0Eu4C1daM4nk20zWEwEL9hJlg6fvcb/d3N3JqOaH8cegZPm5Fx2U/csIEJafkkUVJ0jcob
BL8s3EOwn+O5xPjqWkzrzvLToiI+n3l/EGDeeD67IkNZW+QPi/uRhYEclQPn1sqqn59JrgNUg0RL
j4XPw4fP4YXNHGUVMa3jc6miQez31V78jNVExUULHWvOGjrQCtG93DSG5FGlFok/bJJM7gUIAses
pyvQlK7IPjnSxxtmBW/2QbGXbA2G6gf+hn6W+0TtNnyCdOKLh5+SEeMZz7Ylsbi7nfnhqja4UFMS
j5sbvQyJ7aQloR63IMeVkqAPf96HG0cUqJDFJMIe73eG5z8tb0gAMJLuw6frFzkOTSScO5xUn8EZ
tYVnjGW8TA7FRaC3CUIc/zpHVp1LDTp277EW1+AEzIIzYQjXALkrjZfd0DrLXxBpMNtb3ts7WUME
4ZzidCkF6zj+X7Z0tPqMUgg/38wK3eOhw1u3/0Vc7PjWxp2jrPsx0A4S7SKAp9nEeeLxaDsdyn7X
9Dsb7XmrpVNOkdvJC4c9Ag4dSa32ax3dpfgcwTdrth8H0dwaWXZb4xZ8x+ndCWMaV59iDATrzIYu
zuzEb5A+1hfMzPoYX5LNu7VSOqhIdtwKk6cUdZzweLPspnUAMRe7LA4DoTR5PPyCxknaDz00sy0v
oPWX9/FBoTBtuVmUC0yRQFB6QYqHd9T7urJQHEsAUBPnk8TvKHBNB+uz5iXboJ/hx9E/n02X2z6V
E5UEm5AWhb08BoRLzPDswCysc8p0cly3QwSf9d1Acw/sKXZJdogkU36ql1lDI1Nwg5Myv4Q6b0lU
1nat4+V0+zf2cDSUdUGDtMha3LiBLFZYRWOlFH8wXQuupqYAa9/zWDT5dxQWDKJTCtWCiWngRwFJ
7n8vRbVuud52YGgOnewtC40ql2Opj2MWOEzaGgFNCQEDLDJMZeVh0e3cbp01EGIFOtHh2Rvs1EHi
CDvg0BngJdhKclWHbJvQMjtmDnIdgwHRdGcfhP7+YsCmSn8G1A2ztFy/zR+wo/xxA+YgZJOclZjd
uvja1nKzbhCdezV8pb6hCrUw1wOkNhsW1W8IvuaPpsKjlskEEN+TAOZRa/271sLSUXsjxsNLvrm3
ZEGx7Y7vqp11YQDDJuwJnZhQ4tTytqwH/s2lr5JBuMh2rqFLQ1ABHTIIFkn46TeftMcUc60zSv6V
fm0rAvO3eQUCOkVSKfiflUdYudpNrJ5PZxEvxH9HSFQ8NfDqvKTJ7p05Cm9vjlJ9qBoFxLSXZzr6
hH1bQCf+eiXs/iYgiFAhLugGa/bDMAlKCtUo3gSeFvpYDivd5BhoTghBS+zZd1FBJyPghxoVJeZm
LurdQOXKnut9FjFqSdK9n69YPJhbUUqeYLQR94brjtR7p1RrGQ37hmY0ULSREh39Xndrh7e7GwB7
LoBGsyLGj3OWl/mQdjTOAls0NsWtdtueYs0+Vo59QEFwWrZ4MAf5AUPjJd+ZrP2iFMx3uLlLFlSw
vlegx9mXL7tRHY4aCc8JMlzLx1yPVlIO4y90FN7M8dB25KkQ9RHhE4eH67izr4Q6KVqm8truVjVn
PHirJVcvhDZXye912u8GpwkFdCMl6/X2Kswcz72ImUUut0N1rcCjdIaOWoGUSslrHDJ0eCRR/9Mj
UoiLw0VBh70+u6RbLeJ4ItBjh+8yf5VzBlJvDShhN2A5pz2UIXAviC9WM74NjzR/VSyqFrN0WetN
lyh/dFa7OogvJxf7dxZjNP21N+IaHM4dyrFr4tJ8UdjFqy/a+helRYJiANZTG0aBAdGonIBt8g5o
P5J7YizgK8MgoXYE2qKUCLIm+yDES3a5eiufZYdkO7DrNYNkHKGdveyO0MKv9xSnr8rQbtvc5+Um
x3zk5ab7E9fQNtRxMRhsDx7DLrrA4xYLoo+h3b/wndvLLl5/MyiQMyOGDg7C6n5CVgh62qWeNi4L
9IMGeHFlosaVvAoyPYua2jxRL8FrqNvGQO0TmoUCBhyTbTWqfRWdUWQRuuboS24GbirYCmcDuuIy
YTK3SE7zSwBDEGNicSo8/j3hD1t2A8e60UmC8V0PR497TLXJyLvrk8qmEwfR/d77MT5W3J0XKj3H
L35AgdGAGGBOoklUyEVk6RC6nHRY1uuk180AU/Q3ln2SDFpyy71/dgKUG8/L5RSj4FUeoAKKzQFK
kdrQFYP7JtYWxGEptloyOo/TqVeh6u8KQcq2FvJ3IYLSS6f2+g4if11Dw51bBTx+PbgmzQo0HxAa
TsKblfbe0FjCQGAEk9NgJzUrYGTLnUD6LHu/XtME1IcIHgn59VLFbS2DRLRJ5i+fvx+JfjX1ZBn+
4zL5y8AA8aAN3jvT444exM2fr0TOy780oVyr7sreQNHBMNwT+JWM36mYhtre3ztbLyJOYmQfulAw
fOWVpJLJ88lnTv3TYMSxfJyM0VdYxv60OCFqyKqp/CzfOBdwRq3APfk9WSZAjggUzV9NebRgxPxo
JWfbp+HjYY7vDWzeUBDElcp1ddTflDqA8HXxuuKWdrUJ3WxoWv7CqMx/fu3dXz/LeK9NtWbcriFg
k/yB9rXB3FqSqyuLt5g5f7TbbIv9nPxgBHppPO7LOXwipEx1OJqh2rw+zVK8tYgMSHTZC1KsU1XX
an3hX4FgmVjvHEu7vNNM8mwK28iVyBO3Rw8A4mOb1ARmzFpF5mSCB/1uAM0aGhHf4wcoShLXCELB
7dOI509D/C1iN8UN9rRrM4cbnAj9/toOSHfamL037KUFROzACAyKKt/gHUH8DA17eoz3D/R5gksd
HmqAfEyxFc6VyGueVmx33rTmqpghn3j5GdDk6Kan+odB7lYgrYw/borcRQQt/C4SK1R083+4ijlr
8ZWk8B3IvEWqEOsBPX6ghHYODByhW1eyieW5KiWWlnCYeNajwucrkTmYwl7YYqj0ptyAMAQxavTw
W2SzFeOdAkgYyDCQpFDSwwzKw4nsI0em6BD6xwLz09yentl5ChkVHZSRx5Lj+QnhAvli1RNTKU/w
UQPMW8oOdLvtaSREpaEIo0F/Uirr6oycViQn+bLS03uqJJf1zd++H0NfhKORaMIH0KBNrYMTyV4P
tjMV3mQLhsnelOUjdYnlr/TINF115GKfJW3JQsoHkpTkwFq3H5hvKaSP03/MpBGFJ4sPr6tM/gLG
zyTzgwUbL0pFGIp6LgSPoK7el0vEu+URy0GwYrNgQqR8uwm9ajC7rg4uUKZ+DC3ooW6/4YpC3cdm
Imj4o/Jo6V+5ZkblT5+6nVw+pdrZFm8SBuFKZLPYKNj6uwO4tgCi2T1tOywrU0hzVuvd83DZFTDP
TyUhi5zL3T2XQy1MCtbosWnN6tmv3p+dOWF+8sTqHCMsixxcGg7RHojJ311aPVi6ap/GM8+5hHDs
Frvc7dqua1CLioD5/V1mNNQJ+ikLXB28jAgkWD5aLxhhYZp8rciUqHVsJJipW3vhFo1kwRK7M2Oz
VtixK/1aGIjnAdXQx0JwKcMFveVdErad7qfzaemkj5mJyy7VOZSiNfFgAKBj2PZgcaqG+NCvyF+n
r09DJELQ8XKA9ZXRqq2RP2VM+cbNxfSFBGO0k1kWo7T0Ds7S7M9k8k7aMVDj6YbBATCJu0UHLx1w
iy02/ihRwo69yKSftmmBa+XL/ujiTESjrFOGqQbv6g9RmieAwoW4LEB1/k4Pe8D/LUTn9OUXUO2I
DA97AK+8B6bqXrNjffZvfiwrzaviqtvJ9JOTncK/HdE14YNeqOefk5DGB4oATeREaCjlvk7T575q
H76m0wdM2sXMhgsfjBQAWKUzUlbIESOmziechd939BbxFN1Syse1DDAA7IZHngQWGeC0uZdX0Oe1
q3V/pwAFV0+xiRAtJM05XswYq4WwaPWNy+fdT4EeK2r9KUHIumN4Oj3dJnR14sC6sC9ZVPWtbY/A
j9IIGDIqeXupb3UcsKVwB2gtyWoXN3b/bFho7tcnVHbrPK4LD4yzop4uBu/YdUEXo1O7PZNf/YhU
zeUHmY7zAaBi69Umazft8IRTCD6AzTX1xNOD4CfmhsxAzEktl8lz9fnREunEzw6ZLMZJHZegtVWG
bRnpT1AW3gajjDNmnTYjMQZpGIbkXAO9U4cOCV7WGecbnYF+/yVHj6RLggV+HKIiNRh4iCGjLEOk
CENnOkFWPohtm+zkoZLBMe6oL81asko9xxmxPF4B6eOns1sGkZonVMc7OyyX7axKCN2pkQYg2QRq
0NBIkU41lozSrhUWs47YhGHj7rHMnDuCV3dEFJn23qNGrjoLIH6IDyMRnPQSlXr7FjAoc4YjPmJb
02hPiSQ0BSg7A6geZtsHgKhGFoh1ZDeziMi8rA5PgHBJ8mSBbms0ZGRVq6WkKeazFGE2BFL1S6EQ
ijb2OrDobFaEtkh2dTYc/+gAwtEUitHx1vAdLxYlW57zN3e1EwAHIYcBErHZgaQejmGlhDinlA19
t4nWY7OTgAOSl8GLk96yqC6KojitmYe+uvSwt1Vkf926ZdA2oyo8VHG6mnq2mAAbM1rQ5KVYxBAC
3XaBVCdpJcCMQtxd48GqXsKN6ibMOXmVXpWnHeMsA+2gUobPy6QufwGd/fQt0sSyFbz8EbUc1usB
6t/FOtaLu79Gfqtv5/K9DCwRlWejVdoBJ3nO2k4bW1A8hF4JzFilW1BlWLPKjy8oWhJxD0+LukwE
h9XTsE4lEmH95Z6jjLcchyaSuMIkhDTUM4QHLv5F4O/zGOuzwfIbBu0Y2ez7kOTISs0oRlbpRGDb
EDE130G4+EXONbpcRsLYoRWh4kGXcQtx/HTAWgKLxi5iYvehUdaGcuWaO2VDN7bw59JfzOhSmcgI
Z1Q8hZgRe0BKFvxmLpzBbZ9nStFkKQbnv/SLIMR9ujkNT0PFo7yBHSqvyHL2tHBT6YQk8M3PrE5Q
RlL3Z+OOJF2EQMEPYafzH9jSrs1tm7sD8E2p7tR8nXxe6S4k8XbXQ3usqE2qdwWWhL8ynAgCKfzr
eVf23sg6EoEJjwsVkaMHBa0OB58R/PZog8VxMoucBQTUjE9t1cUD6jvcvFoD42WVqEtiAr4KqPYx
4pzs8HD5/3kZGrhOy3QhWELoTi7ofmxhPgzX2GLggjc87bkTiQri26gJU2I51exdrUF9hydCml/q
vnIhgSlTZE5iDQC7oRPXCxcOhsC/Pc9FEScOJv5VeN6m8ui+fCQsZV8EQA210OQIYKDOqHA9yxRa
GG7yP5fAaM3pQ257EHBdQAjfLnLbNiiSiVKoMhk9ngnZop6VOjVjv6hWJy0Iecj5oOm9tuzwfOu0
3VcwsTPOJxZxjyAoIhdX5CAKM2nSBxKbeQfZnzPFa0GtqEVeX6oPL2381CP6VQP/poDSVNeNNvwp
YoRzhv80WdleU946CtRMFHfprHIdOoHebkQE8rjGLaJlBnj21kj5u7oGb3RWdBSPY7GBlAwZb9SS
xvcNDwFBuFreZ7rmL1Sw9sROhnGFwWPIaHKLaa+/reS2pdVDWxB2uc7NtYWeeE+tygbCdya0OpcW
OKPk9K8IlWl9bi9bGpXRsWlf3MZoj9CxfD+ZcTyErojDX+BKlRLb7KtiM0HVgJ07OZ4By5SasIZ3
zdtZvpel/VMb9kplKoR+CanO1gf7NeHg53cVsNhTxoT7Y/nUBoyhoyUYW0NDWMiS/fUvWS/lHYfD
G/BAy6GLFIMb3VjaAGf1dacp+D0us97N3o5i/9desH2HaNxY5CVybsrxqOjSE0cEAQEiyVTvRpQw
JQTx+9oPySBKqjBRgPKx5TKeJf6Y7giDz+EFD+4vuucMp5phuC+46EnzSQrh/C29Gg2runOce/ia
g6ns4Zq7/CUAp3R9kNGSZ6lgQ1sr2xMVtefBtk2HQmoZxLl9Vig95C9LCU7pOQQi21GhNtHjfgYT
K6Er4u0rUcCunR04wkOR/Wt4Da5rwBDHub7+RO+UDYwdHEr9oWkU3fR5JfdK8c6miBSBLXPwfs6P
HeMy/b0gPLgyufWN3zRwxr3hTfA3NqcS5/RtnCmc2/Mq9OtUUwtXijke9psMY6gFFMY8kJzskhi7
M3C9mfEJezPe9S2Q9jmILjKU/bjLUqgQRSCCEhbERHGbW7BZDJSBJeGLqPlRZOEoAyefnpet+4tl
DHENQ3Brk7P9Gpwr9j4BPYPBIJXSbb5KH5CDhRBvtLg4hsasPyZ8nqWqWPEBRF7hhyVc840YrapN
BAtbVg+2JsFssTr/2xrHssIS/jOIe4egfAf8J1k+zSIov/CQAmIVihu73KbaxjJxitdMHbFudZAD
2JfAhYPVNRGdRleTA1ZkvnGqlCkY5d25KCrzKEkfNlH473zoDuMRHOuAOwaJ6Usrzeu25gAW149M
kU4CdUI55RVP62wodbrStV9NkrdQJntSU86aal2WmP5eMoUxblTuTVDmRNWgrmeY09tAUt7TFAJx
0ekEr6AhuqYbEugFt+4914lGLbRfrWDUDJHy0hQ2SresGe+JqLPsSWf3PD5S3flpxG7Xk8qanVHo
jw0qZ+MKy6vVYp2cjNIdpO3+82VNpjaidz7Bys/67frf23RnIRHiVy9QFrbARoRUICvzO6FfR7+k
tmuKKhuWLpIJBmAXYV93Gqwj/Wn5g5PpOv9in0L49beel9Z5R396VKJh1R5v5p2ce6mGnuDqpwbs
+SR67P05QXot+NZL77SPP6q3Kd/Dq6uoYJ5fwBokPHYPEO3Ed5DB12xZy3nEI4hUa0maQ6l1PYiM
VLisGiC/+IbshSi4MT8XvF3nB216nKa1UeclXv3P42AfkROzzUeHkCCelebbUN2p6FeX7Zv5qVwo
A/IsNKiqeFBRMBRqu5gGfwBtvwQkYjAEGd7/IzKqnB/1I2RqRFh3hsGZ1PeISQlmK98TlMaVTluR
GhvGHYoQ4AQ6j2CMS8V5uSAMGI0YQORvhBjsvxfHNuvxc+CLUYcj3c4QM7TiejQSG2Q3TSyIRVQ9
MRroIWxDSvcy3nlXjdnn6SnLKQaCGvSQM0y3gfEYo3m3IKFc2F7dRYsEjv5plK8Q5eaCWNFp/qde
sJ2Pe0cDmCWH5JiWokOdy1VTvb+ex2zToPn8ocH9rtRCC6BuC27QgRVeHfbVLpFXuu0wnQebrfit
b8drEcG7XHOBBQOlmME4rhISSSEFmWatusrJq5lo0pGtFcTTNYgiHJLnYRgzaosAvGGbOFssQutP
2qL1nnQxmaVImtwmN73e2rzVqjJxFAVa0RLFrZiObz36FwnXmMVZp39dBkycWyG1ZgY4gSH/wy9e
hqF97iOLJLHDFDG41QdaPHAx6mmdpUokTbpcDLQI4IoBxDHiDDg/eDSzSKeL8gpayF8eNl1dnbAm
YSrjkrbwZ6uomeO6EPtma1bCQpCjjHKxCnjvjpyp/R9ZcdRqeWIzpQnSFidi5n5X/0ns3XvSkg6G
OBzqlQQ3DVtZD25oTG7gJ+bt6THoQOphdlH6MVk16T8OT2IlOEB0kHEqaGPrkQBxYOD5DNfmEPj4
EcXJwgbsCAoMWWJ9RHLC/FdDzkwzGZT9+b+qQYtfK4O0dJnN5Pby9OiDzYYGJAU6vnYSrsTwXTvr
/t2+Oi/9lCwLPQ6b9hxDcKJH3IVgAlCI4ngQ4vLr6Tm8glk32j27knoqrgCjPHLmkkAnAQ694Nu8
chaBjqYqm96QfkLnrFIUAApNYboEdDcEWZPBnX2eJc1KpzXjWujj3MxtYWY3pK+m1CxR3/2tXJAY
r2QiXssUp5x0LH05ZSXDA3hoDfcSPh+bbcPaouHsGcU/fqFrOjyn803vnFVSSmC/or0z9pYshrhO
fJ6kEeMdn9YsM9atgqg5aQYloSq6UKmk6cEPyamPyHnpdujyqt+CmHbNhalIFk2bYbHtYV11zczh
4Y27BP/yJ7cHxCEAlfdzlDs6TMa4P+eW3hWS6uUQzRgTXHOAHDRt3nGpUV2SavLf7n2qjJ81aWVk
+Z9EvtMrd/tpzgzLXyo8E08+b5DDkvrz3JrBm0L66AxR6szHql6zCoQ4B3TKfQkgzNg0o81Voqse
wThvsAeXZf9VoSpIn61k3Vfbn9aFvR3goiCTgEZTIw52tniHCRII+O0o2E4wRHSpEB8Se3qrkR6u
nGzb6nO2XSEwiF1/vnb1gzjtnouzDHR8zNe3OU37oDFn8ZaV53r8dUkr7IyGSDC86DaHcXryqLeA
C2LQrpSgCLsM35Uq3XBbg8ylNzWn5w1WkjhuvQLWdx9pPhGLZmM+Iab6nVbpuc8y9Dh6sfppQmaG
dvCS2me2USm0r6uX74ru2bsrTysRlBMIN6Dyd9UMWz+wVi8D9MQDvLnAVLPcIgBrr2G9+M8m6qR3
3B44EPHWZ3ZqqMIMTl6OsZ/oLt5WKzNvHpgVN9saaKBc85/2WFqxmsHJMEWlNjkj/ICEa1oT5Zni
fbJmbLECohmcqJ9HLbaooN6aCUIiFB4dG7FVtYTA3TeeFpnfHvzX0zAZC1KnsIrOGtgZ4HGNIASb
Qb1Db61is1JHDr2tKv4wcyuSTYpdKnNSAAGVQDit9HVkXn9QF+2vahvgrdOIIaFpcCw54JFS7609
seGS2V2rmRcllRCpBb4IWrYDA5ytwWHAciDMV5Kl9dGhd5qoIKHFNBjhOd2sTORRfYMn8fsyrGNi
G3DnfrgslXE494ivrc4GdGqLBgkv4lVzQfmou8Ii+zLbzo3cX1EDdxGSd7HMG10ogejhS9PNHpvP
tNcuyO05aq8rQOUPDXIk+w977j9ddSoxTfbmYJiFbY+RSRcnfLwegLwBPnMIOk3e+efO7RW3l1nz
Gi00Z/uNAlDN8P38noEZBZUAK4rZwBvEXAiVZcO3xNHz9LdmlCI/Hcxnvf4pxNvuRaCzOBmcvs54
hRB6WHPKD5oXG2LImjl+Skz5jCHGi7j6h1Fnyefl5lfZ9axd6lbawODozBKdHY4oFerZC/6IFjTy
Oh2mlut3989f0eq4cHw8hKSGw8t7KiLk35ycPhm14ElOF31dnnQYUjWbmYFfP9/l0vLrg8e2dTm3
Z0QdPITtH/1n4h0Nv16+7XcZU7EheWZTObJ1XI3U7UioQykZhzcgxZtWoTE2QQvRz6ILWj3to3Qf
mQnM6UwMZb+fY/i/oLhj09djh/b9I2m71oZebcRISXsuXaPQQLZ4IqVn7L8jXlxv/67hibpBXraz
hd8qPCNjDhN/1E3NhrhmBsnT81Y75+HP5I+3owbdXmwQzbbKyG1+crKf82J/uJcxumRuliaSqL4U
RCsgP7tUbIJ2fFfC9UDwZko37VubISbOIF86CTlRWnJBBjTCnd5UAJI7PGYqTchPawqJ6lr8ooOJ
vMTjDEBQX4gb/wASSB7cb1+frBn/VVSzR+ZweyU9GxQIVb+mAPT/vV1iOYJqLPDyRTCf22BJo+9i
GHZ8xNJnFmtdsYN1ZD+QKnBvmyqF6vSm/+23scXuLFP6Szk3o8uVgKp3SbgiJbV1eTjwiXafRz3g
pdoTCWRgwM0Rol/Wy7yLEPhvrHakNVpGXqFG+stqnWm9RkC0/9sBc27GtUy80KV6q6cw2gQWEysk
mXGFSlh1SAY14HLzWdLsES4U8aPY2LvsTSHVDoW4Tnkzo+ea25RCMYKgCNoZC1tEZtqc66A0x9dJ
Apeo+Kc+HEGHci7l55+r7lcbGdDaM9V54MD0QopgY1vbIWPymFR5b1NRcdeKykkOcrPOl28RLFIm
60U9Gz7E2A2zLRfAZtqz7IULdjU0hkSABukWUJV2O5BqY9oHHOzNeAev8dZSjdAnfvPP0i4RReT7
NnEVsaZDNfNmzIBD4sTppwcbuPA23p6wMP6EpmIYBP+IF+bF7ohrO8fw5xtIZ7DaGNSJoAY9rbZ0
LzOxUXszMnYWJEGGrj/FYIuVVTn5hgo/X9RFtIVB8yNbSO9uO3HNTLmUP4p9ayVlnsYXI1z0vVon
mjgWFCL1Tl3XsF/bY23BN92SO4UrFQSKfkzzxHhLvWY47K/1tn4S1ALoqVjlkRETAHUjeGhzuebf
SuozOgqgYKeyyl6Qf0jxVVSmci2FFq9Ck8RSCoUbel1CtbihBLSd89UJAgxqKS79JiU1lF7DuEWv
gaVSSG/n0HOv9a2vPgH8wtUcMR60h52foBxd/hzVdatHeHpfHpD2wbpqV0iZcji93lcBPlAt3U+L
XVrNbZ8oAvfu7t/rKWDls8vnXP6pb29BMuK61y3ZnNwAL9yRKSJO95Q6NOSyedVpKFM74nMblA1z
xi14i+1tr20bUAVZCl1uRYXiNfeSlUCKTL7axvP9+z1ogwciqqKHyWthw49ZfuWVYSzJm1by4AWe
888oogBxbyrWRFghuK5+UIWEgRvSSSUFnnSK13phnWLSsXNCe6HWglgCOmUbQGR8QqI1H99W706/
Ovob+z6WpP2XSb/cGZp6DCN4CAnDiPMGQBrQFDWOcWKHK3ecfduEVhRcJDdfBhoRFTWFi45m8BOZ
CvaYYqTpWsrtSC0NJP5IvmOxeOjTTZNvu1Wo0aFcngyjEix1vutDkZfKlUY0OLQ0nPsuV3CgkEi1
p09eeVG25b1hU0FfYu6Vvy945v66lJMxM8mHTcaycGZQw429SRXd6LIPuoylo5Py4/iO5AmtV4dj
fvA9kzUBL3zfPPRe74dMvWmsaucIpIyNEZyqt7s+rf+rR3DXSTHgqYl3sXHtQIII3ob6KCJuFI1U
5X6hgmVhZS0JeTL+Y70nOTfZP8gqQ4BS0DL7EFtyBZRUDaffmSUs/X070wJ2ZIQ5yc4lctO3fdZM
hRmzyZNdI+72JF95BqislszyY1tyCu02pqskwpoZSHiMBXWp9KFU8b8b4gAeq1riiluAzAzm/fXh
3wFT2T7fW3spWQaAyKwb2EwSPXT+FsXgp7ndgUeV1kZCulRLs57y3fzVF2ywfLt9lLSWWFAPVewx
+8W6lNsYxljmEmNc0Dgm/wgl9eXeK2ad/VJPaeRrZM4C4apvsL19FhWnQJDwzO1sKqZlEX9NHQf9
qDomLGXeWXYdRw8tv8IK9cW77KQvipfgRm+QQqFyR2DRu6Cdhn/EvDjUb1kNMGl51Y38ZjSbrMe9
hlWIMByqGmZjEl4A/VUWrWuMkUFB20Qv5tVuQ6n1l9dlENEGIhyl8Cm7olLPdpZM/Jy0bys/Qh2W
bfya6WkWbbdydK0FGiolSyj1IoSV0myy/dlWqIv82/lHP0eHZBYSZx7zrxq2/p0AYqM3rUgd0nFx
IrlGC7SNh6RYr10+jRUEpSdYPV+K/Ev6Y6uz/CURXDiMYQAt3+SO+mQ5g5iyylC9b79ttsfsJG9y
nho9gZsXNojaz78YHIpuKlVjrv//dGk/KrsOB7UUd6xG2R5c5Rwk4mT9/ns+o+u5gn6eB59xVXSw
5CncHe78YYGMGua6nC9kLToxz5iGSBtaGKSKEg1VXbSw+jUNzpze5newAbCNohean7OUXlJ1Ov1M
2piiCXH0n2GnLr/rvhvwVofQmjDjcfnNewnXeOVUrI4czczrKg5e6mFiO1fkm6rsIhmJfFjnkOQX
EHaY9i3sCW0Oa5mx6vfBc5AY48q3fYJzXlwvQHy/TCCwjR5bWZ1fmOgaNj45swh1T+9w2Pum7wBP
OpmzCJjt6zKaGD7JaQkq0Dkn7uVZmrDdeN41kvCC8nUKY1EuWlIHHRk334PwyS8OdmBB+RQgBE0M
Y+k5KjGSwZ27EbqtV0Du2yfvmhLvMaGiaWCLp49XAur2QFA7IAp7CI1l9/msMu7tRxqKDKFxTfL2
LR3or0PqyPxTbA81TAjHy6vEl7P9KiQpPSSPtD+TFvn+wUh01q2wT/+Tmwe24V6bzMig0Deqre0E
Sm+aqzeP3wsni1dbsh6hI8fepreBAIt6BJSVtREkMWEi/kKd/HomC4nd2O89jlyFXmALR9/3z6rm
J4hNq9/KdxOLMMmdYq69U6bMfQdmqiZjOf22TlS9EWTI6JmT/2z07D303hhLiUmBB3XPn/kBmcIs
C6RAYM3SaI+jHcFcR8w8MJSK/ji2AC8g2jH9ogeo1UwuENPklDuhKa1US/Mf8kDRptqrI8XLa6th
URg62hIbEIJrAWhK8M7vVUK6wf+iaNxScmpvY9t0aQSg/CgbQt4gbARmK/jp432qSLBZvdjFv5Sq
lDlzBqRJiA8wPxtgQtiAmF78pslie/WARralcHc59wpjD0L68oNeyLPLPT+upuBWXpOC/tksJ//+
/gcJt29TIr6URoZFtaVO9k6Tcb7FgCrov0czZxsoSjGBE+YeqsSpzUF/wcjRcxXIvUkNh3rfT8pR
o96ENRT8gWb3vC28ZEM8AMlUSzmPPzsgk2lo8DxXIj53LG9v80RNo2l6Qv9cdmVKApOml0+Pfo7E
QbLe8US8QC1ine1iDOJZtfYEWzh+wCpbsdwfvnfkyAtSBXs9sM81A6xvONoLCiaC6BnZ603wXJMz
y8dGgLdqc6xRyPu+JRpAV+cDx8pJQ0JTe/osxoEquaHj/a3s8qngdT7bojPCioNqmy+opi+f9brk
2yH1x9JqROS/GliP4niwLBz9Z6sh3WwmXSE5+nkbMVAFYsJ5qLU6FEMorbw8JYQeRPuk/Ee/NqyK
5opYNqDiN8qF9qFCvj6I876tnYHcMM+ersUYRrrIFYoo3Hv7U13Ot3WX0z5zpXDrfDa2KQ81wwP7
BwUfGidnkmdF2ZattYrk3qpXUEL/6J4eTSzyn/kqntGXD8NPXht7us+YKedqLKG9IljBFXTOuHmd
X01+gf4HtgUDMRb7tr8bYq+P9jH017a56RFSCMogZ40wUXgNVw1IHD+kuwlvEqBx3GTBitPxjAUh
BeGtXxBNJRqbnpL8/iJlyy6dL7KRinSslskuX0bl01HZVsicbhEzFxUJZYDI5YVYgFa6ExqFq65l
ULVsXHWDTHdyks39rDLx/DKaDyKVCJ8deEVSkFJkcRR7rGK8P6EAMPmZgXDRRAvf6hwg5Pi9BW2k
yFrNE/m7ubDJ9LoLo+9EqAvrxk3djiTn4fQ07vcSPmvup7QGT198VvMgV/G+/YLo7F5k+c51IH1S
RkcYdOgvP3dy24P9VV4SfKSofrxeORbpo1nn2XNcINl4aUmWVwFcECSV0PWd5JzrhXEy2L7K2fCK
ZHNC5XqA54vb3UE7lXaVW+e4V+f5cXGNann0DowIbjg79yM55QN+yaPUHnNO9aDSFGC2evytYx4B
VTq6cossQzVCxEMGzk/ZXBuNQV9+66fyWLa7+5/CSNMcUE6idIAJgRLPPm/PXxj0hwbMy/LxkB2N
DfO2hNATKu/YdCzh8qpK2WA7ejGJLBE+3h6tmnfodNi0N44aa5th9fKPry8w/qtTGginJcl7eXW2
XsBOTr5jA97KSRWgqBgpQ1AMXtQF3VEZ1US5Pt/0aN/oyGk7CNtWCi/YA3zou7byn3fM2Ek+CE0T
EMMR3PLUR96SqGNY7qpgpD0RrXDmT2nXIdlpEzu3ed8kg4/TDMpeR/KjY49k6go0MZ7i4JmzSrGl
KeA/Z2kX4OmgFMDKNvtXO6ofrNZ5HUnhqO4O1MN9WVU0LupVDqZBQcLYzs5ieLtUr3R7gGfSXxGe
CHZ6TWcQNawpc94a/rNRGv+IWw/IQVlNDVvYRRL9d1FcBsSy1J7alFdDS+4eVuSZf2RWFDCqoyZt
EEjrD0U4x43ruSUMpHqkvwyJ4togIX3CiygwHWWDGOli8efeSTInJ+wp1f+lW1STwRyBxqcJQmfO
ooypoUm+fe4FXC7mDEf8fLQ6W0tdXRfz1SYrOIhogDOrJb2FcLqGHjRa+5inw7ogn0Nyh8tdUcMz
kWEzRN6vl6was5PmAJroEQWpAwG5zAxckwcTi2BqBw5X1vGx/FST/DW92PnYiieCUjoZc5WJBVGu
rmIMzjhsFFQR/DnfLySGANroTQIL4o71c4RF0ZTIphMQyPsYVF2hy0scPTOALuovm1EcyyRtwuMb
rnqSYD2J+/4DsFlUcgeVMPCXheT1Th4Dq0vckhVwYIfQa4pLkx2C/7Fh0jXBxKdW9GEaNj57KpVD
Hg8DhrPPnMdualQwwlTwMJF/xozf3yQUwBgHE+ua37ClRP75e7wlDjVbQsV7BwLzJWs1GJLrZZ97
qvtiArR+eIhOpWNzBpeligZ1Hi2rmKTV4xemAtPtmb5rXuq7VnJpmxo1ESFcQyIGuXwBQED7mO8J
DfIDwk9vBeAnn+hIrMDzhCQZQF+keP6x9Ja3QEWt7Tnwha2FYHFZwGk7gKGOy/AKDeYMbhRpg/xz
/JUHBwJGVxg8hUUkkl0O1BAeqnLs+z4z/qLw8kRhCE/hfY/O0GdFnTOBZOXTwC+qXrxeZ+R4ol5h
VPSBKJFmIiEhUtYHMOySLYcoZQ4ZxQBgCBf/F4Tjw9M5vYOydtXSlhmMtXXf/duDpVXOYHem2mNx
+/YGzTc1FoIkG9kECY+Fj9psMgGx197jDqHw9pD2qViEtiIU+vOJiLYMinmgF3FAXcLONGB91X8y
yfZHylzfUo5Hz1es0r/ifZ5MCIlRZc3UBeBfd+OL5AmgnNyEmjyZsumDVjKdyiq15NSaDsjUvIgi
4ahzrkNiAWcTTeKR7Q2ETmSHz4tv5KxBW9t9l/kd4efx9qsLXlKDf/OdD1bZb8Pa1f7bLpaEGPw6
gY/lyUbnAILhDe9dz2uoqm7DW5B+Q50L/+48K4dCo9vUzll1HEe+v4SRh7KCMUB3LD/n+/dMCBzt
OLIkZVmrZ+SM/maUDKvqPp/UXBMCkKhrF/mKXGOvsWkN2ZzpCwaOX10kuplFPgWab8ciEpAg6ruI
6Gm+W2vbjPBEO81VrJHfS5+LYyF6AEydPeAPhNa2kP4SRwvA07mIooZgqKhbIxkXcnXosKLdsQuY
XqnOdHmOCsZpDLBf46FJuoHGqvsjZDIko8rdZEuihziywPFMrmTuUFHhJvI/VKkqTyfzikQbvCvP
kzTvA3l0PaLO5OoeZ6po6itRszB/UXguHX+y1shOB83OPxev84PnC7KILlkzmTrFnxmGJ5RZhS/0
of/lGwKbWVedPPvJXoWhUlewllI2sKIkgMPnteEJ/dg53eQmdbXLh0x2g+W7HrNsAMK0YyJvF3Ii
GAAWJ6BTimaVy40DfpzSM+f/lfRLPxs6SfIO7hSYe2hGS5JGiDGYC3ko8knGt/Cnq245m7AcxD0O
xe3d7ZWiT2R66teTbz9rqkyJQBYo7unIQmZcPa2qI8cy2po9SA/D1UcL2PQLFan+l8d5eoeDihLN
Z1QOvA7/8gCcbvqmObf7goirAfcPk/7aEDlzoLw29ovbOWWkZyeEbon2nRXtmy1701VbbgOh4BG0
emdG917Yngva+Fsn1HVk/IfX1AvK5C5StdhAfEc8M0lSXPesz1obABybbqboSpUujW2p1v0oHFSE
QAC/5uMUlGrDeRu7XjYPcd4Vo4z2l/WcR143dgMlhSpq1JXyXJ3zjqZKY35tjfJ68Is1VfLCXV1t
GDyR6UUm94iNmQr89oCnaPGwPxImIsWo1ujikeXZLzWHU3Z5S8TGER2iKH1hGJSs1PYl/cqiZGSD
5l0ffOf5bD/P2dK+Z0Hzeextuh50cv8sKlIAqrI/4yUOQFzYobc3j3faoA5OUbuKmTJ4cyz8ZOMd
cIKq6AYpE9B+w9FxdVt0nNPqgv2pxVHGBycdM7UGhFKW2UY2qsqS7KUIs8BfqfQCy9KZ3sLoKDMl
4RMoHbmXZ/mZf/8v8cL+D87WgfCqzeJ0eaqA4XTYRE02dRqVN6SCAsLZc9EvrHroNMPmDzStA3w9
Sx1nPavJljpJtx80skGGsS9DNvBaSUXYBoElSIaaNSChY/EkRXgi7EIsRmYj3iK4D+Tb8vEtvO+R
hU0eMDL85Ki3LNW2PZaf+9p7ISbQuWmGrbga29r/zGDLvKAXSVpf+GCV09PbK4GAAAhMPjHULTWf
/iCNSf8w1ocWqbAlaCv0BRIwD4CycL1AdNDATY8YobOuIgKpUWGGfDfE6Q1kXLnyV6rzztZRzMGs
avynuw56AD8N+cNDFpwhL3LhDMzFsJOrI+N3l+wWmWM9M8KKoWlC8p/OymvwxkGCH4fn6eF8eSFW
SAxAU+7SayUw00IfBnZS1dhu6FPaLJ9726GTFhzMddAU7p4SLHWa2tVXq3Dwnj75u3oFl2kq6oJF
au9rs9FN7LIVOQiPfK/4eZx04W1VHDcNngSnNcvw8BNkw5s61ihWBVcOhuA9Q/oYG+MDGbXrruoN
InlOCqT2iSvqw7cfn7OOCW+MK0c29FmBkQsDp732WpeI6ieVmCI1z1kVqh3/hQ0AjnoyHPl+fSxf
SyaANRCcrl4vmjTGxVWtOfDb8YaXl6O7P+bGXnfHm5pnhzNjrpmaWXKuw4GOInEf6CrMraoGBDMJ
67OdRrkKQQYguu7Jh11wiAavXDB2TO812amGZLUjSqZN575eDwk5fxvqJMa7hdsiC6m2Wkxs+EfI
0T9UEW/AK+tgD7nOqSPjiN8eJEBY+1Ho+KnTd3ZsdKk5nBV/zw8RDsyYZ0Ay16qHtW32haRCgx27
vy7sL341YO5llipF2x1kOMF+pTFoNMBANQ6tqPahxDPtrUP2H28PPJzZ22WK0kRs/jVjEjsTepse
eAXEXCpShVd4zmtmkzxnijNXKxYWdyvsM0zDZT+jGeJ/CDQzKLlMAQITaJTVjvk4pjf48XQNT9b4
UVzFr9oe+6B4NmSrWBeGsxRTXLMNstV6XW2S4SjrDR25R+o+TxcHrUVm1IIDeCHvq27uhPsEsgcH
fa0WMunY6ToyvtUNv+MCQo+9L5AGELHP3ArbZKHmTGxdDlF1pqZTpGwAYCB8xINkRc89wH6EaU+t
dCOOoKNM3PtsXBPstNzSa9takZhpz1e3Ms53G22SrokGjoPSK2CY2Bls0mPJXRcJpJBMQ6OuZuxn
VHLryeOeFpxkQuetil/vxs89tTdKnVA6TuN+UGdc4z+ry1MvF9xP8jD79+tKX7dZOnEl1BdViFkE
WeVKY6CSXVPaeSL40NOGMbVM6pat8UC8pOZz3cM12Z2btztfyIQL7qsONLcLSyPe2n6nX2LiQg49
58O26mLvQcTa0ljQUe09aNd93sdFr08wHLv79PpMirE5N8+6BmvNwpTTa5ElcTAUQLEHjbzXzSZk
qbnBjlsG7BZXN6DrLDTHMj6jTEOqmHShqIT2lX/28EJtMi+sUBeUu6+BdWMZRyjJ2gzxUCUDh4yU
vWybQioPZTUbNkEgTGDDHT289bODm9VNicMyaUS9qoOabCYWB5jo+SLEJas2Jwvrs+UJA2rFLlnE
dk12VR1gHmCwFV6LQi0RPeLk1ObhUowiJmifxYYyTnBQamKTmFP9YXPCoDZx+zDrbho2WQfjWBOO
AAIamtjI1bFkYva4it4E81wcnqpfF0Yz21FKR9T+czNMOCAwjMvv21dFqUp64yWIs1r2k8jP4XOx
rcx4IVkCrrHd2m4zXCAEQPUvg6yyAEi+PymJ1FIuaw9eFM+N6S6QHzBRH+GfcG+TkaO1SAuwN3Wf
cMDzocHCiyN4g8Yjo13Hk+0lD73Q1oMn30TAmu8r/5Dn80bCz3c0PNiqX5zeD5oetKUBsZryH/kx
WAy87Iy/s/dasfjz60Jdf2kr4C1WJNu14U1sVcc4zkBSmOJKHidZuCPOS1gob6CoFjJZQgZa0h/o
tHzHkKwlFeOMiMYw8GagN0XpbAm6Twdf9uAMrEgRMPGGsBAQAEVLvnQ22jQAUFdLBUYOwHaD3HCl
H1wDeYzSNS27Tlnz9krT+b8yPflmM0W6CZ4iTrQah2bFHYtMqHKYc7itfV7fBecYw1aaRklJJwd3
UdHbtNC37YV8StTA3E/Fx71NGdUsAvt/wVTb+PCceldy0LcHT7utlBJdmXW4ZOUL56m6bTq9OcSs
UyoVW6Q6HDjDDl6Ys0E0Vcn0XNBJvymgt7QpyTj2VeAnA8f1o/PJNnaURuLN/xwATzGmoYcgHbUQ
NY+hGCXB85dmeBMBzdjvEAgs34gGh//N6jaGc3Q3CXe8uel3SAsZ0HBpC48Mr+va5Eff/TlTVdW3
mSYxZeuH3UBylz7GGxkQq66JmtLXg99t3+Eryt1VzPr5N8n15ZFrBJB25CgVI3WY3ygEQij1/D7O
CYZDWTYPULy7FLZwdpE2H4WQOw2tgNoNf0T7zyPcDCsE6rEjM5ZCuHyV1aYRd56dKDngKtkfqLpT
VTIQfVdtXrTqK5hhS/dyX+vmcTHkD1fT3jm6aOQFZvdcGZBW/7hqfekgsf5B1sbWWWWv3cljdPAp
cOaxQ8g2b3iK0vy9F4z6yHFLIclnHeS/+KD8ymwILFHRE0+UyJW8qrYtU3WDQ4ybkOWDnFgQR4aF
uu4edeDyvBbpnUGM2JBXcUrolV58RTDMJnLU6pffCHkRt0F+RFL+Qt6QNvg5v8p87wDsE0Dv0+ud
gk35U/0iCwb7uzOjdwBkBw1sHhbvSvFoev8EG8srQcPlJb/tRCE1/DPtrBrWzw4zHorlAeAIJiSY
eVP4i906uE62JMP7uNXYLGvc+DS227UjjAY6ecdk3irHdy34MKTHNpdaVvWP+xqMQ02wGukdvK1p
TyrcGee0vGor1UNYMqjlAX4ZPH41YRbpSrPBG2y/QL+5WwoR8QVTUw7gFdvvk+lWbp/z6uStdRwV
PfCk1GNGX7a7xYCjXF8Qu2PByvMhZDIf9M1P9Q0YMs1vXyGqdtQnJN1iem8Zq6ekXTndPdPBZ/oa
YSiM/lCx37Kw5jcI6jxy5XGXsXnfSmZ9C1imA7TXu2Xs72+HKrSuNo4ZHQI9VqghoNijiapqPbE1
airdEqHpHgStWjmGTe9wFf3Zooa5dcbZX5NjEeB2gTHakDVTEV76cRp6ZD2xT85BFZdnRA4dkreF
7v5Df/kBQOp37FBhsWPl+txfHmJqj3rE0L86DHvserlvkzes//6bC8O3p5iHP4Q7heHl/ueDMXgV
50NvDXc1UV7ZuKHlK31PUG+39rGvVuQo7B6UF4iG83i9tansCmwjveZLI59V6yu+FoJh9ItcLxKS
txh0jHKdnL5LfMvFCG6tdnpdgMo3qqxDyaHWmGhIGQkvTUbkqCM9TBoO4Cz7fTm35/n7FDSMm64W
m2E4IvAdMuoS+RKoJYa59rgX0PRwdqTVyGHPeYYw6sKZvaaCS5CeBPsHIPcfpSsi80Wf+EXt76lj
jzCwC1YnVkz7XUM1y5bI2M3nLiPQ4Su5ZqQF1CbvMAQ7CVjo2q/hhBt7RsceWLWwmS9hdG3mt7yh
hIDf1l+BhxNKdAT8aBFGg91mieJ7bOvY3jTMpTK1ldEJvGXlhaGZUDffDdaZtbK70N28hRCnafRK
7GN1CM1XEYvuB3FsWViEeVXKfB0yW9fTQR5/16zYixvbrUHn9BDPe2w9u3keogBOB4MbE1EVgTjF
RhFeCqksh08hj3YxaEaujxVagbONxH5sWA3aVhFjU7uHA86xJIYmxvvhAdXdCXH/511redqoUoH5
9bW9ktJ4dJK9+T8qnSKBGkKziWbvva+ZeosYRZnMC9w2kUbjqO87b/X4wuwLGfBrNKokp5odH3bG
lqQQYtThUZYQxkN3sZSbygdpAstZotyJW72jeaSH25hvJO1VEZ5a1fToIs2Tqdw/At4nEA/oZBYU
v3SAqrB15KUuqAcG85d82HeFCsqZaXV+qC1QBhN1EDyAM+VQHDDlWDv2FWJNvxUru6gmS+CeP0Bm
g7cNyzjIR2ypQ7RuR/0gLjcv3uxEXgbdC3IblVlcsIBvzemgZ1DWMGt1ZZEcpjWQTa6IvjiuPdBV
pxWcVSHIB3aOIg0YxrMqw/DZ/+NA2k+dKeyqx9o0pIBA4po4LM/DCeS9LrdyDv8s6daGJNBdCGiJ
ARr6+99e2jhR6Crye+ONOqbgvYBFbu53xQIf3AweMg0LVW3cxsY7aOK3tLZnsFJts0FWWZrerkMU
wbuxVKkFjyRxaIF/OtNAh4acRxazmsf5OFHOZDH6l+jlfsZJO9rcMfyW1+iextP4WT0KMw27WJyq
g1owqnMWMGKCasqXQOZ0jN5EHVPxXSpnxYc/PVFNhH64zT3ccCA0i5Q6pN+/N2JptT6LSKUNA/Wx
OsVEZlh5XLcCCqHGrmGOZtam6fimsktm13pG1Z89JjK8kiSEW2e+paFMuKrVytf1hLBgFBGFYvVI
QQIIyAFy8p1MqkvW0PIhs20OYQGV7us2DTromeUo90bWMXI3IQiLoZTHgKSYOasJqhm1f0wf7unK
Qcxb+f9IqTn+jNfJfUNvFGJXrTsutr1O9N8C2tuOhQVa9Po2v0R5d6TJeCB7spfULcPioaAG9IWC
dP083WJ5TaiQEV/0jRy+REPv4C6HRgo6Fh6K5aojhijuDxEPy8qZUdGFen5geLzhtunBqofJ1z1P
hHfYS+BBtueNupIDLW0QCi2/FdEvDmEf9GcUnKxMXtZPuF+zJMBZ6N6yzZDs4N7/qLAgtntZLBSh
/vXgb7nEKNWpdQcQpmajrMT3/eyfl0v7o616oFoDovLdG+UDKjDNtVG2bdsZn1q775S8II9QUhcq
ESmthtn9qIwZOpvqMgE7wocE3sxv7M8F9tYD9J93K8kHYo8GPliGB5vcDWSSo4AdOaE2sWUdXF2I
A+G9N7X1shPSQajtOfCljRuUDEEkFXD8q6uKnrGCEr2QlVQLeiRS0xzzsYi11JjUNQTjWhbaoBaU
miLXtkd+hTu60UgA9IDwaVCUOBiPzsc85ZxzXCHh1aeuABB0dYMMEeuMAud+qxNBY/Mj9YVQQJGr
Q4KAbGAEenpncfhA4tmFfZ4TiZk4/VVhBnJrRpDs1YYLTRUuEFcfX7S3grWUjjO6mK5qWWbFf3lS
f9llXVZPwZSugIdp1NJYWEHN9eBs2H5Spvp3Fv9AFI5Q/TW7Zl8JaeTnjYxgxSgqlxEAaTaw4KbP
DwkobCtsO/1kN+E6nLJGQFj2YBiemNEOqcrQEuo3NTtBH7wJsOHemG0du9wHkCqxygb2q+4AnxNI
pzkg4YRvLhN3uIwH7VQpye7BhWElOZCp9uid20Hly+fSdq3jHxncsEzxmMubUtaLnsoSIcN3+ash
GusvXHL5/qzx/vrxHUETy7BsfTrdqz+L97chW4UnsDa/1MrSH8IeJcRQBv8frtbUrn4eJRmTWzvl
KpJdVwxBmCnVgOuui98ZxsqQPyKQqww6XkLs9P7h2L3t5jtHum7PFRG2+cHDy03YDr/Y9zpG7Itr
2LuBA/vRuvHJTGtnRpJbNzE9m+1Fs8nCB2NGNZ/LfcJLojx0cwy3fNGs+JuoddCE7VyKIXkN25AM
qbOKtSDHUPZd8UI56cEbByg/zcWoHQPZvi4bTmUJRICsvd4msuSAvx6zanNU9f/XPKX/pMBz5m53
Xt+5n7zrEEsMjPBi7L7/e52iHUqdmalf2Ag4xYeYmSe2KAp8fN2dGJMwxAHL+W9cpVp5PtIH2YTO
Figg65tRFiuJAvqKc1dV9asiFenZSfQa4/Yviv3i4cBnnYHmVwsQlhVbqUyTc19oaHXWOQw20flP
8vQtf1pZwIXKZozPC+3xkDRW4QG2KdrEGwDo8yjysABMBMoq3mxnjClfGErvTYtKE1jHWg4wNXEY
UMcPmSlAdfehT+jyq0dgPonQaLQEyfwAzezVc87/Ee/dHS+p1pxFRISntSp2dF71DRbH/lzmQNJD
YbVagaJMvO+HaIKgKw3903aa9GhzBosZLOOPfYesPsXTjdKcO9L+HyK8TRVtwjEyM1uoYvcmyFoE
nBt9doLbLtz9GC9E1VRIqgS4XS3/R8XZ3kJnBJSdOjO/6fmc+8acKMqcQXXMMno1/SNOyAyJKbZc
VOH6yW2UxO39aJ2l/fjwlfxK1XzttL6VBwxBLH1DvEE6e35ZWeWNKyTVaRJ+/9hBLFPDRawZ1stY
QjYVhDoLI+mW7VSwyxBlciAzTrgcEgbQTplTMuP2uALo7NFOo60U4M29UzmClujiommnyIMFN/FE
BS3PcvFDP5jX8aHKUzH/YkeJfh1tS/+7cen/BD4xymtLN+mnOFCSabzJRTQHdXvtAsmDTRMaIVKa
YDvpfjZq+w6BnV7DE19BgmmE1+q7bkejEkv4DeQZRGUUiseKLPhDeb7ZKMS/oa+byBb44R1Tg0jF
QG9rOIegPQs/j7BmikxuUz6a4xU6kwXxFnTeIZB4bbmX1KuUaT5LfanYfjzXLFmtw1VM8M7il5cy
VnEwTgK9BOyhcSar0DEqagJp8yq6tLLo9KQjtDpu/aYfnXZ81pbmke5xn3eVquy8Dv9oyTUQTEIW
FSbY84D875B9zFZk4wpasGX0dOxT2YMF3RDHnnu8R5MpU70I719YbdQA9eTYVBbX3KGR3nh15pzL
jh9TKf1puE0QcSoHWRsdz8sZvE9uY/LfUKMSXumWQ9QOCjaMRdMSOajBBOKxM0bJShWBUD2KPmks
FPMNqasvDXlgPwxRD7J20eD+DaM08ZJCQM+5BVcYISnes5QvG29HK2m0iDvTURayQftOYOddaTmG
A5hyW1j8nRCUFXPmPxe6W4r0eQWvWH3J7y+klkgm+1jdhYrWjHJWCkFpRyTEaUj4WEKJH2UplNzo
Ms9cyvVSEEEV+Nzt/9yvpEPQKvTOMONXYg/j01zTh2CqhEUSwTO80IWt5LzlYdyuny8LLjXdf+PN
92oiX8a6ROETbxE4nQb6/ggl4N47ZQOIVBEV0BLqM1m4Hptj5Q3M7y+mZbgVHS/94qX0naXBBlqY
yP+WXFfhXC2/wX/z+b5bvINVS/NEkwh1aHZNufJjXJsiCR63mxprmnSuZivGji453hS4QAMxbb7p
Xy5Y5jZFISDi2uEdVRDUhVi8CLf5DqlwESLplyxP7HJ8DTfjrccDvm7SytmQLUKku3WMHci0r5Rq
/50PXH46smvrfFjo4dDWLBC2XSRp4X/qGwd1aBqsaMMk1Ygduy6V5UcDmER9q6THurkmJ5yLeHrJ
KDkQwkxQGYvlWk8jM3YKrdioa/c4Ny1fzF0Cb/lG7hDJ3TUpuo6T/aPeE/+Rku95HeoIbho67pBh
36nJtAJE2gkKzo/2aX/NhIpqqf93kg771Mdn6UaciBidnUUyo8vifApxBeTp488UHl2gxy+0uMGY
h38po4KEOHA6U0TDCtBjY+LyaZybxYRMquf78617a0zwBN+SEAJKNSDMQ8BHaj2vrdklK9ompwnW
0NP9uIkQqeQn1/YfXbhod7ssRRnnD3eiiWwV/VGbZ2k72fmubSZ7vtbkHRe1sHzLd+4M1gRYEeuT
B+cHjXLKPtdHQVOMgUy6fPrGxtYmBd3Pxh3KTPnI5jxlSXPvCPhPvBPMbksqQU27VYRBJOPLOLDa
84pPGU5A0t9BM+zSHi6PIVzQfSs6HGNI7er+atz/DiK1Y/LgZ0mgATsy75XaQWGvOjQGi2PSuuHC
6wYIgUH+rYJAWqUiF80uJVpgDgSZyTnfsG0nLjbPmd6Y2yfRPzGoaQckOrdO2V0lXDchTSbLvjnT
f9Wu6SshJROMzui47c3p+7J1YPVStoCd7yrwgCIPeVm+vx0tUH3PRyeUzaOXi+9uTUgkOVnwLBxK
uhM0tAxk+/1p/cYXEW6NwukB596FK9aRQ7BhKCzFhPiye6iU/qo3bketAzn+wXSbh5NREFfP8zGQ
i2RVPrKyLiH+ap8cDY/aQ5EDDsIZlbxOE1a6K3C8zNOZ72aiZCwVAJZLFUYgMcP2qxnR+fkWmthr
73E8LVQNv6enOMPjBbZ0iZajUTUMe/j/sQKH6sOM8Sv3ypYOl6py1KoitCR+9daKF5r/sxpAPFkl
gsNHhpKr0PVBXdt4ZZV1qkkmbk5XTzF/PdxmKgoffaFGFvZU9o+OD9wod4p9pfh0lcfI7f+f+6Ri
Lfkrpeolt/eyS3pvqlS1z94OgR/XAIavFgtG7D6lsc/j317dWk08jhmm3rotSmMWCZybDlPDB/5d
Y+7PgXWpo7VYiiDKvQkcb600oK6bqecXT6/Troz6H30fg74FGvVXwtCgyupADfusUr9ip5UHnHSY
oyyXBLNB5pWrbxo9Da1gFjse4ztldc98tmfBkQP2i90XBrHyObW4FO/GH9yQuNOY1TUOzx0lJOG+
rDlGb+zUx3B9nhtM0/9Amnfyg0XfZgzQCHZ/EzEH4WP7HytyIpYQDakL+l3gQEn/mLQqnfXIdeP/
eFY/tNKLx4Qv0t8NCWpr8JmoULRWhxyUa3P776btZYm2d8UVinK35yNEmhiv/v6YEXJ71bIdviqL
iXTD+X2dOPXahEd6laDPCWbHeQ1BYdvCKIIs33HjA2sJy78nhoyvvgvKpF0+MMU7omw3DMmcnV7o
Jvmbhg7FyjX9PAHxKiQh0Ztw+/1ghhKlXt7qFqBWbKejZeSV4qOqZwf5KDccP2q6vyGuSmSvXLZz
KgtuobSanf4gKWgqQr1ceBTbDlkbOeTG0eb1p07x5HXwNndOlztqTKafFaXHmdISfO9u8izdHKjt
jZHyTt8kszpdU0ACn0nTvOIL8wgk1vBwpUBd74y+mXb2N8q7X7WXFWeOCXrB0XK0TiCgwX9CCmOW
asdFyXOn09ROwFP54weVkU+ic31KMVqFLKuQW1vgnd7UmuIu4bhSkXEHxveUPIcgIy62vghvURrS
Epa3AAPxIK7Y9+ux/qzJu0u9XE5WIRlwf5dDoIgxcxd42SDkHdLAppYtxbPTxpP6qNEZjMFQSdwl
HNSsYBzNsHDrfY6/SPDZgg/Pdb1m2zRKEH0AV4hKvRB5WTqGyCctsM1bbBk6WER1c3LWwa+Tj6oE
UMF/VbsOBzwEyii17yFQY6dthlqEHASF6OPRquh/e3YY6128wUiZ9ooxGdmIZJSlqK3YY5hHZdWg
S2E/nkPxrr5uUruWVVoNwTEfeK9yjm+KaE9c/vw3za5VQJkGe5uMwBQMD5qnpspZrUgzwXAjk+LP
6cVkSo53C/wZCt82u2t+U8HZ+lA1Rc6GCFR+K6GBTKo8fgK6FINpi+wXueyNAt0l9mvW2L3kiZsS
SUHUxGIT5iEytlAER2+m8sV/rs/BkOpOwW6ty+1JrfmC2iUq8moHkJSeNkbX9RlXSXMtaXlwDcrm
HW84aNHwGWu0gFMNXw4wBHXdu1hs9bu0EHEianOX8rwP1oRC9uXcIezdhtTODTfDINFgbFR4p5HN
uFOnGpblBMQL1FQEtyxvpRlrx/aiHx1cFW0avNp04Xcln47868mwdMNLHkyM6JbMONG0UDixjK2h
0Ryl9o9QvKgfosFBNOolHwnEdpS6YYmHY7h/kI8ualWJQL9Nx+ysUBtqWOJjF1fRVFs0TXjnhWOr
7BG/4d6Xx8QyXVeexmGBsgzgt7z9/Ci5XaOpja36Vna3XBlM0A8Q+zvpvwYA59cJHd6WLun6HJGU
Y/mQtcaNwYUsgnuYKz+i/MzquUStKwum+qwHxDUPlWXS6ZkNH3HHeE/JuSIFcbvjR/GgFCbBNa4K
7rDDrlvIBHTGl7vYszddeOXWnv2uC+yxAejHR8qKh2k0kBU39c1kyjxu6DXxGntKzvTn/U8mVuN+
tYkWz0ynEM3fAhlE+4t0iqPlMFs1luYnCg6aiTTlWV9X58AMUgkM3cSkD2Aw0MFhTJWi27SwKS0e
DoukxLGs4OQrYt0mKBwhb0Aam4PfYrlzmu3I7eI1SQfKRX9q1d/KI16A+dEnvGq5kKxygmdb7pz2
X4C2DoNYdBgo6QLrpXFWnHVFK+sD/n9JxDAm9e+FISQlODEWRNDqjStxJDOyuwG/z9QXFyZksqdZ
sm0fWcoGToGSutXzSYd7CvsQwcsyrg9Cq87gu8aTCxKizVaVnh8qFLO1ffexghN8GBFagUUfh/Sm
CL58qQLQ/qZZk4uvA1kXoUd5h7yps/hNSVzAr7y+z6W8jaoaJ5QvUSlbcRY0k24Xicc8Ut2nPhGm
SrPL8LP2jeHEfAezwArH38UJE3w6XJp+raslKrPGyVmZEDnzEGkARdea98IkWheb2Uo3ukoNwxPD
u6ioXEZLHm2vXFDl4mu4pD74buqQyXQygB02oMYw4Usq1B8TQGnruPxqEQVdZsO40MsRrPrEoLiX
ZlJKvgsrrWyNbmxQvlOoMTe9Cwz9piuwX1KlmgSnaqKVjK2ZN8PDJsD5lnVxCNdTnwC3GSdtO7D2
IXKfnfE+uoQm9ukBBtRZlWy1jfUegCrLXSC3nXy6QSKu+0+9Ak2WPCRrgEcS7YWra/GG62psv/DH
2BBrWRsKd4DxWvenZmQIdCYOAzsUi1073vTEolF2Hpu+kyQtOBuWTn+qIPHLmod1WRdFS+CVhKbx
qJwuja2BY8ukxMBEuX0Pjr6wNLftLs2W213EgBlV8NaeS+tsEtVYl2uR2NdORl/gBbqC3KBQNgWf
WPjc+0HQ6depc95kS4JJqlAcM379GBhMcculuIK1q59g0GJfXAPpxZgpDi5soV/ORDyk1lVyitBs
Uf8oAqlKc/8boLANpi1ltIFdPRDPfvHTbj6aKUVaWew/OfxfjeSstuF8vlKkOQolXJLxYU8eNFeF
ZpeoM5aEg58tpahnOi4qySXQwhx4vtVQxs4IijJIwdfAOjJYaeTNUFQXUneoK3jh61KkebCmnsZh
Q8nKNNZ644VVFDlzJz4WP2yMc/L2MGHIyMuyLIZiWEnKg9fTfsIRu94HEFeLK4ydBWnowMPH6+dY
tHJkULsVeVIjDqkFjQnftwbDILxp3dexMALJ6q7xzoI4TmbEmOaYuz2WUTIDBEWEBa/7aLoVG1iK
X3+pH4YRYyZdZNnVmG8y6Ggvh8ofsoyHM20OlyGJFX5+tmDwHQ9OJR8JAFgJajlrdz0Erxf8M/KM
V+ZTWDSTcFN1DG6I3dokfGdAOQ8dXIhVJhJvXrnnOArodb/1r4WGeyBaZPl11fi85e7AkLndWZga
UbgFeoWquBBuGR1BegKqnPtAtEhjYKWZ+VSoWOH6hemv6CQkNfv94seLmU7qn8gzlXhXO8MYzANi
+TTRzObgIXznnz1AeTjzM7XWlyNNN5Cb2KJ+XrjMKxW7+IwcPPyWbxcncftAEYhhGZpG5BZPQmPG
NSr48Wyuj5sEnFuZSRHXzHXOrxkTQdy1j1UMIxBufBBPzXaYxdz3YXKk8Vzc3yi/bvNmJMgtTUBe
vnYuTZHunVZsE6uGrC1fxeW3likSkdRd9/0eNxm7I1zOS+adbgW2byOeB+jGx6uiV+VbVm63unjq
ynnMDVtvJP9dxGh21iBTH5u0bJtguqL0FtT736ESwI5oc9TfEACZHFfVentC7BAAmayKfLu8XRB3
TsHF3K/riqXBW3GQAigOtbXgHCVWyRiFQBlj1YAjPKoU8mk4pkXds2HZKmTMCJZoJ4rmlaWJqHH4
C40qngaTxnYOzXypxbJs3/oH1p/AivKqvghrMzl1Op/SmrvwMDYaaSx8OJhPmDHmsShGPwqqBM2+
o7e529jRyL6nLivSgnhf53OrvMppw1jjwHMhk54erDSGxTzS51CN6ghbocDADAXKo0Dc0mduamuh
fCzai4wP+4WEYOdDT6QhxJl2a9IqRAhwaOgbQSEvNZUaEjEc7gpU4+ygkh/amkp9LmCldmOSt7FL
QchGLPUNTozCOvOSlqTzPlSuSvK3UgAdHOop8VvZeBRrUOJAbH4+q9YQ9zksGdGrikXRYp5pIBWa
wRhAq3bW3v6riNxSum50l3j08XZ8Cc2xHUtb7CgHuyxY9eYlUvosHa81JJjpjEMOhoPOjSXIXH3p
l+orzTbcvaDIvpvmBntDXD0Iad1pZCV7w43k1sktDyc7fl0UrGhnW0+evLkIzrU49+FuQS/sYZzl
GJ2fWcioCX9blGa7I+wgHfxRtMKFoa0S8bEjcffoddqeZ800necpDkjEL5BXabg2zjLz72cf65Tf
xAa7z20RNb8r4PZxB0QkNIdopFWomRB9L7mtjpjvs3E/Ap1hvESuOFawvViwG+1Op7DJ++rzyKMF
oZTaLywngUJ/4qW7tAAG4jUgv8ioUlSsm4a6nLm7U8ww1MpmKxoY4tHYEdIozbQJN/J+a3YqytKv
vhPtMCUnUGhxnf2Ioi27cXourXxRz0xi9TuqmSoMMcT+dA9HO/RkaMxrikoBHSDsSGlvSc4qPyvn
+Wz/5ozsVDpiDhiLsh3oE/HXjK2AIWz0zoPjT3rD5n8cE1IM82LTHEbzP4qCAdKNzKZp6GK/5NiU
V70JTHt/PRMR7HxhisXYSZSrTdEB5ofeQHwLETTy3NDjNS16UoITmG3wtLfnOpSxJeHJeA4lLjdT
BYR0JWOAjW2LM2oLq9kUmhOZsL7BD/al0J+au04aR3S3eXpt0IZyoc2n56eoro712Bess6HHF/9E
KwjsAr4g+1UETjXlCp/81sUq5quSxx6ESGi1GljeyYJ1ustkTzAf/U3nPc4m6Qf7xD5uRJKg1VB7
1rMq7M8SuBQUWgbGnHjDJ7HAJKiXtxnOkuys9GuDkYZG14I5BAGmGYNfB1C10Is4EvJ/7uPyFgMY
0L41780sSM0ZiJsyZ9/DZbz/r0wplGfJwj/dil5L2GurZK8qYuSnfuZmINPMn87rfcyqyg9s3xsg
Qvwn4w1PSGV9RsEuWyOA6pjoVhepHJlspeou3TRg/rNYnXx2GmG6G6arnu9QNiTl3xXdnfSFw6FI
1q6zzDMPcPv9GP4JxgXNQ3ICJ9tXG2srKqcT2JFENpxBP2Xzd92HSpYCfEsb8CzoFnRFWY132ATt
DMX7qhfkObPgCvOZ32X26tvPH18cnHW5nqAR21b8jAuAOhQ3uezV9nZt96vtNYGOI3c89pmyMirY
OegU31ytx0x/W+9tawqnYiRPiDdoFPxtC7YyIsq8u7oqeE8F8698i+fO+iqP2+ycg5d1LyUQgODZ
dCghdkXF8yu4P6QPLoygZwjfqy3+/LbNVKleHCjBdgcTzCJgj9t8NI4QjrQLBGRXFw4GzVWiuHQP
mRwore2SVa+2Lp7ktl1Etv8NZla7C+gNwiQI0CZP7s3cJULkw3LiuuWJmXcLRSn9peDGasZUfryC
QA+QRG/CztyQprlBIU3Pj12O459ovide+ncMclDRMHOgyKLnz6RH20d8vSL4EmVt+KXhsXRo0FVd
zYVcYis3VvyM5iveRN8vziO9I3DZgTiiLF4N2aNVjJlFnIPAY5V7rL2jV34izLDjhTSSWzB5qhCA
GefKccKY4a9lZR2KV8eJYyhkgL+uelqPHyWYqTfKpzxOHoInVD1OVolcITCnEcOY0Hgur4wNchbF
EGUKwOmN9a+3i4wtlt/7bzcRpS/XtUn5h1i9mEfSRRmfy6K6maJcnB3ObVH4odlPCqk6KtAG7v7A
yL+k5sK7c+yFFez07sNGA4Zi1/8KY0sklGnYo2z5JcH64/aj9/ro68vLufhN92LN7Ngq8mv3qpyw
Fyeu06GPMWBt7DR9DyhHS/3ZW1qbgxvXOKaKuTHdBKNNL9T6IqQxlQQkr36tUgDxMEQgBp4CWcS2
sZlRkHttv2X0IApwkjb08ItWXY/G3gb3kj4tWMpDMzJeeH5x75GK16migHRRECXpAr8vpXNzJYN7
D76cEnlKNA92aT17yPhLjenL06QRiRhE+gtl6ISjqrErXRvNGIS27A7s2jCRi26FUgOlidtLqpG4
q9CJGPjPbVJmSRC7efHVLTecWCAOzlDOV31g48dvKx6s3wkHHVuCHwUex8Bx62ywHCTfxZu9vsAL
9S7MkvaPjc1gCcZswcpFgLQzwmp2hnmuK7s8xLiPTNT6axUwg1sph6mpwo4UsXRPhvHt4zpoqwky
ShqrEAlzPu3kwdc3sumEaUsnQ5Ci5Uw5hamN4Dtqgy1ac8weBCM89wueX1iVH5zYx0QQFr7mF5mP
eygyBTrQyBvYjIWtRmz7/W8oj+/ETpNpCm11kNmMurXFZaU6/wCZT10qeXZ1yOGF6xFZbjarn19e
aOQXPAr3u9lWhkMneXHCsgRs8ivMdmTbcQwGo1oPRfNLxJAVq1MQnvxiVNXB8bgx9kBWh0VW8voS
knVnoPzN82SZUx5UJ5Hv4Fle2vrS/RhlVqh2YkSJnZ1CurzgP85TSQfy2mp91g7XvgAItoE921De
IueshYLfyFfr0F5+faw71g9oE7xSG7vHx6LAr3LPQ7DlSuevbPoHk27NiedkHyd442udJ/fArPqW
NtjetcVsMfWPQ00+KcUdDh2in60HyQ60hIOyZHIud0q1h1yRoe0ktpUPMSENIWZtdQ1J7/DuGOBT
RLn83KveDNBYg2NRm/weh7CnVQkBKsluYYX2TJz4pp6yXLd7Oo9jlEB81pHAn0cDNeCrHj2q6xuC
HT2+aHno3JdV1WvXkCdLzNd0eQ5PVD3Gs9X85aDGdzoJU7RKuI2GhOA7gWNUfrWUBmQh04hSVgdR
1V5BWIoDx3oDGr+8gp5w+VuBIoDGaLL3wkXtnVasuj4C9WI6cyTsfLqRmI47EQxgPx+A+KntFlIa
wLiHBXWDPSbHvU/5sKUvB+6CEBFpnoauRFaGOCCUFBnuyPD4xS0H9T89lLb8TIxXa0GgIJMZESST
LsoPnoUjbNGznDR69iQuKfy55HOdn3qxmOCIIMDT7pq/Jl3P8foVpVCYBMnan4ksCbHcRAtYu3RH
91ktSN43+x9yB5FgpvdxAa2sbZ8u0+667Vq1SZteNb0Yvs5iAkQ32/KI6edtssMrUfe2dsBJXjzB
vb4j/bvNswyzLChWKGZuKinLwmRnV8o/DyZKNoT1mRD+3aJfeWvHM89yHc7VkI731UyHnxXO/RCr
R63RAYVDyCAKyuOTGjIZfjMEyUu4uAZyzynO5QzB4tw3zy8lVllelFNAYswwElwxHSYvuJqftMjw
bVHAfD0BkwsxmGQU5Ijid2mMfTGgUhqIlGLJYeafF3MIyjvhOwukYoXhm5+ZFpja68Ke7NE+bDdt
sDD9H1ue+bw3YxJz2fC8fbRf4toH0MR8JSAQGtgWcoOAYD1dr+TnUBzlIxBkNBHd4W1vyXZPMoqi
Lg6YgZiJosMzKEcUo0IORBCtGdEv0ZzMfbqV1Whe3NOX54JLteQjcUCLeF/15uY+VrCpsec4Hv2G
b65alNYF/qAENcSwQXu9hs4345CxqA3JbYrW7TE8/E5Lkg2MML7wMMMuOnqdbLYOEa/SyeTomQ34
SkBQWI8uLnF/iZ05PcgljmRP9mxIdbHz2BL0z5iUAo/yAm/Gn0TiYMaRbbUvrWJQNgR0z22RzZUy
UEvkWu/0X3q0HrLRndkn8emLBCvvJ9FjpGabP8WcmU+EyJRyw0ne1L6OqergTnr3+hSkZ7gsL+kS
rmoa3wTXczhPg3qoj00w+1LosXWpD3FKxHE1QZ2B1qYyfJpS1GrdjFG9Ye5/Ualnh2Q7uR8Sa66W
TpxQSJbmvkjNed5oufyU8+ekRdvbs+n/IqLxzdXVzCJ097mxoRLUoKdpncrCNFdoJrXpXjjb8hZz
hlhLmefZy4uxPyVuiHBy9+PHRuimTfGDjbK7P13Dsdx2AsMjM84fwxqbtoc82+UId/OZKISZuyLT
uEg6EkC92/Ln9FrciTwE9n1Kh4DgH9vlBLE2XSykK9RIJhDLjOAi36OvbbO+F9HRwvic5i1de3FA
E9pfZZb1eNVDH7gJwxQcIZrDiU3bpJDExprZaKW6S6QmTIiA85NiYqIX/2A/t+yxxI0tRfGjrFrQ
V4x4G0PwANu8aBJbWAN2MUKNhe9aDTQcptUOKEVD608zJYl09dvt/8i+3w1eG0UnWJr2sfiihk+a
FciyCYaCSJqWrSo8as30mx98CHx2nMvBNCEDcap4eH0/U7zq3tgQObIWM/i+HHnXnJdkZyCbEZbH
PCUmV+MDPaU4JgbiztxfSIkAViP+JmbBRkjiBUo3/CEzkQL7zrYauMl7SiL2mMCagvI7LCF0C99c
l9Kw/fHtBvfkEt1plVAw+p16WdKZqXaB1uatwVfDcw4Cyk/0XpDhFxL1cJXSQLdiEJGqr8ATVxMW
8RW10C07EYaalcAQleDAzPTnH/upZlFvl/qHsZxs2fpdCOo7hcXj6dAg81GFyx5nnMVsds3SXsrj
/Kab9P7Lj7+lDfYh6UKV4b+9FuvzK47FrmpLcCKkhZ+hcKDHkXAiooNejMByaGil8k6uStOmZh/W
v8BdCbEjTf2U/4UGrvyn0j00WNHuB6TWBU5m4J/0d8Nr7zHfD2zWFYpOkY/9HdADATXmGGV3TO/1
D4EuuduJShok8WdtC0N17m/NPM0LMMRMYoAzM90k8wqX84Tnakc/QqO8PsmxuF7Fh/UQJbNB8FmM
hS1ZXjIruF4GQhTogl+Glh0POzMqkbcu8hSpHApbkkcYC0TDLZuOEuhjMm7N7225CTeP+3u1I4+D
YlZL5SGZ10IrbHTbdxHkNyqGitFBppUf0vEG+/o2wWHw+ILe6rpqg6WLzih8koiNqqbu9CRHVe/W
xP6ldY3mw7hf1xbJgBvJ9yQaR7Fcgawrr/H4hq+ftQofEJS7bn2ydcVXj/WJcYBSv21KPx1cBzYV
pvfELzqXycZr5aEqpwBwfo1ObMpf4/arpAq7kd7zcOovAZC7eM/11X3zNiS98uG6OHAF6vH/PKjh
35ZhRzf2xMlqyE4D9vTPMkUQqZ9/kO6exOSOAgjiWmYdxyRhDOWng5mESy4OemJXl1gVlqmcf/eD
OWbB8i3e8sPD2QKyitQ3UM5ixoA8UVMy/TvFWBMsoG+FEB6DKlHavnwcz/loRS0TxzYhV9gU1jGm
pXl8ambFip7VAWihBE4YXT1tP0MWK5DIDMqxryJ3rF52pQf9QNgI2jLBXsivJPMZUiTRlbCFYne6
kpZRZhViOZ52JiiFEM0G42SxxSHBe0ha63ugfKAw+za2iIsYvAPa6dazHHMGe8wdw+In4obLZGRo
4ZFOOMizz6U8TW7frRyVd+l1NyF56x9lXUWbjlkGa6+bllaSFb43WPX9c3bZFDhOWDE4Rg4A0But
ToFqkuz1xIRvF7jftcdQIxWIEfMpBMo6Huzih4KHvGGaxM2MMTBfOXIeo0FS6kpqw5Swb+tJB+s2
7cNwD95lqOS3thPWosrcE1xFwjljK3YDKiouoy3ojdMZjxQbFrrx78N0vqXNPTUo2nnwSt0ig+2y
yFIScCH6Zo0veA3Wkiw+n5BN1SOTbDzcEQFGajCr0UqMFMYusO0K8WxqbYK/v4rpBCeC/SasghWs
5L6fy7M7V+lUAOJPgOJDvguVmBUCyRPLIUbD2h7PoyLm3Be2fV8xq/hf3pfMb45z4Su5ktNlxmUI
ZXeF1UfeHdPhgjDdQgjFY7PDIdgmCSX0/t5eWc4PO6AztannN/QI9ManxE+ljRPOdigM9MAMsj3B
0E/nDmys+iYYUf2tQKm8vk0Tuym5mkatY6vhzCqcO3XplKE/JnJYgK9lAS1/yn3HPjPXGLP2olxL
3JOOHQNnIzVKELb/O6UTYYnSZkxr4c3ojAYFWPVlFg2lQMj3t7JTnGZhpjPXsevw2GgNtOpszFSy
ZXjUCUYmveaCByRy5tXD1GBmw6C295kyQqSim5UpgE14CB3KYQ9h1dDxK1jm/OesG+L/rSa5P/ZC
y8tXq3imIXlrxWDVI5utw96p6sTLifRntoFKFhed0iuvDblmoC1/Zy4s2KkFK8sf2/Q+tIibjr+y
WwChEBBLX0ZAeIBweUqVoGXB/XGAyL1f7A6vZZjUQWafGRv88HR63wlVMwGPxegOBU7Yr1eO0rNs
QQ3PTIzLocBgNlQ4d4J9ZbSP84yx8LArGQ+a77qMkHef/IlVWfJ4zYMA/0x/iPL7uZi42MGllEkQ
X+RiNo0mZ0w9ZDBwNHLkIWc1GchXF+/nyX5El9jGXJsrtvwlMh/T/B7mYmQWqH9hl6F8OWdA+QpG
uT/xdiP323LyqLEjsrnvalKiJKYNu+oIeeaMK1xSDWc33tb1owvQRZ+cB6vOzQMnlwT58ZlTNvnW
ITqtVAFP9BJ5bgO5hVWyZh1qzgEVd3VFFYLcHA5pPzY+c+XhRTt3Yt2KQM3JuWYg7JqsHuxa79E5
ZC0QhibQPnVPnRI4SfiIdFiDJ02lYKAxATr/qDdh/85uCmOVruZNu1NYLuFz3jj1sym9Jm4TkOY2
zfNbqwznou+qyfJ07EiI43qVx0WL7xb8pzJDPIPh/7eHZS5sjP3Xi/bBTYRuDW8OBwbqxwjA3SQd
TGINsl8iI+46jj2no79EtUtxWFV63rtcK/MBZh8Vftp7Tu17xQZb1OAhHgwG+8PXFd9qmuQPxVpq
x72fmqb8RyLC8/tP7FCBAFXJfrsMS+5fmYGRk+FIXRflQ/lC5SX3Dup5SSyji2L9csDrojJgS0wR
HEn9y9fskxulg2P083UfXxpxUnnpZscnw0gwTu2s6Wsv8vUZJQmm/6b8LLvBnHh9N5gC7MZ4hQnX
1NoXzGEYnvBCyghC7oleb1hHD6lfohpYt7pj2qVS/BVvcoMr5DrjwVeKP/P8+59BAtnCxrjksFB+
+GJaHzIOeO/oKBpNwQDMukIYEymtdAtwnS479ylG+aUF/r0Kg5rfLLIHjEbapQOE00sTmlWG/EOa
vZysKL86VDkBrtk7zi1TQP7bZ0d79Wh6Qvf7GoEa53h+AjtMgikpWMi3lqPfBzbhDDyfgrIq5iic
eeU46SroorzpefOSmmtf5Tgdyz4RscpOiVFQEoCxK2DSftSAyhIm8sQoRJaPc1+QG0xV/FwXI8su
eev0TT8SPV/GYAZNOYrrCaFLTw6abaHi205+dnBkjLai/2DAXdJ0wdeXzzID8X88zrr/mwlrzmd0
SxntnGxjI4rwYS0rQ9PpP8LL9gGW0rCNTGZ2FWKpUACoRCSHY+8go4lmgxa7LdMcSD3IfyYRpOJG
7BrHwobqlaYP4d4vs40uuS+qpifpQwH0BnxY34p6Nszlb+1x/UO3gbKSKK/ciPV8lTYPvdH2Zf92
LdOYdLu2BjVklEBtSBZKKHqZvxUDcBSQdEh1U4bZBLNrjuue1wnhjmYkm1l+83/FYSB/j8yU40jC
dX2Kd3p1ltkYECf0XVsM4v+W9ITVxw7So9ws2pG9G3FYdRcNE36c7I92u5sHa+7b2dvmF8hTaDkA
t8vc16uAY+5t7jI9+knP3LM1JoJP592/zHcub8PX1Ho2dDgn8xrHPRrSySrpHfPl0uN6IGqKf4X8
wvzztYf7s6tFNZsZErfaj8dHO8fErwHo/qha0fGOlxnAyYEuWe+F6d1Lq0cW2E9mTpkaen2vlbrE
tHk16FhZXP0ojlggGghGpGQYJi2f/z9eBrcyI+0cPLez2wmI6LQ77YedogdQzxR2cWRpcdikjnra
yr+Q8vpRjlsR4NILFtW7Xjli2XWbDHMZD7iUUKcVIRWThR659OdeQUbF+/lwo4vYfqIjcVwgvZSk
vO5fsPRUffDw5tGzHyKJ6w4bYmHjpQBsQCPB9OPZTLvqoNJj04xvGCUgXUXGPLd02MfU8gWpefRp
Wrk7P11e3U3K1ArUJPynCQiv4tX1XzN7YqGHo5vEVfMqsdcEjSPaCtNhO4i2fk8v7UUbDmM+WtOU
1XAlYVOeK2riauQRmSUh4odD37xnllfbSmvigz6S6YzJy2Ktj1bL+iiFntxyOdMq837D8Nsfg9Ki
Xsj0zASp6V8A+rqTLgYgcLbdv/gfdoJDnOMuZ3EyukTFkoAv2gVKhDKORYAwVGB5W8HXo4SLn9UC
+U9RM7UMykwURKQzvU9kOD4NXnoLaq3YjvrvlBa7SpOuPS9byxUywfRuq/20n4J/eSbKlWLI0hXN
UsuAktUb3R02ILsdRleqEQK2IpvNKy7/Tmyg+/K2sLn30AkPi5yX7EROGGR+TtFGfTenlfj5E8Ek
4RRF7V6Ch5bl4zBhZjv7KBbfko+N/bPkwHg0WEMTVZkdJUmDmb/cQqEzvUmysAj2NCdSFawZV4Uc
RdxOt5EPW2TgKtjMzHGrIc86y+wr5XgABX2zXTgjbLPqqAKKC52QKmu8UHaL44vjcF9Epj5zH5PN
7HvK/Cou2cHxXVdBcRsQ9GLK44gYXn03xv2JPdNpWqb4KsU8+Snlj3ppAXG5fag8I8tY9ZdGf1jZ
JysDwB+/wGJ1wmQUYi8bYcHdktazDWNOxKAcDj80RCJjE2jw/MHhg9V20VcvVwEWPRC4y97q1KBI
ZhZgbOp2MMenRO+6hoySPcMwWdJfjCk9aCR4m6eAbTVQT9kEoJZfGMoIDGUGa45pA+MNmWB9Oxt7
UwwH/chP7omoON/AVH+to5V/m392JtPX4AU62EFpyB3jb+PM+ih/gYgblpf779CCVEpowIElvhia
00rNz739wzFKqOBDAXdHUoyM6iG8/A5x1x2i781CQw8z3W8UtV0NW6AXvYbTeMSj4AmNyfJxisMh
O/s+kYlAuikowGQx3mCKu92wL6L62LXWJWmRWVLX+VDmwYhWCS3d2o+o9qgdzqFLIt8DtUarPNJs
qzSz6VA1J+Q3u+yMNsdWdrd405PYnCsoXMvbL6d02sdxhYJk4MuYGgsgoAb4qR9BBixHvSxuv1Zx
8RGx8c0tWx/1j1qh4IowtjN1RxHq/Q/tUjmv/tXaCebusz/bN64Blbjo5XHXYpZmYk9ZatVyKx/J
f+tXZUXEbmEY8YzX9wHahIs9Rn0U4oN1/nnnSKUiJsmm2a8v7GIVr844DtcP1tNAg3xZrCpr4IHq
VMhtrivpFOf0jt2+XW6X7YDua4C5pGX4Ckupg9d/fa8wLWWwEYberFN6M2fPgTsicamIKIyojdBJ
dNii4gEeXBpguSLhIBpy95LJQzoRAokmaIaT3gxpc1OUMWTknaQ8zcAvlPr41cJ9N7+87EeBPJCY
ePWANOo7wruGyak2w2DBPte74/kFTRP+5QqYl8pqsojxG7jjFZv3bRWPy/LKWAJXw+YP4G6ydNLY
nWTYhVMi6zuexzHS68HVH0XvfbUHN+LaB2Fid81bHfkcloTSbb8OvpPYMAi0ppsedd5wG92kMWkd
lnvP19MlP8eoasG+pUCWGAiK0RupI9WYyLdmJ9oMI+cRh7DGI33O4pJg3/bQt14YPViVoHtE/h1i
iMly4X8oNF7qXCRp0dMf7KHyOUUjGGapCewun0T3wGomWP4peDEM4olt+vvjrLsgJQu1XRJUa3xi
HnJdMvDvos3V8/EoGPz8Smke20bzHZSlKQ/Js4t0CqnIcAEnhvzlAL+I1mr96DPJFHDppLgsZDlz
Zt7xPje+vzl4Bzh9BtKnneO1toOMmo7g2LEPEwz6KRdwMwvv9nO1a/R6IIh4L/bUlkHYuODXPm/x
qKIXYulcCZUA+1WnsGiqixATq0mxn82V0FmhJWNyJb9L8BskRuwmblk8qsr5yrfrvyPC1puUf0i5
FAsyRoZKVBsCqi+Inpw1/KguOEMdMBLQK8Of0ACLYTcBSz0iIS+KcxkNxdAh6dIqccpnAkCLGjaO
62ofLrNRIZe0cQ72hQoESw34RwqlfyYxS3IwMmNUcM6LNqQX7nBDyVlCQigxgjb8Qm1NdBens+eF
ZrISivvuStodNZquyNl2CFXdwHmRa+mSVQ5oE6El510YI6rxir6XQQ0y6W5Z9eNuypDFO0RcRima
8h3MQBOu3H0QIlBhJLDl/1yxp/xC7lh690eo0NGU/MyoosEmpM8aQrdRhYJEu3ULNVtkL8Ex9Lel
i5NTX1yUI5xG1DkIdToqWNbnBD8+ZE79su9bt6LoKAzTOt5NEQGhfHLZot+7s8MudpcLMcKepzBo
qjaO6fDnsF0Nk2ciN7SenQNC8i5rv6SX0Iq5N/Awzt2dt4+Grt0VbuvlD+2HkYmI67u9+HVsan6Y
USNLprD5ZgfHdZGn+nXNc5jc1yQS1EGnbQQUP3GIYL8aMRppu+sdWV+59j3jcmozb3s6jtBfFZf/
juvAfdk4aNA/2nOGCNuU70/UOxZYSZwOIDiCbKD+x1eDbdSBR9Gt/BwI8o8js9Q6wof4KTfuZ9Qj
hSo8HWqfFjmGZfRN4qRxdxoxzi/W1t0Q8De3q9TlGg8KunzX6bXauRSUcxNKqXs6n1jNh3XYMw0M
U82yk5Oy3yLwDns9T3b1U45n0lgnDOGIr24mcmai5xUmCW+VnX5lD106Xop2ysaKFDGdbkXg3lrO
y9lD79S/DYthxxWAAGRpIosZLvG9zjzflIqQ+S3UUjt2eJ6p5d7uc7UY6lUzW6U4DDW9OzLWYo/7
YeguoIaHsdEXWbISni1KyhaMcWUpuZUd8VOuxwU1DqdU2WKUO/2BwKoWCTNk87Sh9Qd6bblJmpke
9hJYuo+qblejL1wZBAJZWETNiyR95CycWe5IfbZE3MHhkzdUgPFRrd1DqcTiMoGoiY3jY75AKj/E
Z4T0/djyJCtiTg49rp/6BH+wNe53RhFSM9PjZ2Y3qlfU0ti60gt++VDc8Wcn2S3lnNFvL0QeNEzY
4HeA22IK6xj3yGksxva/BEAszIC9+ebLunuyKTZN4uvKCV648HRXMl7/xYpQeOSAteKz1ro75JEe
ekfmGKPfA5DnOsuJngwNE3wFLh7dDqb6aikpd5wiANB9t3OVsunZz1F3VQANpWECzlkBLW5Vrqlo
Klnmj21KniAOf/wx3bp5cfcia3tUKV8DRzIxF9JGwAtO3AzRsmYh0lXh1rnUccdmyhHkMi//560o
w5A2W4FBz034mglHQeSr5XaZN0ZOh+/ZVOwt5ZOFZqPHvQHyAo1m9a+WilRjDyzWUQcMoXxbaMD1
l2dBKLuIbNibAAjYsc42B0p9iEqjF6cDG8bqHCL5LgiGKJOy9sr2IYh/9Wz9x6ZKH5I+ud1Vhoqt
UOGE05NnMywXNWoJMh1qgmB+AVjvW3CTcG/KotxQ2D5CyE4qjd5aNmnYYvLbU4IMUPK5TkiQkdGH
5UojDKftXeuVhfTW34zvrHdoZAba0cozfH0svGhHAhhJtBYRuEcvjGqeRagcZzyaZGagbX0zhqPD
DgivWQQvhzWXa2g5VBeH1hidO8lDCfoNIF/3e9MVFt/ALOuAip15ra1Azi3MLO3pCLGdaUsi/tcM
bKOmIkkL4ByrpXH856aqpeywRCgmzoxkwBtpdQZ/xy7t+drob4mY6vxQcG+uzpMZRghOfoC31IdY
g8cfLhT+mo8tvpKJxL4PihJAQDJsqy7q8TpIicJBI7EaoqSV+zGh3re0eWeXjM3Rsluu7xqQgCMf
ZiHW5yWUm1VMrKgev1F7CtuOXnp1SIeJcBGTmErzS6mZnm58shPznCkTIXipGGTEZexppVdk0Cua
Xw0G6AxexGCaXBctk/QqX4zxsC7Y1N4KIU6U7b9tr371ulZr7dgq8KBe5rwRcUda8UnRqb+QYcE5
luHxJKFXJx+AOdc/rEAxlyUBGlkjQ61vf+ciLPToqUr9tuZXrjNmpuWVCz3LpcXSFpt6tsf51uY8
WEkCKVeQHx3EAwo8eDA6DLITnhA74NqgbNED/zNGXhplbZoKa2XI57YtLs2RySStvOjdGGwSwQFP
4P164Km0JgxlgkZ0WcnjMorGPijX7pS0o6vWvLuIPIlozLqTgHsM+xklu5Jg1jnBZxii86sRcHu0
vPUGwPTCLqt/bHhD3IPH548Kf89czthO43gFkh3OyZwNQpPwW37QiyC7szhx48bEV2zQsttqgIT1
ylA1RRulQZU6dNQBZLjoVYGZAt9rhP/yHS5fYIeHjmEC9bDN6U9kyXVXkpf/77iVYJcBMzYuhrm5
cwIF+WQbisP8kipcVVKWUC0szGbrdiwwojLMnkb/02mFeafZ/QoAMh4POwMF5e1bHXcWSV8DAK1N
wcBSFGQSGJJjpPtbSrFrAuhbw2DDdP4ljheltGwlV+asr9Ia4lhU1BmBftd1GZ+x+hi3hYPJnpkb
o2ax2n875YMkWeP2w4nVFU1C8VYyRqzDwcpHUxvgI0/Uz0hcKSDb1X1056C4LYhWTHrj4MrzKygw
Khd25jwpYnv0LcJMohK3tx+xTY4VSTf2xiZIo+OVGwGGlUjnZl4DhPoVHP5UvVO9UVaYkoELBWsF
R9ygRMTwtYPvi/wgF5fm8Rb04b9aHz55bBB0jMb2PFmNxYY1b6o4FKpv0M7/dBPpCXRVl8UDUXg4
qHUU/+RGq4KhcKnW8t00Exp5E/2o9lyXCq97DBc9wC5u1lAEgdxpJ2CPIMqNzU+Lm/kQ7vn/X6fo
7NMel0JCxhBUDpdcsznUnm5sbI9oywjwILnx5l4nXk4i5/qd2Nayn6OiQVnvMvziQXVzad2Ydi54
Wxu7Db/d7Q7e37aeBVbXHjjK/3lzHHGDdYiM0PMljYhd/Fub0tuQ6q61Ifm8ohdFbSddxjk+ZYv/
rFXVpJCaj5kXVM7FAPSoud67M4C3xEJKuM3cK1u1tD0H3IEcvf9BQOcgZiTAg6JR8CRs6kPffNom
0XzwbtW3CQHKlvIEI9GB/H4FRoIJ7F/TDeIepWeFs87BCwYZlIdvvxVnwseTv0z+EA7/jOYe127w
xKLNNQziIzyUTmrKc06i/LUopJgSzBT8UzAhk2kN3gK9x32RRDKa2oWHtAm4+Qjvj1+6xwNmGs1G
I2v+uvX9DCvxAqQQXAXEJId+gUGkG5Z9sZ7RFbuXquOJcM/tja/tpnB5vwEsXQnicwc2WAEk+5ee
W75ZhN5eGzcZLesICJhTd0MTh3a1jQuR6QnA6n35+gtErNZpS4hKPgXNpUK/pEBUH4mYQ/ZgBCmT
GzTjgt91GP/h8b1aPBRlNQ2gio8SW9wSlTmsg6iSDguoPA8SwB39W5kzdPDEsLlkSnyxuTqS5PA2
mzoVT9q7nS93UMR4WH7kspJ9YoaINOAnIHTYZLMD54sOUNOUVF3iNoZhJAXrVdWCIrFJCxTcJmAc
D1gjourbyTFzNQxYQzVxlq9u5uhRzJhPNgOjL7Ilvlw7A8tYsGFlb5rf0vBdowE51YLxFAtxVVxc
H6h4kqx68ShoJ737QQpeNPWaNZBBFLU53MTqd509lUkm4CegtPPr6/5uUMRaC8XOAXCm5Ah3RGFh
8darFJPdrUoS38zBzhNg75IR9qTfLshNQkRTF9jdnEHDCT8Z9vVXo38Ok+CbH/YzEzvfZf5pzIl2
zRocGfz4ZBvBFhQyI90DNtcdlJ4Z5+PpEZihgknB0yrriDexDvelxCKeZRiM+V7BtD9o3cKs3Bdw
DR68kDmOG+KD5NZAokVkHsof2BEJw+TbS+ypWpjqTYTTA1LUU2UKtVR3qlXO/QK7ftiV4lveSd8j
W6/S6BgH86jgfZjwwOjg+cFedmQbTVkvzuDrzXEtN6sKYIPfrp9sFEmamitea1VmFuVM8PYm4nWm
fBXnDhhYLv74CJoRhv8m1WZiHkjS+ccDqQ57bxWNCPAgKf1qirUaM6xhxKN9L3/OJbIxPW3dbLqb
wMKY7eRzJD1avkZXeRRoijZqnS1FtxGUD/kFvmLEgSXwH8+WM72QNgYSff3gY3qhU62pY3mkLXNI
MtCDi9lyWVUrpysuNKlJmPpZRfgjuzfHp6vOweccO8UOz03d3aVIgTw4/JNSmdkYZwlT3Yx6lGhn
3ietQsp3P/g56QqIB9qjkWpaSzqFgMp5PvAO08G+V7LjNYhM6FEeuQKl4SYbYGNJoMAOUzBy+vxH
74ZENO+mOqjrsj+59a5LpUHc+7vWMxXm2awPKPDqi579vdd/Rc8pTu7TLdDnXr6ndyJETZwayj8N
JXYFdwAvHAUPEeTsijNTD75PTRgD3hbXbgJhFsNuCSvftzeG7KL/QzGTrTHLvf6qhiaS6Fyhzsw4
iETVqgZGARSSkF56aEY2Ro8sQ0EeDRW3WOUzxSfvSp2g9EanpQ3scEdvZb0ijcA05no2mcLO+KTW
9A/yVrhR/iYOJvtBCzCBhGm/L71rGDiUztLoaq8xhldNXrgPglbYcYUzHTde8s0LZz4U1KTfmRs4
sxCVCUQjSVIReog0Jgk1Q++XXu+n3Bhzw/x9yvo0RGscIDvQtuIVULCuGrWNCVrg7JKG2zyV2upJ
MdUDW8udCinu+wbbtO3hDcKpTKUXsJvI0jlDB0erm1AaL2CFBm3T2Q3aLVR0sN4sHc29RgyhhKn8
I20kTtXdPRKxWOSzUv+rU2v/pZFUAhOOmjIIo26V0cPDJfwTEwhKzMoXGmQGd5/fga1TNpIVNSI2
32fLBzXDT07z5ky9A1Y24UUhUjxisTewjMcpGX3viGC33jy5RIvSPPGDO+13dUsvFKNzKfMKSbyZ
bq7UsS7OHZCe2ht6fmr2k1C1n4nMia98OTGDF2vyDshpWCEq4x7iXlMCEjhwVqttmQNtBWjZoIqk
Sdjl59St9eOpluuehmSoykElY8u0fehuYDWVh442fPKu9vmqbLyCeQX19OgMOVuZdO963JnnyZj7
/RstDs6x/vCz9BIYqhytXwDNzr97YHyM9obqlf9O5F4fQoDMCDP1TZ1deJmGOVMy+D5fheXpRoFO
IqqA3d2Cb9HUh2CFkzJqHah7Zvnmf0LtfL6c9fdMb0b+0wB+GvXeYp9H2OdBa1KPtblwUtcZvv+D
zWY+bn+aXgY/mAO3y0ZNF8GWAQMhzaxE+DVGhd7Y25GM0gIJEjE6noY3YA2RYb7U9A6EJhlthnMB
gZVi8Eoju6V3eENPEMC9ZGBcFDtedxc+Jvxtc3w1LkG5gr75v7M4FGNppfUzi3xCyXRUWWBTzxjo
WO5Rb/YbuyLxHewRlg3nDEo26onl2MzW0Jg2gGEGJwoRtPK/fRoudkAhvx6t9EBSXyQMwhbWZObV
9zhfe66SASuTDfayJY+16VepBFC3haYVE7miuhSfH5RaSWfu3EAdg0tg3HbuEeEwvQsBB11cf4v5
9CLTTZG9CfimvdVZjNtdG5KLI8L6wOzFjyymsKBzBraVaGT47NNIXNnS8Xg+C2kguDK++5MZKMcn
iqWRPDR8WRPMQkzYuffDQb9wJ9cHLHe/prxG4uCwoygEL/SUvKMCI8V3hQ/pyE5O7CrKSk0mki8v
U22dBALMQXIIvVyNXxBkoDT2elRnJytLvmZKKsgZKJC9N43TFEkHlrlutXI+xdIobVt0bljmEZh9
DkkSlfPsSLqi6e30FvZjmelRvSL7qaRrWplUzGb83csNg4fcBYO/yp+nJnhA4R3IoL9P3uisfAqT
EEBaJQrHpuIV79cQ6rSIjaiinilMiabP8nj155H9ZHSjVtf6kjv9Ooz4LhKU0bIOTUIDIpFNK77k
SDPbUKquLkG41KCz5dUwBs+sZGbAXiyCVJ9tnzaRuwHxUims8Qj7ZfD9ZnOSdbF5/0qmW5zvn6LP
6PYDGojraepq0cn3N0/TFVjx8dtsQiDkriRJKz6r9CsN/ZJg4XctNDOLIVmgzqGOyELNmkGG9QwT
TBpTw6xQzjeL1/W34MnuvkisaMOYtQu/IAKKgU1cG9p1WMzoDmylegBGaI3LHKhwgN9pY7PVR53B
4wbHXTZYmBIW2EFzScFdOg88GcLqV3jZss9KFI5TMNa1rr4OW0K7j9VMUuvhhfLXQ8HrjeRc6VeQ
Ei5OGsiO64Onkdx2qF5V0OPz1zr4R1PKpgbA+FSNwmsXOLx8af9dyRvsuMBAAAxe6iqJVYbnYq0x
ub0aR5eDSn0pcTxNkyRxtjq+J5z31amg6J4+QI+nMYtJjUwEzukTDdnlKRyNL+yNQVNsj0p/H72l
i2JWKFUf8OCq+eZJQxiyg/uBKSI1gWbnsz8IsYLrGmzcZDQ8jbDWl8/Vmb+Oxf7XIFJN3Ox/EqLb
J9h6VmbiWEFqSA1o8e80XiyoqYWTT2VDpXEbkzdv1Uu5txAjds2PZoUVDm7Jf5deb/rPS00zySN3
g9GZrR0ATvZzEJ+f49n78k4ANO+BP5h7jeTrYZhg1CIGWZuZe63Gs3BcQAh+KXshZVt4Zgfq6nlg
x6XhBbQmy5u2KyLSinXYqCtkqEpoHHc+EGSk5ZrdPeF2QQbtcXMjNEgV5D2X+GaB7LqDlK5DIARJ
V/yg4LmQKFhHzT5AjusXpUS/Y3099NPsQSJ1sThBWtC1K+2U2Hj0S2ur6TamoiUQcL2Pw+BMaHT2
Jd78FqlKI/ipXSeNbrApztmWNL4+sKAiAO+y1vcwIvmMo9+dwdkCUsUGEKcqXnWsuL1sfOiNA5Ri
GJehdGTF/c1Gai6T3AEm3cpx8Px1mhTksDOpPPigL/D9QTTcjJndnDd3RKdGyGTpufDH4uk0B5kN
g3pj8h6RyNyY0M1EzRSXDZ3U9fL8NE844yPbrIZhNNJsPH43sQo14OfiqEd08Ggq0ATRT2k8abFW
2p/a7+j3e6QhUeMq0AqYv1w5vKC6x70jgMnPVW4xBCXNFf/AGCOPT5Pe5sTczkB1uwEDOZsjJZi9
lNBhoEv89kfaC00ig7a0f01KdChuLk+ra2X52VedfCByLeYWrf7eULAgerG4H/z0EToN9LzqFKQE
RqvJkMznA6BRdg1x+C+QMDT7xUvXiIEbOv/+KqTSNOddhyTZjah96w0PAjYfyeupJKaCKQVGbMSl
z5IZmtSnDx/2FoKw0tQyg/P6fekObqlYI0AIGawcQg4vb2PIb8URDDvsg0GBtZ4ltjfrDtzNfmSs
dl4hFq5JQQbKHFFjA66U+IrkAGo1nKUiY4AQ8MGnEKF/jR8N8RKhG7IUVm7Ar6sYDuvggAiP+YIo
cpMXIQnuEx5496xpomIz6MFcorHDb+ytBNYvo2IMzjdyihp5WPnyqbrdScTnidFKVB/Nmi1RVi3V
6DJVVLu6y+EtUhXuK1RUS419/XA1qfu1sN4oqsgH3fCnv8syCJmNeE6aAAGgOrO5mYTqLuOIjeUH
AtoA3pO9ksecZ2brGtznMq6neS7Sg/HOGvrSYDOVzFP2ZZ5+lblx/U6Xssz9QeGQJHe+sbNNRZYn
fpIe1afhC2iOzNx128fgNAnmRvFpFFk7xRLrUsCuaQNKsqwP2m/nquK0OIJ6yzWyX8A8JJUTcyis
pTMsax4JmYyEzzguoGjxaWdkMxacqRpnc7N/Ym+HZ1jqiN/HKa3KHka/6iCLW8bWHp+ibW2z9Sxa
ikHLRxicP3tPmq3KXNitUlKP8s4Z2HyzbhfeXklrGUs4yJeWGrWaGP+W8UyN4AhtWCipv0mhMhzx
jI+RWOonZbk37hmGBzFEgpqY7xs9EH9BoZYtxfIyeeOuj8jAV9O/dajIPH7G+lAfUX0saynpkzC2
EGg887B188zV4+qeSOoTteAHA+tJ90o0mj609ebZ4uK0q00nJe4XnrAbIi6lFMoEI0E5ZQxaA4W0
ZysEW7ANShmVe2he6J6e7kLEwOh10xgjnqdOsNOQfT07m90LQZQ3A5kfmftQ/8NsRrQFjYND+n/n
JVoGOaMEJBWjBVk5RK4M00rStYxaCdZW7Y27YlPIN0LP7nx9EIq7lDSUbnyBryZQMWORFfL6+sNl
ACKW6WGF8KxWwLBUMKb0S+1Q0L+i4tJNfF16DRyhmmv/6N82gZhgdRi5K7qZlcJdtg79q9WMGSGJ
wyzS3iTuA9sW510C6ZvjLYDaWatFIDRgx1XIJDZWGeh4B/cjhwX04yYyEPcNs92Ikv1T3dgDBoSR
8AwqzpqszDeifjv6Vmls8Y+oax1HDTyYtSrSCdAeQ3JsRhx3/iqeHNJOhsZP7xfvhwz+x04BqZgs
N7WwyIi6B6GcjoL6/K20uTsZcwvLNuBb0QiVFpkhP0XNkvvtFDn8mrNDTqG0T0Qz9oErEXukN8e+
RrF8yX7nMpKzEOfxnbZlz19q1wOosu1q4lOO7oDD5yhWDqwNkLLYLFI1N966B9Fs0/oNNhtoY8YL
cW/+vM9v6t3fW0LHCCIlU3NxLOeRNWtQoN8yBAls2NqadJqQTPecV0wZwTlz6pr1pNJLwu7c7hRj
UJ5lGYlMEByNs+uVqRs16T5BqUtAZq4P9A+gAt63FdDeJEU4zwaIiQ6hoNeZx/Y5oS25zBo0VQ2p
iYNhwyPqMLVmkKevQMYBOTsJgw4s3yHOjpvdLc6DJjnkAkWGNmYn7fW22zQn/pmq0qnrxGAGwptt
eAiPyrWRjP80YTgr1MpWdAgt/WyRpgQzCPj+15kLXlyI1znS1C/BcVnix1XExiUiuwt3Pjeo4BIU
Nw0R7AzBcF+H2AFi2gMFRW7rYzvBmwpuby9kW4+ykmT9vvVIObAp0+SIlPJt2zZut8KYKH6uiUQo
WXCFSUSM0CXLiXWUSjogZN0OH3eQVcUxAwgdJgnEgrMmcYYadnI5bAcezHcO/frnBnMRVLkSCPV4
165HdxT7eGpuJYh9MCvMxYjgzphLVWzmoFwLL701Tl9Mey+MAnfmXcOehbLEGnl8Y9yj3RbOHgAj
TkPOwu6ineKzE2yy05RHsKOE0xdE0ca83lGgnG7nGePlvTNBLRptHCTNgY1Z7eGra0u8tRGhyeu2
UPiNbHj1+z5L73YDGhC4TwLLI4l4OT1upU0f91UXecHAiUC1BPyC5JByRrOD1tiPUDYmumpwzBln
dR9UDgnGQB9MY+I/JZKspq6LkAMEmKautEQ/Cs+grHOb9ub37UltFiuWGfXqcqyjk48ksc9ykHTD
H0KoSWkRE/HGUAOg6j+fEouhQBOl37YjFXpX09Lb1ldwZ/C2G6GxcEHMcScu6dFTlDT//SDKQcxO
V/IZlSY7Jr4NGEcuLxc4MNMnvbVQAdPUW6zhdigA1CYRzfY9NBXzXb+cilW2uLI3V+8mkSFC0JDg
ZenxLZAbDrKuPjsUdIRAEW2PwYQeHePoQyDdJAJVvmbjBMdUFq/W8GVrWoJ9GYqWHm82CQy47rwO
hOykj4JnAQIBkY75y2QkaqswC+2ksj+HCSJ7JrP9udXDliiAC/jQTUz1MMNKQVRwpQMRcXXru8M4
sVNPC6uXaQ6y5bCa3kUW9T1sc1v3sBbkFs/wB7aSVuZrsOsLdMqzxrehST4DU5erC4o5yFnbrXUe
af51mqeosf5ihf8EW9LeyJcBEn78EY0OsqSwvDedm2jLM+bQ/FgrDgAVT31OyzGHC+tUbPnxfYQt
KG9LGEOv4DPtpy5hmQ85qFs0Ge0AkAzuhCsEuENFzwDn6riUk3+2HvGI8F84YZKTrfprzwGwQkBU
l9Zd4/qvs9S4RM+OoOJ/ZvUvP+pwwa4p9YdRl7vTv8rP1WCsy5M/OkxtWPFPO5PtrQb7XAAaHkfp
5Qhf0keawO2tfT4khBtIMZLvLzDV33hnnogAdtn/tvIzTzGSMypFC8/OQCWTuIx/0otZusOb1dsD
1X/xiC/6MKBClNpOJfi0jNVynDKQFXP7ytmpTgut+k66qAiC5yGkmeIwXSTBPvDi+Eyjj5js6G0q
EuXbUe3YVoSnF7VhO00DdUSoY7hN1OHwcaPxvV0yo2QKHCM1Uyvn9+bD6nmA8XYCZjHWGcPMGjyo
kk6ARTt+9K2LGaHqgdvCtZk2m1yzakONf1pACNNqGoUDtnYwsivDFI5HjHCQ3K3ZZTK8KOxPNWm4
Geo9pIfhS+S15csRKT2r9jVYZwwVl9BfvBbAohyd45Ph+H4vJ3vNnH/ZEtRvCyNkPY5g4oGPneVJ
UKUK1GTYp6SuBVTXLGqCM5HK4IoJz/i5kPX2bGBkLZvMqndyKkbyEp4NJkHMDoi9pswuXZ21jmqw
7WVtMbjGVf/Lo86Wkxd2CqHyPTYWxqtO/Tq2kMtjxE7n5wK2KRCz+Bty1eRzEAAGHBp6urxeDZnQ
QIX7WplKdzhI2ihUos69uIYzMWyH/3X3xfVi0oaxM/jMa4A7iLixvzPI5Eti/UdGPzZ3hLtR2JlS
0NTrtspxKkcb0oWebFUkUMJswBFssWLP2PoRPyIM8qyC5VQnD9NZGikzMVJkKVrrjxemUrzShcUV
z1iI4bGeLp9/J1oFHhAsLa0bKoEgko+WxmddKOpTqQKNRM3ERFoR6wH60cPv+izKWDHOPxgzIAD8
+Q+z+0/XBAaqkQbUhYszzgqLCQ7TArKBX47+Qq0QjIeUhSBiq2wCysL5PlhMIrvtkQwjg8N50Yx0
VhIj1Kw+VL7Be7uosQ9UUaTsXJupPKnYF93GYO/HZp1Drxn6isG+FQA9RSkiN1YkzD84E7DjTDcE
MbmyLugnWsdZSK73OKS4kXIGe5FOcQLQrSbQJ956Z0OAPFNcFCfgJeygKY5IJ8siljKF44cRTVQ/
EmXOOTpWujXcNi4wDdlIXdkhmwNfUaoSYA+DHSgLvPOfKkX6mqBufjP6/EPq1+0RXsSz3vedni7W
ehcid/mW3b2mHo5/+90m5+/+8VM/5E7J8r4WyZ4ramXQ5RfJt2pgMX1CCNK/TStsgWkFfPkkntCf
jDxyXOoLw1FnozxeKklhZQTqc+Zh6q10WEtDgRaoMLl/hYQAuj4gNpDfyosfNHSZO1Rxh5jlh/j8
1wN8tvX0dc1EQBkR+vTwkg4Mb8KOzHbdxHiSXaFiE/cdITldm6yIiVqMtKR6VkMwxLPab7pAEWne
65S+zqQrq9GrEe8vjlU12HC3P0VHN0qE2iAvOw1sahuWbSmSXtxXzWZZx8yjHNSKPgoQjzdr3ZQu
e6EhxEKcB2iscQ6qkUzBf4JuZ7xB/qyqXSTVGM09dmcFPfB5Z76St5NnOZ7zjqxnXM/2XvZC7z0z
pR2EEvmMyEiChpvrZ0ikCqdBqH/gmu6LZuzeUFC8ioy57IO3Nyu9jo4eKjlXYK/5jn0BJwctdDy9
O3FWccS82LP0n90k7y+CvvlypZ9P7axHIPB73mLLXujXG35nX0Vz0fKXaG4/PholeDkZIHvVFsOH
b52lPr1vY6dhlvYbkXp6ZqGYu84oKKe/e4rNRcNuBge7ooqgYq3My9iWZbH8i0elCX5WtkM6u4gK
RulbTIwmebzG1z5sCKCD+gGBW3rJlV40pyZJoy/kB+Hz6urZDvMnvOIFo90zaGDWVOdUN4E4+xIC
lAFJ2xHz2CD52zfqypU8hvNo0I5b43q7/dW8AdoajNK7j++HRSCLvhgcKf7seyBJzEU8YG5tdDse
h7l2iCS5tQFMb19vsUtW7tc09UfJyvFAwd5KYKDUNru3AlGsAERhaxR6MzqV/pKhRklM8eJxc5SI
tfMYCaf2bFwz2PnHHgJQ2RmdR3hvxVVTKbO1iG5dQppGHdh2cZhI52tAf4mVaR+WHlC9L3Y8EUic
xQrGgVgnl0U0z7nHvsdw7n7z/+/tykOMJGUqH7MvLDG6qaVnQtHh+CTmPju2gifKG+JVEycQfdLj
9QKIJCHuOQDi/GynNk2QY/yVdkVOt8AKCaCsgd6IDF+eMsFDpDD8NYhMPA9zkC3C7p3ylQatMR0w
9lEAeUh7+wk6y3r8lVHnOR2qiMH4TknKthbO7hySeW4i5L67fM6O0shmXsZPWdBc+Q7s7DsjvDn3
XbhTqsIIDfLhdIj//aZgsvcBM4SXWYwiNMjgSUu4QuIwGYm7EnKfNjkQM80oe0MsJ68GV8UCo+wv
x0UhKI6qzWXJCo9mDt/4N19Zfv92hon6koja+PXhf/DU8WjTymMjuk7zUA1zu1byxRwzb3Bbv+N/
bwimdjbvXGkLD9zepmBeGx6UF10Zg87RJh+16JSOru/anUjw8o4wmmDtumrHr5A5Yiu9TVRwmflz
XUWjVJm/x0yzDBujCAo68QIQDT7GxzkL2Q0nJuOHKuC28xl3i/Uz9fcPYvFmQxLwT/Yl2xwGF55o
040YaAZ+AKIlyqKCVtBiP3PhIb885sU6cGDQoVmMGiJcOI28KVNX2qPCBV+wbNp6BeceNc5GOU3M
wfU0qmjv/r9GEr1ztwUDkV+0pO2B9Es8+pVmSVEdwmTiRq0Zj40hYae9NSS9k6FDaFby7bv8FYwK
/8CEVHFFFtpz7yrsjyVlaIKPXHT6dkkeAsqIjtjkwNAffMwz2kh+Ybbh19A7WjSd+ImhIX4+oUfd
Zmq4MEVqj6vS9rS2mJ/VUDS8eyPxBgWAKK/jwO7p2oNOPLS88gtbTi1w/UaxNeO+CUZbw7UxGkur
F1zSpD7Dwn6jRLfLjcPVn3DTPtElXa8XPLN70/pc9U9mI/f8AnLpw0QuckbSFxrxqMQu+8qamxcD
27mBPZu/28LSXhgEPMjsf86qTan3R3ruVXoQ4atfs8TKp++9dQzP0oMJKvJZ7N1mG/M3eE25F063
0KKdmdQsjA22flhdqtFBCR7zzYzF0y7y6RCBmlzCFIPTEIrBKekqcjDhNGABsKsi//GYFLwgnjzd
FTOdDptnbRK3seZ5PZ9jH/qr5Xb79NIE5W52S2VjothqBYksjupeE/81fs8SLO2rxhk8ATcEQdDF
S3D2niDC1wUFSP9BGnzMLy0c14pDq9XjXnQSZ3QmqXHPlalBOECAbUovTB1jzfZwWQCqIfuwnpS3
vJFF3TehIqvS/7kt2ZF9I/qBnDXpPJPxExCqcbva8YyIXFF7xW1wrljTEWg6DXs3JRbu9UT9M13x
rGAzKVWIHqASmp4/iyZnt2DDyHS5eIQkGM7dtxqpgwEehdwFEcKDo2Z9GlZMZrq5E2Z+9661Pbgg
2z2vjAST9fV5uum6rA4YdxrgndGrjmGqVYVDiJPq8sH3bke3umfD1sKyRsJ/I7CQA5jnlIGDaPqq
3mI9YSNnKBY+Rrwd0l9rI8/2Zc9AHZ1ME5/U1Hz2UTL03BWSIZjtkVtDhusWkE5pARwRnEVgEsoP
D3GGIyTBcBwQ4139EQlsnkUq5aNbYoYmd/Lz7OrWK1kZ/2BqttaHzIaVFMoHBzC/XOrbRx+XxvPj
evLFmGCyGfLd71165KwoLEfbPSgSPrXdgYm7IQrh7ZFeIXG9BzzSFT0FBiz7f4f+n0XkDrndn0i6
FGSndczr0V2rN88oTywr7shvXovCoXUAPw0Tm7UNo40DLyzoz3vxZL1+ZiNoVm6dCafpmt20LUt2
4f0tInwkR8LvpaQqFAiFbwWObFHvV5Ej8ZDI51wF47Sp8rKv74xt5tPbyyd7+LgezJIVETq91GAP
7hWdUFTpaJfB8MaFFYE5pYlfGNohShMYh9X22U3tZyIICd2QpvtXNqbWAflQ7RTq7o/EdQ7zoljo
mOlp+ZBY87WCz0aQ6+wrqhMqvSeLRR37ls2jFhDkLkNwaXtrl1d2POfFRCBgS5yjZl4mmKs+Ip/v
0rlOIOT8XPapIoD8wvixhLW2xGFsGp9Df2XovMTorgsEKy+VmYdv6lD0GlWlZehQ8WmhNDh0tC3H
69awWoHNzE3HjVyxf6i8BawHUzt3MYRPUB6BiYlsjV0wwR0bB6ALnkVdQy/eL+J1IvRf2hdv2JAM
JMpJ228nA8pqPPSF0Q0FTbgF3nCa/hVvIbCom2DBpXOhGy2PVqRgHlFxc+c2gpbKhLEPHJZwdE4c
4V2MGdJU7LYLVvHZOWzI7aS7DPrnjMpI0/6+k2w3VmPv2/X+wZM9zCu85leKIaji6IJWWuyapc76
kmiwNxtcu4A9QLceKSjt0PUrEzo8vOGICVIAkuepQlux5ZwkkJ5EzgI00Q3vmEebYlnBSXLTXO5n
49b2yEL8MolqEXzwImmmwMZR9TWD4+T6pYL5HSV7V7XDC5om6QtCzkMOAD0VRPlGXRBHnkPFt+YD
zIBBPnlix2ojENQIzj1EpEsBHFGpBO+EJp8ywGtO0iplLo2NzGmwRp7MKwg3i6y4bB2j7y0ei7cK
ocws8mauQbGKKIPKhC82tHC6TSLiV019wSKz10libSebofdRfIyyxgqeTkC6dzQJutuw9GxEwILl
82F5R7PCGcFPsmSDa/GZtCjSM0OgthTi9e+56BSU1gp2FlORojx3bK9m342fs6rT3Ck18AaMMHqh
3wK3FYchdcPNLqx3o59LMQDrhokXj6ZfLvvkd5iAyeW0HRjHc7NByV8CsxYk7bR8QAELjcKjnLtw
ak6+oj7+SokvclfYFvU8fVF1f1zz6KbOmb6Kb9F6UysxX9u/D5w2g/5l4cl4siCrWAQt9WDfcAJp
x3rFcHOOPWlfOsq6rTEoBtgnGc+wJ3WyJZYBZ2o/8gPJ6LSxK/ssyMVNNwvqfCP6RuPOynSXE6By
Ndw5uqoyHkYhnCmq0vteLpmLABdVRqFj/1jnp5fT1P/FSHV6QvW33Heq5ZhO3p8rDZGloSPMhRu/
M7veQ7suiqI+axYs4encbtj1vIdpkpnLDapgQAfoTAqtEX8yqznx75xESE2oNk7cAAHyWLBrLd50
Rp/vgYt0qvVIguW45EmuhM6qhtnMGnUZj8egfM9iJCEzyypccvfNoW/3ZtKo28FCw6DX1ZOrM+88
+j0R3pEs8RUsVzu5uaK8NCMgP/iW36dBs6YQ0CfTqMRrY3zf2caWCHPZxJ/ysT+2Iy3vsnTPOc5w
wuqaL7Pf3731FyKHFLy894nhHzxanuYuFLvBO/G2UOGBXHDO/hSdzLWQQ7uKYDYwbwoFR2SqD4O8
plaXhZoUO7jtub4uBvy37aa/TtlbCI23UjefjNRACFcZ6igKJY8gTZDSutph58+r+TqzdHfM+Yzi
Y0Z2Xo81trGuzJa9h3Ms1lLboibhFIafmINjC/XDJdJ63T431DH86k1nOTsBsTwIQ6rKzeoy9TD2
dKJ3kirQzXmliK2QZUTL5xNOxDcd6ivG48C5ITPbqV+ZBN7SrfvvZf4gprGUo80hREvjLVWzEpfZ
LW5X4/AbYSor74zOvsI1RXkbtkMxF9+q76LZ61uxf5tZ4grR39hTwEaPLUrvmGc9sRwkLXkJ2Gau
Gv9LjHZzxJCpVAEaxfW2IWs7soirwgnqT6oP7cuvJdEyl8J8TCAcURura9jD/47ba2hxWhny0647
kGBwWN85iet0mTWnhcHEW5hvZL6awBQvYnJ7G73W6uEA86eGEYxIIFQQJHE/7pqKhVH5+EYOz+SA
n/48z00G29MaAEpx5r/6F8eFcWo4B6f0/w3FZVc4A9rsjsIBILpPK6TbpY/KHqRC9Msz2a3BDKfp
d/cNKj1jGCadaXeyvC1Rfm1/PKH2ObFW4HuGpZosmIQpNhJfBPK0uKeBWFm+c7dUXcogIK5kUGmY
/p310FBm9v41lcxZZKThi3LGRnvKjU0cGI/TD9mr6t8jtvlqHgXULIUK+W0x7mqec6HVuAmKnFcA
los0gMKipdd1mYWNEpiR5F6T4BVeDu7eL/gnOH6Dg20j7g+6zjvdl8U4jj2rz54eoBa9tbZ0mpG+
XpOvgapHBB/VkSYNOAxn1txpSA6VQVvL7fm5bCsGThz4qlzvuZjYHzH47QSD3SSfADhqSgSlEoCa
dHaWhvJP01WMP0PCYC7AGOZyTKhttKkaioUbpuEuLbn1dA6S55inSuqr78uh8PW2ZNI+P3JzAT5K
OmznDdPbIcnQN9+qN+PJ5hQHQbS2SukQ3exfJ3XkEjm+uZFRQWgOzQoCj9+68twFySv6Zq+A9Vbn
vs9rAM5i6nUG6Rs/kE3KNC5OtrR5gp69WBujZWXSWuulV4F6gEciwm6OeGhc4Yqf3m90hNJE2f9o
rOH7a1mL+ke8Sdnk3BL782eb3n9lfhD/PYbtmu+3HGnpSDGQw+Trw2KYtNq9b6IBF6ViIZaU7QHU
xlt5ohi7J4yqFB/qVp5tSNcdCD9/MrcXBgMH/zp8bRCH1qcgrwRGQ3/Bv9fgS/Z0NnVyrLq6NWJ/
tG9yO5uF3wybzgoUwi0ZN1DtO3O3fx3ZlqdgOrK+SAHiG7oLseSaM3RJY03pMWapM8bPjVM16J5U
oSn5W4Juzk3jCozrGbxLYFlAySd54HHqULfQlkCYdYsbxooygF01TbrZ35384Fvexsr3Va35jaG5
JPgwPqcgxtzAESOxwiJfn+FAQfVkcCUTrf92siKtmQ96MsU+rxXCoLzuY/v3vvz3mQI5+QwSfgcM
/cVDDCQceEosLxCg7o7Tg7S3HI+AXfHGNlPb62kTbmY+jow4+zy1k6TuQIlBb+IoIZp3uaSSuqS8
GMTm/+eevHtshvmTPxvzAz7sC5hCe/eJUFsu4gxd194PTKYDkW8jzXycxtiaeKuk69Ild/S9KIrt
gK4lvmXa9akkfDdpNGUnmPoxhhpFQxtLJj+LIXZYH4FCimqvd2L2AiRUhuJujMrOHHzfYaKO4/gh
hQa8DO+7fV/nsEJ1j9FFtE1L/NgiSLTdbf06tic/b2J+G13Yp3ZvypQ4ROXWZlY4ovjifJU70/+F
ixAhMS5dNUbgzq/6wqkQa9T/zocZhUywO4URfD0CkAPKhCZEAYRITEh9SqH1UZAfPtoNw2Uy79O3
QRcFH6tpWrw0wyYSejA/UAt6gURHeLw5Im3zzuAG8l3cOD+kR3bqlEHOAQ2sUDBPq6EdvIE1HChg
FpOwjF9+lrv6aP/zfaAcmy3twAIcSBPs6p+KC5wfPORryfclxaTFDvB+uI/eNVyapNLoT0oCIO/R
co4Sh9B5kGDCLZJVcXixkDnufMSNfV61fXWrlBOS8LrnVX+CpIHs15cxCXsFTOA3QxJoVDm6c+ur
AYWOiKu+V0TqaMsdM/+NVoG102oX0xXJFpz2bF+FwX2NUsWeFtYXR6aTl0J/MwF+YMMOCR3bda99
JNbT2nD6TqMqbVVBVxBui3K3gJElF4Qah4/0I+s6EE7A6dq4XJkfPgqvU0ssSRmma4i+Hz6hxZ5a
yzQ8FoUJpWNr+I7NuskonkXlRpG8q7Oz076luUqR4B0OkeFHQirNo9koRqZzG+LbMaf7vLZ+qogs
yS1gu3spAj+7j7gcOkTyDAoALlVFrkFA1bzxyNS9CjhBGggnDzXXbX1unnFv5uzvn8Z5xQJP5kE7
jtTiaxdQtRgG+WMMWQCOoTXwPneoHNy7gIRu4Tz8Ba4is/sdhj03oB+DwH5uBqfPpvGyMnYArTX3
z7nrWpjOFD1fwKcfu8LL7gq0OdNNSRBJjGT2y+OR2oOQoaagre9xAutPeRLLjfZqFrlXDK1TdOfr
A1XLAP9CjR/8g9jZ5j9NdxmJMIDYqbkpAXpt4mPdGwop+Qege+wyx4zw6DLs65PJ47T/5qD3/rG0
5TmNj2w05Hd9w8JB0uhPi/t3vYSSrq6B9Ed/9KQ3etpArpQJpovHmo2ZnrixsoNtQK5GAYXTkVDv
5zKKe3Kgk252zQ32xibZSMgDYNLllKvEi6BECgUTpWYWaWDUUncQ2K+E+Mr+smgWeDgP8pZmDd7B
rUFyAqmq7ab7owWVaqbLrxH2JEtS47yypz0GYNbG8igi7SqZBGIBuqzte5fALMvURTnqXhrh6cEo
WEGWUG/lpLYdBudGcmWyxd3iyg5ki5QWDuE7xD23iPvqr03mVfyUmtWKfx/FP0uEQLQDCvhZwAOf
vMf4LxbUflAENj0ma6eEnRMyZjqGelcm6tzttm8VMAgpisLQuqtwcSSj54gCMWt5sI2sAzDhq0+o
79Qcd6riTI8W6iD1smwn/8xOfe7wwfgxrLXgw16NF1itEJ/tCiMfaBfhBx7tlHi5Mxv0Gc9PJPvZ
00FmMYQ+xCUA93flW9ApmiIhiyGDhuo5GaGVbsJzRF/juhqrHbcuph2BdRaFZL/JpePGqel+tAul
tfGQYprIYicRm06oGb/ZPQxeY7qmFgV/ymzksWPm5JziZXOtIJKwMFDUqKoTpJ0ZfoeNX70mtohs
eqlyzAvq4kMpc72wLUxwLrsoTUh4nLr4uNvzyKhVwWp3bU+6VTGHBYJhttMP9UCBEP5d/2khTK6e
trNuw3ZDoJ612uC65ixfkI/5KIdbcLh+43bzp0he0HRns+cwbBh1tZrRkRNEkzwcHeYT7IYf3zsW
fHZE9G27U2D+XbdHVcqFCy0LXH/lPnpNaVhQpxHYu3YZ/iO+3wfGJKW+iTnqTGCiBG+Rs3EZ+7BW
L3KQpsspRFvEVys2i3gj1auKF8FEvdFu33lzXiPph8AJ4dyHO2q4efWbuxUG2j3RaSV7e52S2MOI
mR1WNtFNGzgt3beuZDEcK3ufnw9QiKNiGwt1jaDwtjRPIE52rAMsDYXYZy7rUJWQ7ckHrZkbpWVd
ezKu54MA5hqXSRcb5yOWU0AiE3iTBpKPkkYWxlrklLnq6XDgvIY102KW/DjsJ44QzSgSXXug/iyT
S6kNsugve6sXb6WUyAdt8LyOb8J36USpHxkmVj5kP/yHLMDiDPxRro9c5X/efoY9LdlmkgyWQZ3a
4RYWa7I9Ul1xzGfyUsjfqy634Nrb0MPtvzi9rqWWViv5FO3OZIGJLME+eDzbTIuZcmaIgQDMw7D/
w/YYpqsZR542xEfo+COJzUe5coZxSCTUXKchOdZGYGlVQ0EJ9xf6GQASbck2YprOAuTotzkBZV44
kt8yQyI9UjW1iGjPHvgrNhy49RDhgvUOyipOZLKin64N0AvYgL6i5r61zjYksm6D4UV0gUgri8rq
U9Ao1GyueSBW35uIjt12anPUa1z0zuNHi6Me5ModJlF00z/ys6jp/t/WVcmu6FwV+8zhVnXGfFRb
Qi1ZsDUsbqFRfHwikPVcOPpsaVXl2+GDkHVwUg/HqqcyI7srm0jQnXI3Owbd7Gp3/dn87FE9ILkI
nPUJGSO6ykRk/nnkkG+5sKMwLq9tZMR1un5/I9easAJse0JYjEUcH3zd+kgJ8lFNTW8fQJJKOJZQ
oPuHjNVadw6P1/9eiT1knSnQ4szIxngFZlYsN0v6Yb6fSMEUCgqNNKhFcSjrzHufgArdTIFV0f2M
pcOuaYeqw0aEYeWGittzqTlczGlQmWpw7UyqfcrR6QmOVpAip/jq8H03Fh1OvXryvuU85/OCbcu8
cMRtc962N8h1Bir3T0yVkRaMQeIVfPBeG8P6S3beVi8LNu1u00LMr+v6QokKB6nllgLQ6oDWxsfv
S3hUo4Aa3wVldq3EyuBvJGV0RqYDdhKOG2f0LJXv5k8ge04d91V6i9JKPH6kn+r5EEqR7BAwCqkS
IGYVDqnFBEqEQ+bI7uwyasgBa2GfiPPXve3es8BYicUw+J4RM5NcxWBmTSsJa3DVp+tlcnIYXCnk
a4stEN8/e5y7UXZgIKPC644mVfSEnQUeGOkHlUag2JsFiW9TJ7NWuONEk/z7svMDxAIbwDUDnrEf
abgWReMMF4V6a0WjEamd1aBZNCq/FykrMkE3HY6JfTpRv1sJELhTmAgxxQIddnJcE25nPs1c2xHf
82exY4SYCzYrd5dZVS8kD7E4RXbLyJRHDL837gKK4/Dzr1H+t42O9OqYcnYnhVeZ2Z0gcKRSHn+y
r+DHXg80XVfK3LiTK+ngCXFtSDQKouVs/3G0TgsBnF5TG2oQsRue94ixSk3lZ4/wv5WhmiAiQ/LV
c6637KdB5NU3yD7XsLAay+JJSx/8oFkkke1cLB+nDf5tqlqnZJHh5iBoM9aJKl7BVv0B+Vz/BQ6R
7B3Njg6uVPxwSpRPjYcobkpNp3lP/7vmi4hNoVP3CUAmgyEmcv7Sn/oUMiXiC72JA0PpTpabUSk1
eQlFOcz4vLEkMJ+YzwkWx4XphayUq2O/W5xS7XKJyhO1i7h11WkvVDiHHJHDgluY59EQQJd8COE0
ObX6/Of1RfBIpQKsgEHPz2obkrGdfNtL/X9moJ3sF1k1j6QpiBHGb194A+L3/IkmZXVWG8g8CdjW
+troiV7R0jxulnbwIMMuRrf6+avZZnuV1U5cbavxzbIJLbVsjtAu/rCwThwaL4CgZNd5ZaV+266U
71U8ux38lNFpB/kNHqGvtxJnHhetd2CgD5C2PsyJHclAM0euQsZrozfBqhrkksZ+iartyfqz0vMw
UjeeAA0WiOsijHA6dTLiwjEWOL84rPBeQ8DIl5TZol8e/fRFON7UBtiHrj8lDShbNrDqPb+Zo+MW
Z1/5uvhLQ0pTOjDHUxT0XXvf7bsKbGksvjpXxX/Z1wC2IwWoiKWLOTplO8F3pHx5ONEIxSXQkV/5
ExinwC9ieCTtEAwfpFpSp9ANfB69CbI08Y3TzILFslaQuC5Clmpx/DRAUYlmfasGathEDkFQG6Im
Pnc8vbpA3qSsA0CIfAZ45qjxgV1JM9SQSXexZyIUNK3LNe3wTqiBpbxSDWeqbE5g1uTcY6zDZmJa
5gDMxAiwDu0nDSmvxc4YQHysg7SkYscWQQtd8zR4xuCv7XV0BAeJkFyGFP7i1si5jMrXtFzeE/7H
qeagOLAz0Zolh7fHkFyT7rfFyWhDjifWYv62NZgC8oFwKMJyJqYDwAcodQ8lvds9sKF5vZG25YT1
/CizTFp1a5MT3kww7/bQ50xe6/fiPFhDKefVup1WWr02pX96V3OFRytmbIt5AQaZtv6TIM5/oVvi
s56xOpGWxr8GBsibaPyRMzX9GaNqsEIU9un2zeCzYYT7QLDtzn6R/lY0Xo3KmlT3vfruUaOMRQOL
urnnX2qsRi3TFxd7dBtoHeec0ruRZzO9vMz9q6xB23owvCUazFPy3bLdIeDNpKFuopKPqytCVp6k
YZsmBfcSQG5oAa21Yd56odFRZBfBRaUWrhzAFnfqUS4lB1Tqf8fwp1uPQmcWbI8W/0Nx+/aPDmub
IVPxVhS6jAVEwy76aAygGMlNLzZerGeqrEtgbSn4kXfVUC9+K0yQuGyfQLM/QEIMuqWILdzQDqye
N+dTsj0Xx/tLYuwVivDN0yasaESwIYG1mpcmpcaH0XRnAzsCtjGVU4ibrNEquQiDAGB1fXnKCVnu
T0c4a9FTRGkXaWKi13nDcp2fXmR+2U/lY+gD3REhThtRO9qN+uPDZIjT1bjeGr0phoi0vrK1bEKJ
OpJatU48IWbT2USTxBZq7yQrfECMRe7BYg1a4ceyE/zyAzHQP9yYdf/N/DZaKIO7pQqU/vtHszOI
ZM596eRzsdUf25wuUvEsQVIp3ROzDUFU1/Y6O1+OhvTE4X1lXMwTUJuK+PG/0va1m6iUqknFlOF0
Aiaio6lhqjnv4IvUwuhesAAMJ89ooR+jzVkLXMgO/vlvV4wvvstLYekDUsTgzP0UsBAO+ETk0Aww
bxxB36sXxhwIbcHQUK2tEnSo5SyAofdzchwI3N+8Nf7hqzFk4+d3q6Fi6LQXY7fhzFZfiE1eEnIW
Q21aQtp7quFUxaCdHa364yIC0s6yOjmCcml1BY8XxGIidNPTIrQD1Vxx8G2qQdy/YRFc8TlOyIyo
fbK67CgKXy9JiUy3c5+JtUQXBEQrrJILnBIE+5x0PzNi8BPz4o6evY7Bzp4RM5zKeQF7l2FOAl3a
STtgrnDxJtjZJjnmkYAuvtUPVFKdq9ljjhtz+3RmNeRzNQXR+Dp56//5sSGSyhkMoOTD3Ru7F87b
Lv7xZ2fEYQQM1UP61JPR+SgPv04p+UVs4BiNqlv/P5TEqFaAtJY3UQ+Bcg+hV3vcAyjeWq+QFfEW
mcEjNTATQDi10fHkrjj5o0fVvv86MrCSOMs3n6+WOi0J9bZOJYQK4HSkNO0olz34qQcY+OQLusiq
TIkMcpEKRar8korYVXjE9MwJ1gZZzFJtiHvTGWX2Ye2FURwvdROTDJepkQOIEtkF5En8sa532liP
bS07hyF3/Vk5r996QREtHrSYUinOb2IvMV11t0OIqKXNAbXDRVBAkt7gZDur6tEkKxEoBeg62kxR
1vAn+uPrVTVzMasgF4yjDIvVn1p/YWQWmei0+iJ6nizNhD2LW6QXf/6RsrRDgpTyFLblFezlAWaq
OVA8H6xqR927pV207x1bbE9w/f3I4reOd9nKtYKAGElAeqVJnqB3DKHedUkXGUA8vIEpg7/LAOBO
qQnUs5pxG7Ay8p9AdfVxFVZTmzdcPb544lsbcnIy1ARLCRNBL5OHK7D4eoXuoFB7UFF9KszXDjw+
5eYicILRifW6mRV6rTzCDhQwoRq5k3dTAGTxhz8oQcIQK8BES141w18Gc+dyOLLFVjxniJ1XnoaX
I7MSnnSfIQAl9BqrmPVj2aVzazBNHUe8f+Awizd5FkCb3KUVI6ayxO8o+sLSk5kQgy+iDITvFu69
+nLv3uYke/W6rxyR/2iH65zV2P/TwBNor3E61GPyjyzISdc6MQ/n3JDQlBe3O4uoiOjX4/7nJf7y
RAyjlMgWgiI1s0telQsXzUsw6pFFQWYRnBq4owhmXnNzCGpuofh+uUCicGE+qCOm7r6gdKQ1tdZa
zJ4Q4n5w6mPRnAwfQy4mknk/K/b5h8+EyIq3p+IgzX7kI75+FmU5/VoHB2+HZfB+3LYB3u/Opxsz
UjpZX7gRQCs5NbX3Ll2NmDeWhXxrLAxzRY1pqoYkD6aGEK8iqYFLxRFhEWC+OzETR37/Td6IzMUF
7upVwwB2woEJtazbvpcx2PPMaTT316MtV5uHrN48rnaK00qmb93UyTin9Ufy0eyW1GaRUoa8iaqS
2wDkISDEmDcRkwIHVRSf1oA9RRqbCodV3MNRW3qQzJCiZoQgiZLvu+jg/d3VTciUmOpUIKl66G2W
SDkE/vUZMA8fL88sGmlFVhGbRogVYoe8YvVIlgpenGWJ7FAshwahss+D3m9TXmJQLjw3BTQEI8EW
yGHcTzhEN9IUSiNirZwyWnWXpQ3s8ewM5dqIjCkQfu7DvNvfKbtkgZDFLOq3jH19jD7GuLXl3vRq
VyPE1ytREnRRDM2sjLQxGtii+7OdJWQnqE4IshteOta+r/+oZfm0iH52SThd9WwieinA2cWftkCt
YCKYuTgymG/R8r0KEuXrtNlrzmJb06M3+R8g9PYtNrqG7pPkyx+dMAqQ/9pgQBTA8ra+JdrF11bk
3pSFZX94Rhl38uCyZtR91pKEveJpks6Ydx4kLGJqr55/rzeUWpvZl48+yKwSTDvw4oUsVuhxllqC
QNdGyqQ0f6qv4lpIan2yxidLkMgxzveeeMxAqNhTzC2n4EvfvdxI046qks+7T8KJcXlba29Dqxze
CR5LYjxU8Dy2n5WI5SiPFnsgxCpeqoo/X9snTlUBZV48QGOILywXCFiRbAJ3GvuFIvqPtVK/EZPF
7VfdHce65lu7Ev8j74et5+sNcILLYt5TwyPHgzqi6zFAsXRZMwedl2yT4LPur9aKgWq03TNydcPq
8n+Ynt6BvZmVCXNOfPlyQbeyrrYMn73pkqxqtmgp1KPFoQV3I0KYBa1rWACowBUKsV6h18JLwErW
05gu0mK5gALy5UsWcHF+AKqubO1tnPuUxkKN42MsUCm2i7zug/oR2AAi126ahF0Ig2qwkIY6q5iL
CozQT6nrZ9Vue6lx61Ta/lCTWie7MWFRp6RqJUu0E/nJb92/n172dwl4zpylBWUwl3GdhkR6fKxl
1oeen2FrtqkOImgylJ32uAOuVPG4su91wl6nZ1doOhlczv/9ZTOAyQgyXe/5nhqwyMcv52M0woqQ
6H0pm971goBKNw5lM9md4pMqezj4CCXwpGPEY4k7cSujy0c6lJlFNsTwrnbb9XOMG1uCtGwj7OXo
lxVDM3JAJQo4lru+X0D78PNXBXoZtlPFhtifVAeZ+poNhNu5cpB0idmyNw2Muqq/2mFdk0qZjrDh
7xBYwuiYVhgPiIK269Pov/kY9wylA+mml6cbwTQCH6K3QlrgKinfaCXSFzfTseJycX4H014Sc57t
YYZXL4RwgNkJDDz3shD9e++moaE1MQX9kB/5FMSoir4QvVOZDOEobP0jVjt6THvF07uYLjrzIdiU
D4680xFVRgSQe7OSLe/r/RNh8LS0+nPpCvkFIAIoBBItUFCG99YUAxNc0+AzNhrOcKPEoupFrch3
Ka+Oc+tAj/VNKCRdFbIQzPX5yidNxif2L/PhehsjJvFy8u0fqQAcje+0LZlTbns02H0llt7HvPwr
EMvBkk2Q/X2qiaQN0L3ITKHdp+xZsezA/ouGysNc1DA0cBKjsV5Yxck3gLmITASPWTRTdqL1ZttS
sb5lapYQnjFuwD2hVJGUlgCFCzu8ndhsXW7Bi840/DpgMKv+LbK8yeP++swx/CDMSXR90g1jAZvg
DJNyOmds1TpT6Agin3rdJqI2i3S1PePXOryVG+0Xo+t/0fnhswBMt/q5fK+HZxV8+3ay39RfHC3h
ZFWr0DmHKEk6Qg1N6mU0ET0toNb4kRRSnFzsioghEOTnx0Smga9PtI/6iHpQt+nMA9cE44HEM8FY
PnLrvbxH2MkiFdnamr9JulzfQ+ClHRn+e/b5TbQPSYOaKr/Zxw6O55WuvIyP6uIKexDALP2d4Aie
KcWn2HXR4c3PZIoMtNE0hdB31BGnwVCexaI92+a6GN9yB09auiKmak0OFCKugY7/bLPkTvngMykM
/7+Ijjgy8V9mcZkN2ODuze0YS4y9eGzxqNud76QVWKhV89rFnYKFTav6mw5vnsp+/0lYurQ6ixVT
Ug4YwHosTWe/MJBHGAC0Q/M4XNNpVc/lqXWKxLPmz5yjt4k1ogiX70kAE2S5SiAv5Jf9bkr04itu
79OA95TMBEr0Q6WJVJQKcERjr45QXkUoPG9Fwe31TEtrX1hDUzsRtndRL+9QUkl52dIW/StwptP/
mYNmyq10KtJwdjpXjKqz4Lo1LJWzkDRa8NYSLcem57pl9/qgZ1gAvEwTuj2oauOKgTkLD8WbAbIT
yNY0kE97EkqHC97CSzDan82vpSWl6MQvPKWZDZBSTY5dUQ0ftSM1bHEEWlAs1AGrz4JUuTH3oovi
EOIMBnabedSwSA8v2fQrRbI+REAc6EIEeG6k4WHIq7/05RzA5AS6Twyf73uYi9ys1iAqOF7epiWJ
Vi5inDqlVXyQGrZXd+DJekYu2+tNqHeuMtZPjhQxCyoPkxQ0d/KY3NxJbm3yWQRvRgUIzzgNnNRQ
n2abCKo7SuMytHAw/9eLIdLD1zkOqZDOg6RRhEvruPAUDxLMZ6ZXDvAA8kXM2J530VzJdyoF/srn
kiJTDuMyHyR3njRK0gmvC9Qlvr7xeixaNR9U/980CXuD4hl+IEDOIKR/Wo46A6jCxgMQKJhLfwlX
Sjt+4x3rEphzYPgmP0iOKpexRKm4sFQW0E0udGvpYkTxQhsYEMfhJ2OKHaTNeFigjtFYaM8G9Hjl
bbKBp8HF7JsG3H+5DvbAHyj6syPAN3f5mkBLBuzVjACDZsQTzW/1MXkqJsPsoiRo91oX7Ec2Zs3b
v2ZtDI8ApVd5W/OU5a3+fWJfsGr1AsItyswFgmv+vVWYZmRnDLh6dbNssAjZJ9sj5awWgvZx87VR
W0FHGK0As/6EsJrnyW80l6NbzEFzwZZzz0AeqOTZsv/xv4IUmijtodc15vNPVtKdaTqBhG0dSz3R
+hoZc494yhUR3AXjioPQHORJWFqKNGMpKQVtjaBpNt4/F/c/7y6zjtdmI2Bc9l7xJVT1Qx3YwORX
9ko9NjhnturzJq39aL7JEDpRN4MqijIPP1zub4+CoITw28WZ3iJAM14NTgSJRLKQAkUDfGST+Fdp
Y8HLq2I7LpzyVba2wM7NVWXDQ1Daj7ljAipF6/qyYodnzLguEO7kci+JOaYH0VNySdmGN5pB7Ivp
X2a095YcEqR5tplNu8H1qTp7r0EwwxzyHHgzL1tO9RLtpZvlvVKlCnYhio+hjGZod8ST1/1Ve2oV
Ua2rxfuhDPXjOYTHP/Gsqjrxh2NpZDSRMf26brB4Vyu6uktMQb1Oq10Fbp1h5jTEk2hePk0IdisY
vEdHtk/J0wsoWbKCmtjHaE9AjsE9MZa9jfvPeLKDCgds/XdKIPJ/eibt7Li6CC4DgR6jL8otEmOs
WuwBy63N4JmvkvO+f5R6cvX5ngKZKyUq3BDhJJ/TNgO76pwm1jCPCXPnain91sV3hb9gRalha5E+
RICOu1CIrIBoBf+fVQ/D4U5UhNQWXtvvvD1XeEApYvDnQ37jSPcQI6x8ew04qrQQvjBv4li22zHP
VKDOGf4LsrcPtP1EqNsY7xYFxzmfVm0dTWP2vuSoQEeOZ4/U3oCnwuY7aF5F1zVtbKxckVcYWVop
EKk+Qc5fP+KYVNcJX01gFS+IX123rD0oox3c4UyHU5tIs8LoN1PDgYlmcufMnbxsAD7nQmp29Byf
qt26C9AJVXkWllGhD24B5+s4mTUPeWQvzbpiHLXoL9XTGaxrgbDvyYFQlPGBLaU/KG7GiBpt8aMa
0bD0xSDGCZCx4YaLdq6WxfuOf6IiBRbL5rBmFcbNuCt1mrfojQ3fBlOtcjQ5WuHhEp/MHBVFPfa4
2NMQPmm6+Zjp7nn9y1GE6a645BPtGSjiKQfR5LVEQWBP+yffSp0ZTUztO0U+3QURZv6IumIYq0tJ
/MGlfR36wNQjqbIaCY/czGo51lm+YKcrBIRnrPTX5Eexkv9DHIxWyDPf9itCv9WuValaROXJ6eNJ
BEzpz07HVO1K6tTGXUSOPz1IIQZVmyx0ANwznmOnsWeXWp3Z4mD/RSQCG9dFmVjEB3Fz+B387CAH
MlsaeHE6oMh5W14Y8wtXDgJC5Mu+R6aVhZopXrsIh+f7tG9uZKEtQRGoHstTIXS5yv44M4Xz4WWW
KD42Nr0ePSpEaL4NM6w6j6Bz7XABojTfJocZDuQ7ISC5Q+GsOgrUcNia8s1WzTDH3ut5n+HhGV7Q
Pzcn8VyxbzmIdew2dEGfBlNfCyUb0To0LgRXiqrxKHkMAtGiTpSOablgZvV7TX0A1r/XYC9q5cSF
0Mqt2ZO2zNbct08kVBEgKxe2tu0M8qmg5kHNUwg/suPiIVeKAlyImfZD5Bi8wqowsBt5VpJcAPvW
hNmqQ5Ex81jOCvmbkkrQCg/ra+Akq5T2k7KA10tZn+MQEDmMoQ0IBa37iVGFOl3tO5F6lUMAyW2o
fW1rtglLPVRM1obL+77rQPgkNzKBVGVn7knClZ3iwkl2RCTEuEN/JgmaF6wNTzdwCTZAcOIqjhgb
U57lKUS4aU1RwgfWY1PaYkrFbvb4AePrgEIHWc3as1GGys/bqLo9gkIMQYRmWy7uoPLXgt2xEzlg
pkq49GYCcN0MVjfkzpL7DrHJh1KSx98PJttrjqlFBX0XoeHHP2BRnA6SvXl5hD4HC49pX8T0mSiu
esVf+Gsj5Ovq34oYBOpmXn7It/hFgywxMMGKeEF5XP+N5LV/lgdJ2n8/t+harAR1abPB/vbp88Lb
59EodPy3bpd/qdiccHkEiOhVFDi2KjyWz0ugRcVBzk7DoDsKH88AlOYmlfNM7kXwQR+76Jkp4h6d
LrUoR6XPNkR3YDHMjcupePo6kPCDL2XR73Y05QMsQzeqL6Lnfhuaswcz901jfpf1QhYQPnKoIGRI
UEWo00OcaRC5AZiMlUo3p5jR4EAS4xg1vOlBAHpZx9XNgMrwD4+AxNpfIixdveXNZdkPhhsv5o44
bJPLjz+picRfGitrA7qZ+c13MaCUpFEEfEQ7/c0yb5GNOfk0/Tv9x9LYHZQMUkvC5zX5OWey1qnk
frdMSJUymu53NgXSSyv8tyjHVQQX+Px5Dq01Ti6+bUKpGUH2EDnXla4ueRB4Uff4Rj7r2YchhOcg
L+T1y6XWKTnYOPaBnYUMdEDBbkcBB12QhaORO+wjFQLCHjBT/is/kRwoVDtk3wwuoMuMsX6iCoCw
wD/sBZGT3dju6zEAx0UEkE6jcZkjre9JyqjY1gjTaj893l8YSGpkzKnZVQ1BMspJu+vi7mX9pDKE
LOkW4Iw4Jmh05opkFeCaHgU7Vu5C4DE8iAlT7nct6sj2uz7zKItBgDOK8ty6ARQRR0JKCJ3wqiWt
ewtA7HX7BGva9grtiAUT8IMZ/QG0uXRfLhTbJk3Io+140SNh+7YewRHKdnEzhWFXqeXr5t2hfFZ8
+QXHygdw7rMnsmSv4MLUZ+N4+l1JLb2+5JJTs9ihmaEcBS0+WV0xffibKrRjWylX6APZAImJRX6c
ifFdJt928bNChzedOPnJrI3g9rxGmeivRCHjRmyhP/y/z/nq3L5H395jqBg1Mv/Xu/MwXP6JfOw2
9RsAjeQKY3fjcOcQVK/1vBgg9SmvFrR0MmXbhu/I3PoX7ezJ2UApiae9V9VI2OsXpksAPjTVdMLG
s19tye3dBAi0cElyKVQuk4V9HkcUtTTmQGwTNgtrAkwDC9B07jJorUXU23eNOSjcB7KsrloR5lOG
ipc5ZRLoyllK/shW5e3MqLMgPj7lH/4pjYAyE3YNKC+xxporazw3GAMfGK0DkqgmjmWZVExq0ZIS
CmSU+4xtRm3ioulCyLB82hLgyIA5GEM/BIvAJ23on4lWaw6kI54p2PWvxbTRgG8UuwopbqRfi6pM
MmDT9p2VKQ1GZI2kgrfMzAlzZnGU4gpjftsCEZU3kp4LQLgIfO29bjO5WT+IXyPdXmGiOJBjveog
Y9KFakKBr5VPjL2Id/pU1yCa0t5LSczUPcMF/sLXF6KJbEJ4R5nLU7BwsQhmrcwyxmxyvI01GaSw
pzeFdw4+oIL5JesmUmXixvJBoEEA8EsKwh/fX5C5nRNVOw7Iht1lh3Z0Nk3UK8NyKu4iu6IiRAZg
GVMrtLUvzGphLthz0I4g7eMIgYVjgK8kS06P+KOuPy0yuV4QiDpMLY2urTmEZ4BtB3b0nS6mfPdX
ktV3sx27/dHXOmlBYmTqz3LFFcEn0W9OA2T3ju0va9eZOuq9KagMDElJ80fGOSB5WVoi3quHO1Cs
Jd9pVJyUlSbAoeryVM2hx0/VBHbElPoR5I71e0UtPre6Z4GLv9YN3GitEFirZaetBdxrB9zNS3w/
YZzInjx9e/JWmuokxY+3CI9VwRBLRoj6/yj1O3aygdfNcsCCUqoVyqlT54rX6vHyusBcE3zzJ2ei
C+IbWOC9t2KkE8F0mF9ww/UxlX1LmQvGINZSDPvBTSjvn4wOojdTWflIMG0IN3XjXAAI5Dt73qkF
cFjqkWonQo6XhED1mC0B0oc1SDZZwXGwaaDVc0rzYpLD7PSED1jvB/faygWNygPexXDOZQr+VJWO
Yvv9CTZmI2yzVB/N7yLlFjgIZOUiTfMfEi7XKnqHjJfAZBZFe5P8qqpGg57DOKD9toHpgCv8VV70
0vL+mP+Y5MYfxUwDfQZT4RHr8fCO6wPNEp6BQHLX1WhV1IOFGrFW8aiwpJIHEwR3vS/xZZ2Ytf0e
4MuS0ueUuxU5SY9m7SSGdfKrBgOCY3VbhFMQV6l7rWAD05oO++F/3PdMRTGCz1bvcexompE8xr/F
FV/u25UVtBREDv5SX2m4Kbs1DaXwkGItRyBnLBhn407jwZxARyEUr404YZNAWr+PG4VIO2Mk6VE9
MsUclv/+jo9SOiGl/R6uo6FGmNWO8EXSYDB6+iqd0KkpyYy7w6uQPKLK7uNIxLpFNV10k725Jupm
F5o0+PvukhsI32C3XvU6WIhl2H1q+3sq+vDbz7BYZXecRNabj1LRT0HJeiUzkyZ/erlgC9ipbR+g
hDnON3rlfQAW9I+smUZR5umviQkUsBoIWU72weF6zTZYw7pLricllMuWy5ScuQEOHzyrR3Myk4f2
IrZBlFt3UbnwgN0CkMcsIev/+UG96fDOsd52ajjVkD/uok73TdMtQLYO/wlu1kegb+/cEWhF1LZK
vL5hCGd1UNBCnc6FKAgmdNQa2jMFQzlM9uCmS68c/aFVrdWDGQc+mjX+fYcgRSBGyeQLd84XrZpU
3AYFRpkgi1AfWsR0a0TwsT2P8naEijd0ByNAg08lTK3y8x43ILDmiyEWugFuAWekdEay/lqNh5PV
st31+pYYAYGc3l01kyDC4C1cFpgaZOWGJRgaRzsncKFb+QKko0slzyoq8udmmSZA7HltdbomPDWD
EfSHdks/MEkKuParRsbqVk5VvqPoU0+1A88Wuw9CwrK2w0utWLQAvxTPa+TGArvZIwcbAAp1+vk4
Ydqo4PwvrTXtiTsxtwyf7cPa2U4+La//df1crZOmd94ZivUWf4gbaonWEBFJV4b02JcNGM9lr/hl
YAy71JRS4L0X78SAZnv9IqS4vVpvKsLuPfCUihccExJ7BT4AgptIE0qCBTTSCTcWlTXd9FUaju8j
xBjZeOHrifX33i0TvorArS3NsItRitS/Vvj+D4xTEQ199dGIY28FTNN6Jk2rsgAEjXuz/zM2hitJ
HVraDF0LtxMoVX5faxhfpYbFgE1u2l0PJ0sYgdrH6HSRfmEgbSg9tI3IP0CLc4NyB0j2erqZpyRz
yZzcIaCusbQ2nu14rPJ9bsBsxX9kEEzjFj9y0hbYKwRlFpkfUkGV3g59Wc/wDYg3X7n7Qa9xqY6k
DpiCKVZPRkOTN6FypcW2z9D7buW9YgcKV2fXOWRJ8uu2ePAyKLP5GjvEdCl/tlkzatJlCgDYqMRt
wbxGUFxX3S9jFbFiVYiv27udFM4mgKbPUcRLoRkK1jXqhu/usNrjEP+01vO5wGZBKoY2jauiUFni
5+8L1bB6tuPl//UdB2BjQycNvHZX0vfd9kxIDaVr/wb1PgUysUklxtgC9YgUD/DzjB/29DRIV1VA
LsgobB6DuKQ9B7Cg4C0PpKbNAXadhcLpGJRCLBd6ZAfz8a/HqV9FyMHaXog/4OQsjuMuc1pUqXKK
UHnJYwnN9HLZzZ8HwTkjysxi5E6LBMFXyRsCxjMt3+M2qGeT0Vtdn1+J82L04vTv4rp36NEl2Sjr
L0dcmfcY8GYrNwGVxYmxAHS57fFDBofswpCabouwPmNZIDdMMbd5XBEpvomX3HoxNj6jNwd42kP0
XloTT8XWRYx092x6wwDsM39SnLJXIaJFmtLevBmnlvWWhGuwWMSHQNJ/Dd3OBCWyJlaeAcEzTie1
Mt0HURERGfLKdRfP0qOpYrx7S5558QiMV+1/7qOkpdROo3I8wj11/t2B+fLmELw6mV0qsUzC/gO+
I5sSMyXyPHZCG5DA+tOVsVElXcZphv4Bw+Xg2mS3Wit/wZcWVFEEGfR1gOgFR+Dfm1C/R9ZhuSLE
o3Eij1PVF37Kss0ggghq87I9lxmIvXVmU9idqJyhQb+1fMeubKi7x2GrYPic9sJ9HR4Drh82D16M
efWIYRW8CzV/fvTLvrU1dIDBjORAOHf031e4+6n6L5m/GrnUlZ0MZw1wKYoMMpjX3R0uO1kCAQrW
30oFP5uWhqdkvQgpqwDyxDoYNbAJy7p+NmjO0wGfWmavVKCOyIA2ZFSg2Hlrq2LioxWW/AG4V/ZM
lBZLzMfuhx4LeUmG9UorYmktNjhcqkguZZasCQYCA7yX4JkbKExTaslWBZJ9o216e9UQzDSZrDEm
GfbI1I+XiDF/REt1l1t8BfECLqsoZkCHZuTzeNrERdWVFNQZXKy+GUFo5kxKMf4QC5Le2/PtLw3l
bjWRTkEVEgdMptO4dS8FgRYbcCDfk2vUF+IZBO18cfWlL9ceeNwRdJXcN7ACRbAwnfiPLgSBLIjZ
us6GOfReJsgddlapD2OJZyT7O8oL4RFiPuvrfgKuIZ2PPsFhb6Gquu4wKmYfoDiMROYCQlE/TiRK
ALhELvdact3kZb4V7ov2IziTjx5vXpZZRUGQfGz7IyZnXSvXzyeJi7PQZlYZZwJ+pc7AxVy4/KcG
ztCd4cgspbE2OeyefIGLdPaPagdVjm/+cmtX3mgMFkki2qKGoE6URL+dFNhPxCflo438K0zUGGOE
7pV7/CRZvIpgebTIWc77f5qMZSFg6aH5u7kw79Si8nQP6POHemxO4HuFxdD9Q/9XAS8iFN7iFlmZ
Tlq56dvDDpEfz8E74AGsMqFUf6/3ZqKrNovocJYpoDCZ8eAhBppceP+GxfAWUxZLACKnAU5h/0wq
ddnHAFG24frX9/BufQQuuEp2YdwWESBvEDwpGDc6CEImyMJH0plSHL4ReuQzFwZcwS4CO8kHBBsR
1GfMkVMmi1ZP2aTOl8xLxCxyww1NiYblNYNw//NX5KbyseF29O8EcTXLvRM4hqXDnTgNDnPvNT3K
3FD4bC40bQ6jkPFUy5pIgeGLzHWO2A+tuLhskc9W/cX2GF3zIYn6LqWrBHDBsEY9RrUlId3/IGal
PSIC6MhLjLuueRx12P2nMVYHyFwsvVcOfoPxuyAQX5pSgBi+H/wE2S1slDDyofN9nirJs39JI3F7
Mkk2U9L7bCHw3zJaFI+bL3M3W4jMgNzcYpDjvEMbiSi2+i9bWFUmUGZF4Ze7WEAhrTLPdHtnB1bQ
+a+yaRkpYuuMTVWd8iwFbQQLSJ8bsEAW5v3DgrQDIBijK8PV+7TLd3YPF7EXpUf+Qcka0IdyDP9r
MdJaZZJmSbfeErutRYlRzq4na6N0+X4SaN5CwNBI4FZi21tLXUHvTlgzHj5VAqqRqPq9U9ObRf3S
KAhTlooQvaNi+i1iVZzBpaVhKAsGIkdEkRuQe9dU4HDZx+EbAt7ZmnUtpAqCowiAettd405U8pGQ
KoPiFRnMvJNIAwDC/hfz9lWR54lRy2RKnsGUc9XkP9onqeUjEzt4R9+Ln7TKzP/Nb5Z57J/A3VXv
/DyaW7XLmedlZUA0xwPQOV7aEprhp7mLStWIYmrac8E/vPorZvEoYju88r7H7xUgsym0qYeNitaZ
pvqSkeYwwsrmn9s8++zB4Pc1N0yRHY9ovhY+qL3OrwPgZnnubr8Jl9/t/772cUCuXcc0s1lgEBxB
eG/fSHGsbjPXd23t59ZH01DlPOQwkMfTRAV+zE12c/2qQJkOspYLViwUvIiMvJTmvl/hiUCyBTgK
Hhmndu2M2XJG9vkLDp/wbEwbkGTZuhcXSx1YUumCqT0DyotfhC1wcnw0polkZlm4aPKkbhRJV1S4
FU+O27/e975DgGql2v6IYzYnXqv7RNQiOoQB7Ki1S4ly2telP7d8OPumUBpyZTtCVFE7rOUIAyyW
51UUCXDmAEP3U8Rzwd1zUX9RmfzJl93f6VzTRer/qpj45GqGiRsX9Mn6P8FSPq+AKwmUeWDhvai7
dg8TbovMUD7HsOs53ACmzKMc7W/6sJOGQTA1iPyvabYoRVHd82wNtrikH/FFtDhWbcHJTVCj4G6B
tbq5ZCPemjeccDHh6Nk94FOi0OVZwuRAzkjl7qNOyuRiHAoqHyjCktPD/2NBklRgulxmuIvE/BwJ
cdEohXEYTcjrMa3s0M/pRZhCuDgYIA/U2KXLjiK90uPkipaimDiqzGWXF8ZAEj6cFmLURNhIdECX
3yGGqKGRzOKm4ePEDfRGLNur2i9TXOTjNUxNsxYVmNcXAdimKuD7YqiVK1PIAkgIOeGzUp+9QvSs
lI17RYuSPSLbEy0lOC7tZYX3KCAnD+kh/gbjjhJYox3U5/m8C1Yonn0dfGZbepm+C65I35ALNMA7
DJ0mNMmKwMB7P+og57VxHBRc8zDXkIyXYwg7dNy9Uvg9rVC1tWX6WyRFWrvpG7R5lJZ43vs6h6MG
IddRf3OjiuzQc0n3OJBy8Jp1zoitqB7J4ox9Ia1Ioly0cAf1QEDu/eWmJEfcTOxbGbvHsLXO54RH
zodNtMPx1LyimgDrrmeKzzLQx3Xy4aZFfj1YSAXFrWdhdvNIzVCGVjBQhcSEMX2IJoxK+kX3up0x
Evn/It6SJsQHQGiImAwynrrPMzh21aH5z80JAegJqXLNLlNxymv+LwRnsJTKw0iV1LZ09nE6M/vz
Z6Loymm9rlqKt9VD1PiQFx24xB9zImWsrYv7AhHzrJ9Bs5fshvRaIUg+r/Oiz63dcRH0icPt05JM
BcBfM0MxzO9Agz8ZDlMaopqbhNrvToKt4IhTeQT5/WhCqsp52M1MUhiOoGYllmoCkO4n32tle/7W
p61Q18GcqX0nJoNeRHiDHR6lIxAmAPvhjJLdzc/FCZUc9wF4omK4tcSU3ogpxhhTxR9Y5YfAZxZ5
ByJZX+t+pTSbBqRbPHF/L2D1c0iqU+RJJDVa+aqmDYUcc4xtk1s3oJQX+yJTtS9d+Ac1h2klpZ8L
rhQG2RW+awke6BDAdkPd+S7WQITtmeWwX0LiWimR+LbKm5aqC9CXTx8Xh1mlAu9eKGUD9cotYaXJ
P6Fr3dbddWRj0eaALwTGQpFgpRhOCzZYFgFiVNjQ2AHlzMlnjCmXq+78LIadn2pQuq9oEenY9Gf3
agil8RpJcHiD93CInyQZsuNZ6ne/QxzhFT0iyvwwB+j3zvCC9A7rK/p9VosUyO7GneZziF5IkKdD
NWpjycq3lDracmxu4RnMju7HkdCRfQlAG+9Kxw5VoaGRGcu8LGfk9n6QWTD0IB04lIq0PGyLjTDN
SDCjqpUUE1pP19nMmbxmD05HyPyInh/c3JFBcAxNeccNil4P9xgbL3zDldPsgKXn4pIrj3Mhhp5D
pOaOkV6aa1CvSGzngj60ev8QZtUFYz2CJWP1TNVcWeVO8I3dEbD9ZS4EZCXW+lZoAgoESbar+23J
5g8W0tubZGlfB7MdG+D73OuRpLqla3PdeoxWEiVphMIGfmzJQaeQ0SsO+2zA44a8eQYfaZaaa6tQ
FnOaYZ0PQc7Ym8NllOQAdFsCco0M9Ji7S11RM8cYNpFLLX5R4EtOG3iKYbHqN0zJPBJC/XWoMCKl
7zWRE7hwsP3AvNMyed+uZeol3OHaGcIp+mnsnXPL8TSSflMeM1TgMeRQCjrX4oJWCPMxqw9SqqSe
MNLw7vtP9wvNbFFGy6sIaAKXJDdTXV1y8NWW+OYoz3DlE9oPkuifS/gRVfGBJHqp72wcjpHVdnq+
Plw2QiPBChz3SRVrwA/lUBjVXM0mdOcks8TMExX6uCK7cLzMZjKBUkUchNRzGHocSZtt2pcZVs/W
MhIxAGmxiLl5MVyOIEJ/+Vr8Csogz1TRcFM+TszDNw09bVKIllAPUQbAMcyQR1Frd/Ncf6PtPGpA
wE2GPM5b0m290t7Rd9aPNhgNhk64IuXa2QHwK0/E5qEkZGlqxbYVo+tu0nJ1twLtvXEMgNA2iTkn
nwUC+tgbhfWWvYj+A0hoBajKQwNPTPV1YTw9HkVdVdrEPE/mmuj1emXllO2C0AJrciT9VefqkvAS
7i82m2D1+dW4hBM2kCkkqJHvekXZk3N/lNMWNLp7K25G5dEKyK1jmlUW3J3cBniuJr5WW5Jva0PA
pQmRvHFoNMCqiv4aNvBQTGVAh4O0+vlQs3Dl4aCJaHxV/0j+aT3qmgr4KaaWn+1Iae9o11MtOETp
iKa/RC/PDb9lqFd73Yv8MxK5g8qeOJ5sONdCGRMmyMNljvbza2gttXrlyv2mjKV2Uixd/ck4cg7N
5WQBwv19+af5ootmIVfS2Vt1zGqrDvUArEtbrkXdS8SjqHsNy+6HNSDk5CuKBD+RI3QKZ098biY9
ErcLImDSlZyH09EsDCQWFA7eph4mwIWimYvI5Ik68932KsCwBhTmhzj+W25ejXruF34PmUTX0FFy
/kXquW9tIm3avKVXPNnZnFe8ksZYpcnVgAZK4fcB+wnnHhzpqIyDLzcx77UoM40jGzyYxJluF+uB
DMd7CjaPb6rj/wHAMhIZO39FAnvL/VfUN2W2PFR7MpKbNfQ/XytBm1MX7xcv9BF0KyyolPJaBD8c
NmzSuKpRsQ4szMm2lu5xxe42D7qsjKWCCIo8CncCpq5b9aYjP+zFLEgyowCLwlwYIb50sCg67RjM
DNaZaTKEjbXRzORu0aDtG/k9DHP6ZuupTgOxH1o/k6bN6YrHXXAj0tueDVF/nIxMJRLJcoEnNV0v
rcIzSf+UqA3g50OufgRimlSoymEXUTdHkjM5YyKW/r6nEqlR9kndxCGe0N/4hNOAqKSGCDhYIwCc
VhAGyuHQyuf0uGO+CPE88uEq65S6xjm4PTDuXNccrWyj/Xckm3IC4PAEebyQU4OijlS0pyIHBfLH
Y7qJZ6Vob3BHchQgauGvop/o2Fn86yfhiwPKc5FSgeerkVjoe1t35uyMdUY944Gbu5of7GjEAutG
P0O1elWVuTbWeeaAdbzCzayAxUtrUVzHZSwYu+SLQ2jdOsZfY0bvOAVoxp7g56BYIGdvs3r4b9Vh
g86CXIfNsTwVmGaU63RJhNmq5C0fwwhWvUe/WtNxLaTzaUE2zRGmnpEXDo4w+mL4/TicoFdGMaUW
qI1vZyrYYM5FuIVrTfiFisG1zwYrsrbGYe7rpgFvtpOofi3ex1eD7m7TSYQRQtXJpUhhi8DPXZ+I
Wx7NLCS/UiNWEemq0cnWu+Yw9vz6hZHOnIKjc1RSwNigv/otJeMvWPG05N8G64E8O3i8fyXUw2mb
89a+/Xm/Bvbj5KRBSIsjO5OeFyxPb/sGy8mNzvzvFz0rrbdzIEwOnVgL/D3DPEqa2HBtWR3oL/Df
PX1AKIClrNPdflYeVYPiglefZxZRyJJYi1YowykVGPfVgfuvQImo24ENoMKklrpBs4w58iWHMzZ3
eHSQ/VS3ItgToLynoMj7Zwh+OAqFk4ngk25Y+/9EUx2a6r39BgagdwO3EPN5IXfvpQhzrLAM0fTl
hMq80F+nUrbrnJ1SWLsqRqh+sVVxIP0LltXyEIvMPkhtu5+W5hNvtZajNAga5/6ETRp5OZwPGMvf
sGzeTV/SkaMke3BIBvHe4fvNPwBNX7C5ps/OlzulxrJgnf2R6ykUnIsjuHcSBXRyHd1HNmO3WYZR
AMAfgZdbhhMZJSsOhwSgATmo6ATz+K7YvBMSb8tjIlD27kqooUcROYCcbmgWbiPIT0pfcEpIpWug
dyuWyqAG/UohzX4TEmTYYqpPXjFxMNlbypwUIZWv6UWeg91z01WFJiwZxfVEhzNKx7ulpuh++Tsd
R8cHZkS9HlJHhE8W8mwuzo4DCjlN7wd/Dfcam2YMs/OqK4h6Nei+rrWuunS4GutTN3bhMdH0HXi3
OMLxxO8IM6Xjeh/vXDHMklDy5nwIyUT8I6lMBGkh6n/eVrP26a7B6tqhGMuOoZrOWkyxf7DPgU5L
dwtehF6sTvR96qD/HnnRyImgQtUMRwznoeL1J8QLhztweH9TbPa9irx6HrfA70BUOUz1RQGHNaAi
wYJfLe11tVUa9icvwdx77yCB9wDzDWgNj4bCgDBrW5+0MT4TmNqQtMQtZ7/7e9+jD2EROnxj3sPp
uD3ZeasqulqPAuZ/JsolVvsXlClk7t9z/7ECWOWzLK+9F9UuiVezupAfbR87Wd+Vl77v8qAfBtdq
Z1XrDV4pTwz0wSCTh5E35BzHDK65k53huzqgMnE1ZEgy+DOKmTSyRuoThN5MQvk60fBFVHsVuT/P
iYzoeBfRobg+5rJ90b/F2W9ZhJ4N2WDc5rcivRNJ68WTeOLOpFh6zt9R3C1ahDLBDetFhWwDrgsS
EMjDPU9UWicwFrloixGD7GOCUPhfp2NrGsyB80CkdB0WcBlrNcWQmjZN5VazTFtaCyyxe17fYHHS
Vu8r1yaj4yvMvIU7BVRhpAqnVPOzigcHOBLsmluu36vbL1uzsFJGhc2WXKfVidVSiCkIObPZtHEO
OPAPuVRBgM76PtkLig1gVPVzLfly2K/hYDaFQLF/m9avF297rk28blkDkY34suRImPLMe/71XRw/
p5PeUZEPEu3ob/S/A6jqH+T7C+c4juNvjir8Tj54zMmUC6P46TQDhz4x+QXA49oHiTAD+DW4v6ys
/z72UrSX0vj5H88Ztv4NwoS5KJtXrp3XMcDeY+V1kxoLR2PmJRsE4/DvUdIUFoUS9ZVUIOD/LMes
Y/aU8vkssusNHYRkkt3gMu7BFf4o9LhfAgeEUF7Eumbpz3xJJs1jCna//6Ms06PHOYN0jI7o1/ss
L4mfoYATJPhBryOqrFH9Q9JIDE2In74fld3Y6GGth0Ov8UQo4UiyKucXo4fgV0B/ix4UjIXRSbgN
s/XxgqoOzxbuqALPAwDqiX3ug2lq/wfBEWhR4IyJAF1uA9PpAiAC1Hw0RIKXsbHhC+9V/8ADevxK
NIV5QWGmtnf/VlnwloEJlncaxl4wUrBiTTk/uYatP3iZ6VZ5YO8fTg2/Jcxw2NPRPxnLMjEQPNj2
hnOlfKz5mU6TxSP+NYhekNt3psGwprZ1VXWrsaXtDUcqULp3vbajbMuBcsMQd3iGjEfj/qDxRozW
DMyjf+GWe2oNgThWet7BpYqFdWiTh4dtIplWHjV3CQRaGfgFWAi6RDSaeL4Q81RFOWs4p//paBGc
u3muKIKP+0tY1MmJlc0apWV+nz6TPFzWvkWErI+K8TXWMZACvuxBTQb3LtNdVoSOh4vYN7Nte2oQ
ldBzBOluAA/OEKD7RN5kueN+Lrr69Q5j+XZ1ucLo66uE9a4oAjEI6fyXZVhiQUFL2rqgTPR0avJ9
hWeZsmA4wDsjJBt/IfoVs9x66FMOQL165jlXHkAujkkVpNGkNwlt/t1tq2+bpBun500fLPhY8Xzk
85hNJ+amDdqX75RALTcuAzIEeEzAHNgmoBSN6ODzVctGleKAU9a5Hy5nOS1303OE5tRQkNxVgpIi
p14Zc/rx/zzF/oAIl6u+leWspCIhNpEKlJ3xK+1WKGvEGkXUTPKb0KnfgjcqmQp4unA3ZhCSrv1L
8gur1PjrFe4bfwLZh/PbVzo8YGDbJWd0YAlHIsMzVIHz3PR0lX40I283fIoooA9/Jc/maDEkHSYu
pgrSna3TqQbp+UIv9MoQrP6K7OoLunpt/nlHYkqO+atxDWhv5Xw+2YOBwkdVWwWyb2PIKSd22McF
wQAPPKsf5q/+kGqYwoKrau9596J3TREfkDLv7cCc278FuPmm31g2/6JE/EjpYKx46BONNaOCYCRn
VdZc+J2kAybKyGFmczjV/lGappgmlW/Vr+78oWKyu0mXL9pWjNxmRbraKwe8MNwPKironBiHWWQR
jA5yHsLlx7nsE4SI0Cr05+2I7FoQBBA6q47si14nx7VjpffJygHPTw1TCXAq8oBYsOyTKzse2HLS
YH+IWsjUh707qoAxfi+WnGAmx2mxqDVjr0vEanIYiJ85bo3AUCLDS6poi8QLeKMOp2SbWydOLpfi
lVVBvYeXRDcWBqLUJwA4lrdy/WhSt/nZf6eYwTvfkqfy1faGurC6f19c4ozgzT5jVlTuzxQImDSn
VFUNewDdO6/Xv6mNRIKrWU6kgJ0odEGIgfYFPLy2WkmnzF41+dzzHSnZTb36kc98xKvRx0/l1eNh
zMYQJXz4/0d10NTZQ1KVEwqBg31JyzNPU7hMwpp/sZEnvwPXFH/PLclWw0PT59jXzJTsSRxkjioY
OiFUPqp45kXpkJGefFRVIMAhCkdc/ZlD4e9FjFNLi1kufOlRjAhZ359Jj+GsvFYjJr4TdgkONUBH
Qdnh6jcwO6Pz4SCedAFp/WHlDh5WZxZrJyP91IquHExRSfzcECsPLkwaXIBr9ahw1t3st195Md19
jSjLSzNtMYkwRhfyNhiIAzPD0gt03haupABMZfWdD874P8cX0nVnrCS7SNQGpXRej/knyRfS/oue
v+foqCexuUuOKbj3vR3porSqQOzs3PzrHnl8EERSW/sXDpwEGhZlIIqNfjYc2woafG2jdzfMRsNN
Yik8+/0q/zrDoW1MVs1QdVtnfrpACPfhUrgjUEOWysaspa4erp4lUZQkS0d0ps7tFUkdwt26VvQl
nc5O1emv6eSPfkzmdqgdApKNht9lpSj+k7YArlrfipX8uHkfJXwn8zPMJe1D1KcQiimzC0W/rnXB
mYUIA+S5tlYtnWwhN4wxbF3ivRpo+GHEoRpKm9dqMyqp1Xvc9J3GFmaRczvmoZn+zkmX6fvLl/Zk
L4UHGhE+F+X7IjbUWqvJ4it5ANpcrRy5BnxnlnrFAV7JQ5/8tcUDRuCnOZ/yduJRfuxSxtU0j0pw
uQx34YP6pEUnzk5Yw8b+BlCOTBrJZtdoZH4oJMkyzasaG70xjl2dT7SQmw1fxu3bzpGXoBAVfq6r
FalPwuuCc1jwsNYvUkcIOtQAhzMpntBr2E0tKBIO2409QO5JCDinZUi2q7mUlWdSNbRZE2zFPVBm
e1gvrWO+TrTCR/C4EsxoLT+NpAvrpE5bzQLCKfn1gGdNE0DD6b2SY1QLctSIokK2OcEG+bI/wcU/
5Ie5D2reTFXdDmJL0roZXd1r6Nsil5FxLvxw2B26+iHNdcoaJUB5tZ58gndRB351jghsAhOLZVBX
N37ix3QqUiEEVNWDEiVlyTwIgvvbOstFrKI3RBq/McQ5T0xXG0P5YLzFl8+IONhK8YwhJL1EQWEy
uifPBY2JfYQlZB8tSfPUGmOBgmS/tYL1IxEGfFLmTmmgNYDsGdtY8tku5vgKzHGl6rmHhR5CyE7E
2O3HMaWKyK3vIbfqolSdTpZQCxxKWcEGHk1h3fEL21gnlnpFPEqpf9up/pdsKIjdFTZrgzqzo/y2
Uu8F2mzVyUkL6jmxi9pxURELzmffBqsY+ssEQTDXzH6won4PAJ60iSz9j4m8CtX1YfXmH6kJtoSG
cBImd1MWhDQFgnSUvZxYYu0UhBKAgWuzxd4xhtETUyT6K7cWCH/ef1bXhSni6+3kdWrNvcaJgkSr
R3jb1b8iE0s3c+bLzFnXySbd/zph4FmKUTIVFbHxkb7+MbHnzb2TapBSCz6QIhbW1DDGYD6U6KuE
xM0ouZI42VwaLDHCrR5VuGYtXyiikD6bDMucmw8h0k5M+/pzGYdLOPb+oaz9S/nQdkZYaXjrbLag
NI0RBA6KfAjplqdTTZUc6rv4/LzuX+R33Orgz3KSVXyDNcFcc/IkWbuwu3PH76721USWeM6yQ9+F
H/cmYlEOw5UnkimT80uatlEQbkjxl1kksjy1MFQpZ401YnQFlnpaXeomx840KtUonfe8MZwXHmzf
OSlXjMy5BkhY3KBw2n9w4SoRlDfK3XbLx1mR71I0K6Yo0BT9ysVbQQ2TVxLMSWacRQU81MaiDlK9
Ut65Dt/vqC6oRx87pGtdednyQto2fR+IRi7fPaqOZWF7in3smQOWatQJxpI6m16yZEQsnM9TIDhL
QDZGtxSp71jL1takZsGqu3Bu0wusM39xpG8e6JaG30l0Rsc9afYJ1xPHQIoI8wEdPDHulU5qdG7p
YkEPC1ReDSru/qoL47NSDwx4SnAdI9Oe3IBhv1uCghs3LeKQAFt3FmwH3EWLU1KPqHBxfl3jQbsT
pJgaSqULHcsYp7iug3VJoA9uP6nYysmKedth3RooQXJSIMM0qenrrcVy2Kve6m1J3HjYOXXo/gJR
HTa971T5iVps5w8RxClFVlal7gOFLfY6J9HmJVheOmaPE9WbXPmCBuEDML5Rf37yFDpt5nf4Vk8I
XCA2pvikaXEijgHC8tmksa8jNz8TGaoxSayErW9UKTv6lqPUFHTdqBJ5DbWuL9z37CdhYTWaM62W
dh2DZAqUD4GqIKjOf42qmhNrAKX/RbL4KeJuIXdoCvJg2ZlrXQqmpwndP2040ZFLKFFmGt6nUw9k
AIwHmMi6ehrf+hR6+ImTtW76/bYt7yERawgljVtjbyuq1dEO7vffNhhSNBklg2DiPZAHmLqAmVwO
TQMfaZFh6uJlhdmT64jp2da2mLT8fkPD6AwnZKR03VAKk9g15p7tsrQ5wLBtH2G8qcnFxeW3c/Qc
bCCQSDvFOfoYoQwmKGrQRXeAWy3wWLUy63yNyXdagGrFMgxPkNjea6RcjDvqmIz/rfDJp4J+U3gy
8shg8ODvCy3eaF6VdG1koRR5ceRFiuwiQqi0bRGR3nUypwAcca2ntROvePaE4HtgrOtwCIlZT3KP
gGK7ZkTp9JhguTeSu+UVo56nlXtZfiReRre8pgl1ZDNywp7ugpNP5BFGc6FLYl46Ql3S5kRrgurE
vF90QL4DNwflQ6ZVtbOCb6BbTwYt60HldArRWkee36ILDzc0C8RzvszlrFFKj/Lkph5SVQQrh5h1
UrfaygSCs2R+IeRChDiJjU0O8aLKTzp5WfoEHrTaaGHyyx6w2rGiIu1frOoxlDz7oL44QPcHGeM5
IzNwY3XoOwCzYkyxk/CJoJlQWLtWpjQflhqZNDE+pAyIiEUOGdU/fBoL9nuCYi35Uj2j+zs2kazN
etCm2DFhbHwV/zO6osJKsV9rwJ+vThWr6VRYIl+mDT/OF/3qFBXiQWj7RRidPuSWVu4U/R8Ial/E
ruN4hIXL1PSAgItlcCz6RP4rlnWuFmUIs8HXiG0CbsDBVJy3k5Qr9aZqoFnGEkzD1BHJt2XMNJ2a
MpFemDXvjfpxTQubHmLUo6wiuPqPileHDSTforyh/t1MqyfttUzK/4Iv8bH63VczMK9XB9R3NxgD
5Q0I1wUQ7AFzOLmEHx8IfxCEgs6JO572u2y6IJHxnJEoUtLADXIbeyHMjoeQq7Rr1dzfVmphhEpw
N75wmHBJtUHvSBfSG6jjoy1BA+6P9a42CWthrcVyRNGptodWnphMPUFlUPKP1t6wD7pxMku9THVE
TQU0RUF+pDbHgC4iO3IyxDRVs2/G9EXauj+G+UuxUUBSMHAlPEqXTHRs3ibnANPbM1+YDUlpwNLN
Nqp1iZstU4DqEU4GR+A8nOMHtIeds+8LbbG6KmmcPDUg3rh4oGbhVmsOBmc7iZj4mbxaAdtvMIYX
UdIiGJZJtrHrLAqsRCb3Ybw/ia1ITvY5xm6yX03V3zyOHZgaQmUffNdHBu2sM4/TTVESgG3nsIQb
vNRVDcMon4wxsoyA4CaqwWlnoM9u9+DzlXlFEIePCFJ54F/9IqkNgFQesiGdw72VxnQ78xNi9MTc
rwncsVq1ep9ZCT/5fSyMKA9UguCDW6mFIZ3uKneFbDMDge7NV4iS6gSxwWEU8aQOLQAuGAbwMwxF
fJjytRxIU9FTtd9K/FXy9djEfXI5VMoI95Sr47kyRH/vX0K4hd3LJCylglzK5GQ8MspJAA/Of1Zl
uwt7H/hA9MkW7Cw02C40vttI19KBL+E6MQoS9G2/0szZeiujidSBA8Q8sAVwNH/SID3BIajs0tQA
k09p3SCt45o38L+ER5hObWIlufX56V15LkMCY5mT/sR/VBbBKu557xpRg9n0CluCFGGwXgMn5zia
hbxzTP6AfplAg9Gmm+LuHUBW7bEmNJg7vUjM/kwqpXQR8SlLrm4bVqTF2qFDQvhCRLMMdYzB7hkM
5HTOWqJPCrthiypHs2SVpq+qLIZRj32NU0wab40ydx4Ofdj+cDzU9GFEzzsOD19PbTzBHKkySFs6
3FlmhUxY18xxSVlnodzbY+TqU3HMa87utIYirtuF9r7X1heERxijXtRJIfvcztiSzoC2QoQqaYqT
awMZoDOO7zVssEZK+Zcf/VzOzUpcAMKnD6RjioS5VwCulgAf0vAHS7f/gXAGjMaGTSRuSU3ELOr0
AHGi16Ixz44MtdhQSdTmYZejcR56u6cTkNXzIRtwGsdf0di5Fl2MIFL/9Xz0BrmKo31gAgcErJeN
taqDx06WJm16j38RYm2rGiTRo5SMacOfKSjldO8MEotsrqflx92PPxdorw3ia0duUSj/hDh5jOzz
zrV2hjmfNWE8rIg6T1NCUDVzUMRWqmrTBx9XILDF5QBMq3sKRO/ZmAu9elBgOB+A7b4jOX6qSi4r
KifiBzHXwoS5Xr66Gzi+6vnliFUO+ZTcnQ7Oo87nre+021bi90IYjiqkOe8DekpKbcvDbOel2o6X
N4uAR9EYlkNS74440ihWmS1ZC9HfmR8hu4LmrwRN69+l+nHB7WJbAyHqdaZEWY+rCHCwMVPqPL3c
hlalP+rxUp0VCMvX3JcEgaL1YXAG5fAet/O7aUDUaG3AkklcGrBQJQqRS2APL4mEDt6MfURx8h+2
DEpgMiN0bzXNyg7ZbmqIW12mJ0i+kqA7sLa4MICpStPe1SxHpYnWn6nuronb2zNpiPd8JsjzOdOu
ES7LDwYY+muG37aD6T0iFONVVyQbn6FbigReBMZMGR234RPa/dRpCxcR7w+xV8jfz3RzWnUsLeNO
U3Na7He1Q46SD3dfqPIPsgmkkMSgDiGWgUvvm7pqGpmH8a072pEuNRA1BDJG8sYTxdq/kRT9H51l
JVuvJRrp9Q7SoMjMUT2UA1CLp+pel9dDo+p3RYADKTokQITe1M26gQjrNoKgAwC3xs/8aNP7yZTY
/R2b6TtvBVleKatrarQyFgK5Jeppy23EgyU7Ti1a2dymkaZzhHDECWBt3HOnq6rH49741I9OSYRE
cXZVu6UQD4SG6vs2pZTHMueay58SD8RoieUvs/t2HggcdY8/Rc3kbuPUVWcPa7noAZBtaQ7KtdRJ
kE0DDTbycj5xc1ykLvUfkU/iCVKaFTCk5xZQGXrtl8gie8Y91vlC9UOphDsfjwcEcxVvTsSTyuQP
wqQnYXfs0bATG3HqxSUvAaTWKBPo7MFgso2ciIsBVFsZVQuOyEgd1oM7OOEvrvkU7lilgNOMGZXg
OkUCjDRXmajTP07vI9gI44OpSrJX4jATtUMYvxIHb9b8wYDNm5veJEWfnNt/MDAteNMjv3dUoIFj
TeEdmeesYvzrNQHjYhrZOEWZjIYOMNlb5DfANv6YJNe8qEAoJUVZJgIw2hVe+ePfXJ+59Oqq5K6e
kaOhkK/kBBGVhE8K/En+HQGyRlq1PN0u+I54YxzaRqrw6/MbFTnh/3/58CV9G0Y6xrdwS1wPXXh5
Xpe9GQpC8Akg4EOOWjwcfQYGdzgbMiJ9Y2pSIMm4E5TRDqiNyH+UDG9QpKPIwjAJevTQTP6RXjmc
BT8OpUuOBo9ShHWBvv4KDsFsMW6Cqzn6T3nfPrYIBg8JV8IAT0pA68woyMn9+AnXNbdrocPruJt0
Zn5uQzm6SB3JCoVSesWrVP46K3fLY7PVRbv7L7pOoswYznUm9g/RbIz0pD7bumY7l/kRfAhAg1V8
q01APw9tdLc0uLXJRV3FfoKmgbYXeNVLNj0sRnepF30icy3iutxG5wKGvzKhv8AHi3JXUkIK/2L1
3r1QcXY2KdX5QJmPY+ApwYAk56ahXc8rV19ARnMEmxYRP6sYPKBaqOOGQGDTq2H7IQGz1ctEmf8P
H7WYqd/+Bs6RN+tv/xerXX4U8EVnqWzi7/OZTcD7s/c9BVwUojznTu7wmbUIgLr4hE/viQAonvym
iuhHSoxsbtZU9JFA63uC/2yV3NXHAQkfKkgbudYuf10tAl1k6kSTJBsNrDc76IkftsgOKLSiRRbf
wkNAkjIb9ku6vm5iUFNi1qpsL6njgcl2hk/QTvSjIxWYdB2oAKonDkxFHWvQBBQ3TpWfC7Dr18lh
ldzW28h2G2zuy5kEiW8xo99MDm9BnT+iyn19XY8XFaGdTJb/wjdU8e5Cyka/aa8i6MRjq3X7Oq6z
C6tM5/sbGWCRCa1SIyQspMNuP2hfwK2M4GoSK6Y3gC6RcRLJPa83Hom+FdW9+PMNISJOl6lAfMTY
qcDG2VtWdkX7rxuAVJHn9Y6+6P8+CQ+w0Qew5l4cYopubbIu8SIM3e3edrOjinRqJSV7J8Vkgkvj
Mmo8rl4pC1abWx/ckKs3jBRjsS+Oxrb7w/E8rWE30EFbpmvb9ED/Qz8apF8n7CdVpw9SMPkCXPu5
VCzXyVi02MmuU+xubv2u1C+ukZi6O3u5667PFVyIZ4jzY81UO0IJMq+ycCLRjSycOEbs8UV+4lxu
KxtWWV2lIaUCThyIr63H7qRomjKqaUuAGvd+arRsUuVkDPyT7NtvwLlRKyJ//Zq4ZueeXaxs6TH+
dHphJz5JFe+1qecXF5CYPQyUBq7bAsVuEy1K/nuh7hXD/QBEczz3VF9AZC9sp9ObzZ9J33FCHIkL
AElt9UutS3BeTzFml7IqZvEkdAovYarLeh7h/um9V2kfB5CVDIKxwJ6/SPTRXYlz/K4sbfq3aPVi
SvsKH/tq+uX6PXN2kJpHw5uoil4nmsWk/oSvPpgs5cWZPTDMn9jwUfolHKlurdVRctmG1nixaNqn
tM+2iVp8QNUtfCI6MxluN7YtDA26Mwk6N231T2BOZaCabGV5TBiUDj5hrEoWcIycsSP7sjlDCL6q
vNIL27rMbdqZnTr+O+/kh9wpQXA+kfEFQW0jynJONeKx/GuODvkgsKVFSm451FCxR19+EEDEfxcp
gZoGwObejS1sKChAuOUHyOju0zFWlSQXkhfUs9Yw+ST+jZJqS+sLXr66OT4BSTbbc4TUpff8azQi
qFNBxIKlWf2kXILCe5Fn9RnlpxDueZ40yDlpV2fAVI2rwNFSdgRnOzv3RxYzGKo3oSmopQY/dEpH
DtUvY1G/x4w3XFkq3p3R9yByYya0fn4fdRpdJM0QGl1crw9wYkq1f4bq3BrfAViiSOuKmaEkzLsh
4NJ6WQ83P4gmrG9EbApEZ0GruH7nEV0KTg4RnwnEqT+skCq5opD7wPdTZU1KKY28mEOd7wIISI4E
YSEIF3p+0aJM7MHahXi6rRZgmGizi+s8UOfmsiW+SVxoQjxC7vBZnSWyXYCGiUDpXqOOhc60RQaO
Ar3W0E3R66tAHk4mUtEGhrERc0oMElR9unZm+hgfLpbTa5MeEYi1lPMVxGmPGq9sfPoYAbaBP0rT
dtPvm3H9HKd0OZ1bJSL/TCy3jD/3Mz47D2AyvFtU+Y/zgJovJFv+fymlmmOALkOcio/0sfAN9YuC
xQHlXMlxGQUUtU1jea6YWVYSWi7URgxT6JeVPwPoEqp6vkaEeuYpipUVZp/bTlOYcUbDV8/tIJdr
w+Fzp0wMBDkWih3rXNU+XYYlbcQgFRuNlJkpBLNlgh663fUIE33pLaW6CmEoiqHaNRiXrM4+690K
DBKIh8TxIBwJ2fOdINYqPA+TcP3ftetWPNOGJhu5KUGR38gIZN0hUZ4e5dJ4Tf7bDcxnB7qE7itC
nr6HknSw+DOKpFbiTeoVWenWORwt2E/NRxd7DtAdBGVIxmb+KGD05qTv8+nY1cMUUJP8DDxeR+Pu
5+66fpRsOwmAkPSJVMR5JUejkBmavYPLX02fKFUWW4C1SImGE+ytysVkAZ8I6xusppgsPb6pEkxI
6/2evVCJ4IUsHILkSQqBCIlhw+ip1+FyqfOY7xAIEho5DsAhi1ZK87igLUSX7z5agLdUQzhriERX
9hs7kzjPzdZ9Hx2sHLOBYqY1uO3zjzk37uV3/wsyYolRIosAfG//1c5DqZkBsWCLsjJB1SmpzLeF
fjmRMBoX3SQx9I5Y8NnXsmSJWWQVe31RtnTTna0z89XfAwnvV/8sDTB/d6/q+H41HQy5zCYC5DCs
sG6i1+i1pDDN2kd3sqZQSYm28C9XtvXrJ7UudlpqxJ0xxqk5bGSbOecOZZTC7bavEu+eMeJC8KeG
QqI0vAz37cHL74loCwnHIqbfLa7FLIPAOiAHykAw5VbSUhAMZZdxsizjNkaTprUlExk00o3AN5KE
uTc/HgHaNaTkZsAShtglqaZ45vJoIHnLh7tG7vtX6IQL5Y4pyjdlnVRLmobjwrXSscnY/szeA8xA
t3qfacWSFA4fObqtoV+3mxu30F9fbHbPzW593TS++W/mRocxpKyFoRdu2ZZOWyzJ1LFcvCD8RQ1D
Q7+CQiMEq6Wl8n4rK1f9sABVBslAMEr8dFbXz28y0X+I95ZOe7DuFkzHyPk4p6AcAhgvT0Flix/D
fq1UyviypjV2A1sUvzIiEasdgryU1PgRhCJWMD7jPW4we1sRCXFws992DgebNtYxMGWF4pGQ/yRE
PuLfs3xVX1IPnWYZd14kAf7u93Fhc0LNitYcRtyfrD7DuSYQ/3KVuEg3JuC3VdQEkhNB1SL1ONKl
gzV/O8vSuiOM2LdAaEEV+Lz7gxyOe2pfXidHeUR1QYi1q4WGNDNEPGRohDib/b/J1A86fkYbBrE8
JQwstbrJ4kTjaUrG/zwY4xwjtBni+Fg1nYfnZjvt1gO/S/z7FsR9zPoxP2Mwx6uxHFTP6DBAfMLr
XH1xSfJjsBaHAIhUIZAkE8e1IGQPFnPO+x6ERzS+/YCS11ETm/0MQpJwpWuTNbut9pIWzecKAPdg
fUvvQzWh4rZDq1uqthy/IMFLoRKctiYCB/Io3qIWj8WbsSk9EojncOCTT3a6MH/1Pt6OjEorxC5+
AnbEs1AEkhZq50dyt7Qkx5/J5lPWZ6uc5cn04y99k30EjvmKhwF/7tApGW/sy8ehVsSoNURzTHFq
jvo8jSO4eZ+ZGUIEZZqCh+JXW9I44EuZb8EkYh+8bCpjfmqs/Li/fkbOm5mGluow7WbW/dA7/tiw
7y2GQJPbOob/pJS3RKf13WXEJcRKuNJJfSbiK7K2Shtc8GFE42F1VEYDc5v50krJUmvRnpIpHPJo
CY7goOw3tleP4BAzMW60+JCtVxMinn1nmzfOsvwtKfrJ5THU8ulRt5FRYVbpJNU4Xb0Gp4gIGTzI
uUQ66dfr2+HosTepLxdiYsarHEo0Xke8T3Av4DrxMPmHD7nnJZiJYIyoHKjzBQIQGgCx5S4GjLjY
FA9FQKm7xN++nfbOQwhRP+2do4s0ryzQoVOZMOoKVAI+W7D2DYCtV+DC5vP4wtwb+cKlr9ykMmmA
5poJI0l+PpOFCu04+Eu5PkaZn5UU7Bs7906pNbbbwUpr42PXfWGoz+KszSv922HiKDq0meFAXrrX
Zkmhq2ta+830y8dzyy1eRb0LRVWS/s+2CknuTvNYgQqO20Y2/V76/chTYmo912bLNuqWQoGkEt94
px16pkw7bIEIQ8YkUqSeIZgP2rpyLt860eD5i7Z/35a9NoPHR5CLDbMeggHSUUa6IWU6TQSHdB4b
eNZEmOq4J5+HFZraKdBKxkihkcEhjqkBxYfIOXPBDnyTDkER5ZNKZ4Qh+2BjK+tQ04Hm0oPl0t+J
0IPcF/Cup8Go0uELDrmjhnFfD6qu1+0BFU22u453AQJknYcAkqZ7KRxXqcIYcM9uR1xMY3DsxTfo
Gh5drEuUgnZ2Wmh4iQKO3CPtpC1oZCdrwDPtE2nukNDz1n+iGxDKP7Qr5MWae2LunqEBwTNw6QCl
B0BXKgKGA+FDYnwxNQGi0OaIikPcN4+EgstB4ObJyVagKKojrokFkkqpZxp1yfKVrApfd+J1oeCh
N+UYf+mdgf9KtUh0kunaCaCnRXRU5FqEYZdu8BnacIa14xLBYLR0+i4Bu34h+6qrQd5r1e50lR3O
hZji0N03qUITvo6ZZbwDWBPhV70GYu0QLjGBFyr95sEHm+Btl4VbnWiAYJGDAAy6f0DweaEUm5eY
li7A7jrHdZ2rnbPFWuErpCEVhYihKYBB+VxyUdaqGmES8RlXaAn9iKdP29z9Kh0RbMaDvntrtsuo
xigSospiJTrFF1K0Ns9KGf2tenz2U0OAxC4zE/ODqQfdmhfLzOs1Gtaz0T0C7MhcjoZyzyuICi0b
vRLpwwb4KHQtiOTu11MoZr2wf0CfSFxx1cULuY29z0bTsVGvYb9j1T97+EtYbCcVUgBDoPSNND7J
UDGKoVtta5Cos8SIfQgWndgMU+7UVPKVnj2MI30i06ke5mqp8s9X3sYXcVfLWmEf7EeSPgZgAdc6
DfgaVmCK2F1cok1Od8/c78eBy1FcOzaIDotHLmjN1vyxyXBc3vi/1NqloX2kZgpCFxNHGEUeWRnd
ubVQk8V/cPq8WAVJ6I5d9xywWw8/Bo8GtSurdhBiGOS8DlzuY9iOth9+k5vstcocPigSPvtyrkMA
LeEGdLPxe5Ju6TtV9SH8WpeNA/oxA3fiLmYKrCFhTrN6sgtUiXrqpf0B3uZ4OelrmA9tVjmGkYLg
WFPD42NjqkzV6dYyzO5hdUZEFtkV+RSsJ76tuAQcrBAkQT0WBohom3c1REMx04fOdupE5rQxBqn4
T5yV81HByPrZUMHQqZWijtmZKA8ocOPv1Q8i8auNNvpsUw8775odsL8bUGE9H/2VfxCb8gWqreU8
luQCOsEWLFHxF1qmvo76e6wyNuG2bIXd5JDmjYBNl/+xFK7yXH7TRS6EuUqjGfEf07C55xqdLUjN
zysFjFE8QTvRU6qfIkCUuGuh3qP4EKrgLatLNMBh4TmYm8BSXhH9jo9bTzyF2F05GurnxWJI39og
L+fLyyv2IVF8xr+b1omzD3SUBpOm4wXB6S4jCF6XeSbPvV6ui7MrgWCDOW2B3IA6jbMDlnoVNxV9
Ik5NCAgM1fWTxKURFNadne3g3MF19sc8e+EHQjd0KITukL1cs9j0GoAPLbSNLTpQ61+HLBL/e6lZ
FfVZ/fFbLDbE/eKeaAagsHklwARnGccngxzyECqivJWfAk5EWi2hSwwYsyOEXJtewyYuGybzgqyO
cgLn98Qd8icPGvEaNejixLxSV3ZmBbNPxHzadAyD2zLcyUqNU9mR77RxEuK/L4mdnD2Sqoy8MmWK
44nU+phK1jpSYVUAjhAEOuDihX+F+KfMDGNkvCqmJp5GeLcFmFxSzzVvaRw14cCkvHvJf88QdXLD
igTC/dIZFu5oqbDhJRHqSuJoYJWh0VxlSexM75wn9TSzBSjLimApEcpEJIJ2lCfuhLxxYUcNRtyM
NKG6vM+CdC/+YEb1tpRBMSNGEcwDVMa4uLuaV9WSZgt9o8d3kioEPYici215DNxYdWSbrhH31pNJ
ErTejViSE3wJoUQ3Rb22AhvONQsx5Of3H9zKpmIsD+UdhQ0Crz20N2TbRrXQNzaus2HpXHbhDsLv
D/rkuZ/4xZ9KDBID7RIkcSBEMBViQf0f9xN98i+FymY+c3YObe0B/HPPud+RZcsa9Mpo4yQ/XI0F
muAl0WrnC9w4GRWVzm3v4uI4+PKBQGjXfu73+o54n07jMQI6KcuREzKQAMeRQQNSAXdfis6tJQYX
nHx6Kkb0qkdyDMKCvOqcvJZCHdjaL663y0RAz4mn3U1dzoN+7CshEmOyBlFvy76pldcsMPIKq2ny
V9m6xY1/Mv4f1s1hnmWd7EhrBlcw0IR+mCMTsYK4uvwEO5DS8H7gyOYScrhBntvUbzzDeGF6usOc
uA3jVAHa5OqUSeaR0uyT1ING/2q8ajoho7h2btCWD+y1Oh5EcW229t8aI1VY6Bz0/x0PlQtZnQAl
9qLTxZZUmcDCRtg+UzHl050+WTnBkCwCooXN2lLLZIlQhAPJSbrZ1kfa6k0UjJMoD+ep5777g2uC
nftU41ecemXJ8aZqTg0/n+sBZ0h+WkTrUs+wkGlMLl7gjtZNcfpvPrUIiA3H1lcCFJMFvOHvR+Cq
19EIS4PYQXIxg6FgIvSm6SJgiFWSVMAeMkJgNKQy55ZpdTAfAekhYOEHWvNE7vKWGVYAT4tSfLSZ
COrN7C1fKOKDw7Xhj174dWjVsmz7hkMmQHw7qWDkJpnkWfoTPyIdHVjkhHlGO4zzat/8B4tUqv8r
kN9ctet/5+ivXRCEwWk13CudlsTz/wdTZHPwIOxzqQExMfBrvKEs310C5H2Yv4cR0g7/5OtX7B6B
3YRG3lQLv15fEdbyY/Hv38x+U+RB+6Sp8OHR+3yK3bF8CMvMk+7zrpKW7Pdwc3alCC4KBTnlz7ll
QmZynGTRF2ijV0s8P3EDWpA5VpoywnhW3Y9J0ShTo6MX8MjpBfU0nmvTdvHqoO97WF4on9STI9No
Vg78ZSMoRVI3ZAjb3jwvOzpAKgQo9ZBo8egoNERxPVkYLrmWAOsuRfSQVWlANj30qRh3swSKgKru
ISIM9DgstPfxkcaVMwbcAYPfZKqlGAX4PtpMKdap9BTn8SJ1WWRgIn2JSf5WcKt9o1nJ1Q3F2sjy
G/MoA+g5ZwWKUlBuginBMhFw7DWeRpmhdlkoSVr1Xn7ssMmgdoN6c46EdDlsTWoFlF1mHUhi/LTd
wXLSwQUxZeQ+g1mmRJuaZ2KoB40ZbrdwJKKCcIEqQ8M+3xy7oT049jYvfY3biTcyRVqp2ZKgKmiO
gg88EUZgcprBgvqrC5CSF3dhw4//A0NsbJJCsHfJDBfon9O677u5/JWfMPlQPYiSR/Vj54CKmvlC
E0rRWZohqntnPFGTcmREMhFdneGXglDIObdtNwpdAN6g4uX/LHok9RUDNWJWOFiM7X5pQRcCMrt1
74l//FXanOJV4lidSpwqm5paKyLU98bp12KFjcp4QKbItc0wXjsT7/z9w/8HqIvPYkqp/ZO0/2M7
SoPloraA30bNH5rKHjSdAAoRHYJCdGBMbbHM4STQVG/nETG6XVpPpsoGJfaC72VZyDNvMCupHonx
1YEmCmPl93R9BoyjfTnrVXClp2ASuJny4WKRb5wyHixkT02kh0xbF8Zqog599+Geg5u+kmkSJyz0
MAHfVfrxov0odsL+wkJXusbsSz+rbGCqsl2w/3vb4T/d7CY59xPqjJQQNLkP2OVToncvK1UkpT/i
PXM6jXnvdjzeN34DqTSSKt1Mt0jItmbywARONRYeBRLTHgiJlRZq4kWCZeBk0OoUAGjWmfvBcIix
NBiSe+tL8j1rs/IeJpgWca4X1Kb9InEMmkeZ2kQ7QUUpnlPk+0xsppwb9RnpDyydlBVfhWIN8hp3
VjkmgoBjAx6BCAv3AyGtQ8pbJMtEAFb84tcUG0r5UVks8lCf7uFGnYw5cXfRbNmV/t3rodoqkFRa
/qaeY24JQjlGAqtfO3FPAUmr75rqVyDH5/WjcQMikCuYK1gZX2xjwjdgLDasqwgNU+WeyN3iH81N
MlkS/OBRgpt4naKy5hc6kCRuOJ88DeuvqfYCqsdb2UqFE4MdUBNPLqB8Hsu8aifwltarax9icym/
IXPdeSHfNxJPySOMLE82SYM38jsV5xqIPLPSUb/HwnycI98bDP4kQB4ULy4ruXlytOu9IxoIGg8m
9zJnzcq4cwLNY5WIKNof1Fr3tPLdEKPhNDYcCrA0qIVZm5266xx7NRojgVdFWhnI1vN52qpIF/PN
vzcoTfKKXOE7Y2NFHq2yflX0LHb+l8bTa2eXdQilkrVC0bor8EwFPD7Y+346RbL8mAcm4ekbkAgL
8vBhHq4lcCr4G5nRNDj02WPcjb7YgjtjUBPVT0De0POOpZhW7IylnbPgbcKZqtMm1H6Svch50YS7
J3PClVy+9e2XvIzejZ+YpGBigrCj/O3bzsai2ccBBm71jpZWTvehTBioi0vkgYGkjRBRtu7sGMAp
jPGfahiBaOq8hTzlkwKK3JmjTv7bYDrQYPnvGXMf9ebXhqhegMXywRwj9uU9/Lq94OteNDGvupvX
tA44WyBNGRbbYShJ7XroM5UxyywFGCuhL2ooBrXGD9S1Kix4VN4ceA/CQrt6OGTNq5TSWd2yioIr
2kXwUMobLntKqTcssNLCeyatIG5k2lsYlxZSYn5VgSNJfvxLL+WU0ZNDCojh5uTVRVOZPq2UO0Bi
EmqbRs1yl4OOA38ng4bp0atO6NozT1rezZ31kTvDeWr96GefmdKqxRpjqQaHBsdFTd7/WRKhDARG
kcjkbokTu4ZIGIv4ZYoy/SmJiMEOUlTUuqI1w0pgjLKVAPmfyxLBot+lo4xUStlUl29UmDlwNDK1
SwMp/W4yN/0NfvrqQbKszUtryWFYFh/1MhiCZ7kPtwPA2OF3whvI496mrzNJO+djd/dmBfZuXMlT
Wez2Wf8RMMhdcGSaes0PJgGnFtAP9fLN7SoX8mbH4xhh64VZS3esVu3tBjDnRDtS+1Hg1uPuxaX/
H1ZFg0HrCe3IFisDGa8+VWj55HuzCJjSiedEocX8AoAAQod7QW7kWbDbkNFINUMa74/q75D+VkN6
ldgDtt6T7C87AA8qmNPIlohjfdFRK/1Gi88JDBFuQOqrCQ6fHp+gZXjN9THmsDfFszvjJonjpH6n
Do2WOk8wpwHas+ixWnrbwCTr6ET0f8wGIQZqvKIkGBSJ4hljlHziuNvYbc6vH9ERxmPVJ3PMB9id
ouoiAd4fNPtK5vK6rOeeHIJzH/pl7Q77VQGhoPrvKE+xCYS9+nV6uaP7cTF3kyl1XnIZbrkFYzi3
V+P4ZuE1stuI4gEntAHOBoYtTVeVpYyedoJzhNDxZenEYHAXKFin8H5uvoIg8PKOgwibLUArKEPU
ln6dpWACzbvnYXyIPa6cXuM8aFIgCOgeJ1K4m0GMqMmILZ8aqwJaIlfbsIS7Ibdq2EF07qYgaEx+
idK7BvWKhxrqTxs6VJvEgkz/5wKKsEhiBnEE2h60ImaP/Z29AjVeptkzRc2A9lqRwa0UqSWiCVLd
/op/u4WIdYTleoxG7XB4lPzp7u4wK5ryGzvWIrJGH7j+aTo1ZV0oCunLdl0cRjklCTYmid4i+ieN
toDCrZN7YcVLEejJCaGa5rBTXfGEd7LiBXHgsFonV+rgVTdqHYb0zOW8F14+rPekS2dqGCcf7dd4
2Vy1jVHBCSzoNLRcV+t8EDhLcscSlFFLUIiH5OMr+pZD5V7wozTOhXQzraEwr9zV4oQFdhi03CF3
lJqvTX/Fjg42G14yvbU6gKoWLwcbpgu3FgDd36FhChGbsnKs9gTKiPFy/MNuoqYmUGMt8NoVDb6w
lQWNA0Vd8aZxkay3JooafA71q/hwPjejjCENpAEhagcmY0CrEYhubFG2B8frXgYKb2bngzVu4mzL
rVPq3Ws9Dze1xpAGgMmjrwzodGVomDBYLgsWRNBoP3IsoSpqmN1mTc3qqd8XU1tGCvfO/mr5/E84
LNHELe8r++zIGyBLcAx54DFTzn/iUrMqAinl9MoxiQayydP+NzVisqKNN+dwft6lhzyr7qvIXvWS
9pQM5t9JsSoKRRb16ja7oDhPklW58EX8fVHrQL3Onnakor8c0XMwI9Fy2CaXFfjh1lDNdmII1Ib4
oDSGH9KnwMgT8qPlt501uC5Uw2Y4lI8utEW3tjRnmM9ZDCHGtlxK2AU6gx723MasETz88k6ROJBo
P47PkJE/Bznz+GsUe95AB5oeEbKr7ml4Km1D1e/YDTK0vCU1sSLCkdhcoIk1Yiq0unUKACAIrI9Y
Aiue/ez3HssEmG3dhe3WEo6oVh5tsAhxEAwN+UhSugUbruOBkdPrLOHjN4QxitT2cEP0yhTvsPM+
RuqnVbYB+eN6hiyZ8xSY8mZD910MFS9XX8bJCYdaMXQ+iMIoWEc6NLFzukj2szdfckixPwRa0OO2
P4/qROx3De0WM8SCvQ8Qrchc+EkgGm2w/w1YiqwPA2EhTh3RtbjaryNDsiDyx5icEJKHnrRSmuWc
ghfoL9x+EQKy0ZLlZtXt7uXcIXc36Ec0bSkgPTgo/jbqfNMf4ZLlMAHzHVeYT6BPdy814MV2+nqI
qb7bJA/jyQQ/T66fZ7JlH87K9OHS0CycTXHLuSDRIHQRBKXg7WH5ewNxa6mg81ovNrrFrxDa+BMN
z8ydV7XBf3E2BrPC+L+LnTVfewYbOE2gZj88pIJEjGDCkb7075ju0zDZMMHxCusQainI/hBkM+36
eXuQJgnN1pOqxPZMrDibHmpld/8gUdnYxJ+EQfBM/VmM6TOl7aZvdbw8fYAQdg4OEn27Pd1+HQxQ
GZM3vOzOafi7L3HLRhxiS228ChlNyXqjqNX4Z/7tceIQmkLDUdv2HcBBkDboYLzmZYPlGNUBFE1V
hXWU7gMLVxrvcJHPvsfXuB2IsVWfIa3UvZv5bsBls8aIkZh+6dFd2ykY1cPicy9g2MGhkAZuGaAo
NuIK7Y9DeJTVL9r3BOqwc80WJUhvtbt0mBQYaIUKERyLrHhSUoHdkY5ODdTtRsroebNbNV1Whc4M
6qcg7UxsWrYkKxzoQT8gSn0baeV8G8Uh/BTBtqeGSY7eHE3oZ36oqBOS6VLC6mUa4V1yv9NIcn2Z
3Fim9Dle/lA4/jPb28XXaZ8JftE5D114skB3BL9LCeIUVyDpYqkKt+26Xj68KhT5l0Odiyn9qvjh
PyM1MHKoLoBomwlCV6LbHObVDem/uLXxQVav5z8dcl1wcCp5UdqzXMBX0HpBYpDR6H93MvN/jWFE
yrYK5AmDMaJFZb7jeVOu0L8TtNj9xlElsYNEnpCGizF6HMYQBu2hxzIbFbEVxThfMBVeauTW2kVp
uf5gd3jPfLnm/AIG5mNTNe9FLzJ7BWUcREDk7opJwGq4a/2FqvpB9vPMKlku9zc0VNUN515naOYv
+SJFVfcBvq4HVO/LR/aGBc/kiif7f1RekpRMhjEWUI8quvA5oJB92AWiemyAtsLzH/EuYQrRsmnA
7oCt6MzX2sgZNioQPzKnvnzxHi0dOvHE0cs8qde0zVcT8sy9p9jRBl0Q7BW1ZrFNA1wqPqvR0kbW
VpoRLt2CdWy15lGyD7lOqz+SilMF9bKHVZ8p6TQLxMZXk3Ou/iCrHjdeA5Q/+kCzFfCTgTgAvT4d
tlLYIrce8Gu8haKYnni5ILYL54GvHcbq09a3iuhJczAE51MkHW5S6+kawDb0rE+5Ng+ovcprPpTm
3Mb47rVpZx9ZiLZ9nPXPD4q7UabmSIRFUya7kVoZKM/zgrIxVUgxzkpqGR27ytNVmAkNcio1c+EP
EMwxgKUoAJjIBi5QHMk+T2LRswy85DBS/SvoQLwx1Qv4bvRKfFc/s/24zt/eFzqku5LatWDFmAPn
TAKqs2vGCsBOCy7v6VqDridK2LwBeP/OynrUhUvxRMM2Qg0paWzprRXDMCCiCSOJWuzqMA/MIpjV
Lks3SgTp6IAIakIyUPGmA2PD49s/uvpr5jfEGwmeGbXRgOdgXO5rFK2gBMwsrprXrb4C5Xsz+ls+
1sceOA8lel2rXl7Tazlz6og6cFBOo4jjPuesDY0B8wnfOE+oKz9JPey/afq2Fr0FlI0U5DjypXy1
p2v61hZgHeHIuiOBNUt6I/nNUWaA154J2jprBKMVbK+NiUKaOnZH456UoLVIxliJ/EY0HskruC44
tnxxXazt8KajXR3lun7kWB7XEVJWcNsweABU2JPZXBFvQIq0p5FsLXja993SXiSJb3YA2dhkjzhJ
IVjh74sZTadsEsZocWT9RL9AcV+yJglHV3RYfhk1cHFIehQ76WhSieZsr11wDOktkV9t4tYR66xn
kDsSj/d9khC8agxMs+vjsU8PUR1aS+QjUcngemGxHRn6mGNdtJk4dpMTu4U+pwDVQQu/383Y2dDs
TfvgPe/Rvu1/7jIju9o61mppkt4WW4y5DcJx87VL7WcNbamzO7/9c5OwwLrBNnR6bVFnVzv1d4su
YNV7D0voD3pwT3m5iqbFdZpjE2RbPF3piHhpceo5n/JBmkDnk/B5iOT8938zggTw8RVOztZLlsMF
0j+zP6Xmk3d7ogpmKuCLFOmu0VVIjGAnvT2BVLxSPQC21s9nFobeiAryVOoWwMchAWwFn+pY1ows
ILG/s5/PJdiBRZFghyQEEeHEU7Hk1TJXQHbMcDeNYyqCSqNsrJzQzt1EwCBkF43HWX+HIWgjVmEO
H1+GA9n8+jhdenipFJ6BcFFXFz5PcWcN5LA592MVupr+7Qv+RWmmzr0V0WXowEys0btAT39oHgTX
xrdgNrNyiZQ8cZBA+4zUdCKxxHGxYSrqbS8Qyld8ogaiIk/vYswE4OTFKSKdHWoSx9UwX7glJZ8A
b/MmTECtz+fMsGF1BmvrT1mg9d5LklE1twxarXO5H58xQeeneD2O4fudPFLjBaegX6AMNMj5yupx
ByXj3A9Ty1Yx08574eCoqB3tgHKP3fInkFZV9REq+Eu/8WXj6FAX855OzVmnDkbA16BVpq4Oat8n
dghXygKkRZi4NwYTEdcPncatW3vrQKkSmmAZDmG/iPCIODpOJVQjABJ41803pQ4r8SZfRy14ve4Q
3y+gcVpb9KRA1tiEPzwJ+eZKtMK/Tkm5NfTYhIjeTIOjllrW4vUjf2EG5a7qYJuBK0N7ZYvitGbe
s0nUEVpjy2Sbs8p50kjGh90ytce7TmEMd9v7SR9u8684orpR0/sCUIqhsbVkmcZWOdDj/zYx+EDS
Jc8t7wPez6KrTSHOtR8o1v5qqLqOY3cHyy3pXpS9HsQdi0k78jhvHEJmCjG2Bn4RNIktk4uAlo6R
UJebY9An9+lBDGw2yZpOjly3BU+p4AKJJdgZh3rC055S51Ejhs1y6UYH/84FVGoSqWb1dzwpDKg1
oQMRObthpAv/n4BzFd1WeI+eDovVz9prH7M2wu6h/S3cuvvfvj4NJD7Pc1tJ6uMlaJwChgVTEexi
kAdzhWZT6/fDKhgf/gGF3cYS2MJEvmY4jwC9Kdj/pRHXQ/BaH5VM8+6u7fduonEh9BquxJogET+c
oy101cD2ExgNPg8Zkgwy5z9YVEnul01LQw42zCL3zaycqxA3d1RMv5bslBy8MY1p3IkY9XSbq5D/
6492yxTZ0w3rArQCza0F9ca9AnmMcytbLYrsL7W0qKX/DHHq2bvm5cMiVsHvBtSW86gbzYqebjXz
vPFDjayKpLh1i1YKxM5ptkm79rqvndJYFQJY8pQLi0kV+pE1rvub+i3nVRbbmZMMnHkIbeun5AmW
6LELXz+IdBEDkoUCTgoJVm5z+AXOIcFYP38IGoPAACqjFvP+1HVKnCPl/HIdNlLUTN8zlhVxSDn8
FTd1NUwpRLIMtfVp7s1JfOoulbfSPPiVYA6+3/rUbSoLagyvA6y9A5LrwsJut+5efNZKGFtinQ31
VD6oDDuZSkFuzC8D8x80dwhdR2lLUibEO1qh7Mt81eA/jgfm8E0As71PeSzNQ7IAVe/++i+qHfA7
R7zcEYIfyISKxuSxNJH7ZAugjWdy9/InvazkPrCOzjAhpJhV1gchpmtDDnTLAc7dthQtlQEkbCf1
t8g/z3d0yzeK3YlEbkMu2sWFTwxJtYYTX3759ZFqWCTNSu11iOHspCe0SHwCKOnW8HTooAarajCd
pgMZpyqz4xxcP3xdTtaJJK9wvwA36ohDzlrmu5reT6XmDT2LIxjGa25bcMluUCoP0vXADQYpNSUJ
YFMfTb7jOhtbqnJRgpCuRijrU3lBXGnI1gpARViW0FMEwh2i4YYguBKiLVAkz7CV4lLN5LDFTOd9
ySNTCMYRrKlu1xqk7CchC9KRVntsU8nN4cktfFjYpIRE+2MmJClQY/S+zGxx/ONZ+JKhZ4BxtXWy
n2ONlwf6AIQC4qlxTsGeId50K04y8c+hXSn/viBa66prhZZsR7JqZe+aPZnpm0sjfZ9d7A+zOMte
4S9TvzuKjXQzdnj7dlitN4NvGOUBwuW2C3t9xabjuyxkbMc0uxxLKJXsbikXJLv5iXpqVF1VoSI0
1pwO5M0pBWqwuGMoe1j+hsxkskh07WVXkvU7pO5lOZF76t53+Ud+YPWAk7XzPFVvdRm42fzkacgx
H2ZInNnWfyofDG4bet1VPyCgKV2KtFRQCXI0IbBoHbAYRbXgirqewknsEmV6L3Wqmsl+LqsKcHGt
Qs6FVDdalBxk9fLB5I9SpWbwE8iU8Pw70AlM/ltJs/qYB00PcoulkX76AACtTexBZEYC4nMyo6ib
JOoTl8lNqfDxIVdEv52EqtFtpEG/djKl2Mk/jaerxcbMWCQZ62lxhfPINi8paVeZHEWWoys8YkxP
KxVi8dxWimVUT9l6MyhJXiOZLd/z3KSAUW9g1IHQ4kFzQnl5iEbQms2D2s7v3X4pvptgnM84VF/t
qeB4xdeaV34lnumuPIFGCQPS+11WGe7obRo5Jt47sQvOfKgndqQGZ/3uOHc8LDggYahacpKBalRO
/jMExc1+hm77c7eYd2FPGF/CovFgCjucFdp2egRaCUGktp/b5nZNV+0GGwXOmNV/6GGh6KPmP9dD
+kXYU5hxQi0YRSVT/xTiyEkcU4vaXE/pQhOlYFpbLFKS94sbdSZL0PmBxSuDzCWJz8LanTpkVFqx
XariVebf+mYSwDbquKVd2JqhUMgtESyaB7c6MsihqHQc1IVKmvLg6W+2TGw9iGEjgI4HAg+csa+X
LEtkj85oouekcyq2hQZdjl08jdzlakgLcbRGiMhnMPYT45WAjLkYBbURbaA8wFA9txZkZTwj6/q6
XytNf2vCoiW4FE5sYIyu9eFs5F0q9wTv25/+zQbBqQRwosWvbe344Xst6/n5KGLRuDz83P9wbTXO
Ub2fX4Y7NveuumonYR4S6O6A2gghs/REv+0ektl9YLn+2Lmfsmqn2CwW05lNQQIE6FQvOaj1Iybx
Fvc3yf5JdTWrQsWeDx2XAaChLeTgdmBj4ka88JmC4cFBk2SJO6c6HSH8ysoMNvyiUeVnn79C/zjB
DrIc9cZ5nbi6+99JeqyDRSPOthQxAjIVf5R9C9L7PduVp+8mlpWOwjjsbryIORj+sBBQLShfwXwg
9UZ0cCsfY87shvTJ49QDwfE+Uq170IQ1kjRBOuXv7ShsQSdVMiAghs/8qQFtjTwMJrjJAhiudB6/
HiH/HvbSg0tlOOAXJlubyR3n4jAwg6lkio6ZvA6HczQL0tDK/mLSDkb5t19/hyqnbGSSDNJ8l9vV
4Wy5XjvEnGIQ8C82TtFBLm2tuB1TLSA31e7n0u2txPGDBrX9Sb3v+Yq8k1J/HWqpozdTaIhp8tm+
xk7FjAuJ/GQfZbocgK9+9QUWP0HfEO6GgF41hCZWGZFEL+ptBtu0Jl5HqTwE8tyrHwg0Jr5qbxDn
DbBM1PUMHiXsdJTeSGbXTf/uhAAA+DB9gel+vlb+MOn5uahb4r/lDP89oCVN2VrSiDFRB9v0O0te
0BX/KXXE+exDjWFYtXx4Isqqaoadp+Htdpdeui5yto8n227ip6YC7SuvRqwjlmBrorbKW3NssYas
IPGrTBrTzL3AavJoUPE4CwkbDvVIyhJiU2OhIEcCXR+Spyk2vTRHNwMLEc3UThiv3gNOujfv7uOF
alvn8LJjt+jeKZOFOr/+rHuFCdAdKANoUZ+C15wccEb4eBTxbBWMfmAT3nRafGR4NkqIELMYpy58
CZQ/t/YgY7zkqgRuQA/+OWakWxoQF0PLUMnR+l+z18ZgWR9urimu3pVLaDhEiQ1SYHZHd3sJhJXI
aamBSOIj+ou50EqL1XiwnU/2vYnygRHhTAaQAgp+PFMK2bDgG89QP6HDBZabKZOz0dshTfwHZbUw
d0UGGD87Jln3WXB1UjmcBHi+XoNBNCql5geeGkAVCC4D2G5lVh0GV2E8oGJMY+wJErFK4QbGa95t
7W066U26LWCnahEss9lBMZ4AmOGTERbIuokwcERx+nZuW4to8yhG8fbcY0tRSSbihU28Riv1v3OP
91JIfszZHjMcyDFrN6LPAtJ4D8jE2U8kEB0I+kIb/1a84TKGsgFMh0S0V2kC/+YVgYRu/sJGmkRS
FKtuvkGv5vKQCVzxrgW168Ljs3OVoZvzbA7duXlssiTLLLmRWAHgak0kvMDYyDxxGDgArd2u+gkG
M9B7XtClKTrZiZVsWHuN3GXjcPaY9jDfyxAPav8HbtdHgzp9cdyanomC50n1PTViNwec139LflB5
bA/+0MaxVl01DXE2XtL1XQqogbSVTi87AxknHZpxfKfQuU3CgP3DpSu+i3ziUBSxDNOKZCNvtB1p
/YEoOjkJ2bv3+P1xRVrpHCgEAz5659t0mHFSluDDfxKvuR/RrOVf+lshm6BvGCSAY5bXZgolh8I1
iZnqefRwXvo4tx5pjiTEtfa7BJKkzq2XXHp6Ll6OtVXI2P3EhDAHHglNHFXcM2phvGzabzN7oRCr
I9QHsELhZUyuiGPK6ho3BNptmGVvl2nRva58drF7qZeNfkrOf7JtTXM72XUiG+gxYxU6egoESun2
7aswgdMjkQZVaJVY5sxZ0JTs306rYv1MCPgoFXMW6MUa10uAkhmDmAZNU0JQDnICQ/iWTAH7NHN3
V5T5fGEXayQGBYrq/lXf859tCvq5ex16/fZrMY8P9G0xdtuBhUh2H/YNQu6AweT3kYr14ypv1WPT
xa4AR01l/tlZMlbyvKs5+/koC5uznytaYh/DGlbH6ZPQdgnbIERYOcCUuSpKcW8F7qCox1/XU380
cVabNyYRUBqK3tpjEXrhKWSPsTBufJ7mKlYPbGqws0rFq53EXalNU13QJXmEJJr+j9Udo38jHD4u
qSy7qc5RwVMmJDxNrG+STFo4RcQ2w3+4sfwSe+AJoONzopezNEpew180AwLVYI4xhfSQr4FaBCGp
jrmdg0jjHPSZOuItYQPEtWDlQYF3FUeeD+aNc3QDAgUxVrrqilDEZ1Rs9NjbYshDawz6lI70PAt4
cwvqbMyh1CeUfOh7E+EtKoje4VI+qJjmXkLLhlD0ZDMbgrp91D5Q9kLtzcDuyqkAgb+PfV/noNxA
9Z5KcKTwbGwI6BLOOt9s8CKo1nDr3FxibXxntoM0R6AEDOQGPWt7QG8jQ01jbFWEMyX6RL91bfXs
u5TSrZ8W+ca0n9USQiZIPBwXkwsQFfYybibcqIC+Kk5/PNqae7m17Lr3dxy/a45/PmRf9frWHjVC
2//YDYYpSUigRDIswY8PHRAaUHXJTJA8H3NUeRYY8ltQmDTTvYGp2qRAx2h6ZbSaP33ei+wZ2IcB
j15n4l7ix+Kg45Q7sg8PPz/9BG4UmpftlXmvWUNDvvpXbHTXWXZMLRpsmBFsiR0g4InQ1sxDEwrS
SKHKb/Cs73fb//rsMxTEanZW73BQzYVLfBpczHj+6wbneHnGP2v2XKwI0SxFShSP/2ZcCPAFLc0d
hGQVlsI75uzkTOvzR+wCUMhWfwdGR6f5yVRukgAR7Li7PKJk5zsxb2M8Jz3ARg0cdYosp+IOE2UY
Z5PSGAA3CrONDU0gZMGCAGVhbv+FP3tSTTEbMBLUnyxsT4Jai7DrS4nNqoRX8h3wqPC04i9OZJYh
qC8D9CJzfqot1Qs4jueMHESCTyoVUgCDuV6/nWgaGNaSqQWyuvmfIaxWTNq7gbPqy29kjGAKZqGe
1ROYfDEiDFmQ5+KzM2V1eNWxAQf3q3oRAZQ3p3/KrEZKntSvPz5c12b86L/RvfUX7UoTpWVGF+Gg
OpkSRfwGwEgF8zV7/KFL9Ra1G0xchY6FDnDKB0dBFokSG9QWtLBsg7hWL3DXM1kLZ8i6mcjGNJT5
FwG7nC1ycak/wicQ6k3fXE9ovfwkXglXwlpUAPNpFyzVu/BSZaxlVIGHUHftuGOJRyXIYhSg12DS
IoK2dNmU+Nz0wTpWZGW3Q/klQ7EMsLEGLqrutGc0tl0WUu9F+EaQhDjSKA+norhH3B5uycDDFt6g
amX2RSEHF094nRGuOY84xME6DLoqh3gB1a7X8DFOIo3xJiZIITanGhCyZFlOreXbpjA7KjHGlTYT
lx09fwT68r8c882a34c3HeBtRvm1zmwo4XYvwbufCRBg2LZKRFv5GX0yQejnul0R/CVsNqL/pRpW
QU/YDsv7s5+aN1HVgPEfhL4miDDLHevBhPhGwDW8AC6hSSOp278Zg7G7GpDgmA5As8E97ITdoMWL
8vZWl1OaJZHmMFfuWZ9hgGBiJHniLOLs5yyPb63miWaViTCtKHKtZukan2zr9ID1wlnHT6MMQyd2
ygU1tRYDh8DlzFSKx2zQqAg7aR16VKtqnoLdf2/vP0SuQeH+ifWqzrzPCAxWMq85tfNLpEezaQpl
06N33i6zbVlqh9F9Pvqu3fvgwRsIAwJC57JUo1/gD3JVtUyXxVD10D2HqZ7/thyUk+rjgFpQylot
6dGOOcOKlbHzgIBt4wjRfBET2zdO7IltTMC28uUiAvD996vVm59GRa0HBcTaXt1PNhcYD5/1MAYl
5b2VvkbR4aOUuTR6Xet5GfdokJOaYDgI9UjcQWYfA1j25bTrGm9FQn0rsxjQYsjR3DpT2Lc6cRdr
zQecGNWJzUnhxXC9pvSSvWrr80WT1cLI7mXRc4nIe/f5AT30lBiyCwp4EmyN3JJNSrq2Q68sfcOI
b4ivPH21XjP+VkKfyt2Dkx2T9ch4vkgygxkNkfG1CsMagGJqWH+VnxWIrZcCxxk7k48xxtf6J4g4
2CPPLp/Y04xy06d7i9CQ/bP2rdSq0S1py1HFoYACpEhdCNvo0bPdMkMkvryx9hCK34K5qEtCD0XW
UPP++0sagXkXJkxWdULKf0xPJyw3IXlGA1P5GBcQdZK12YgRGlUgc9axI4wcL/IQQMbifZ+R1BSh
Ael9J9L7Pw4aZVi1WpBq37qafofIhO2FjAbunrkrkI0TngEE+oi9HDFu3Bd3JVaV7g8sNSKCkC1G
YV5DifkNGF3V1RlVuZgw4e3rVADy+IJ3mQJj6lY1gv3rBeaRd9l6w99dwZMFhBz5Kmirx+HgstGI
u25uVmRle9NRlLC7+59g2JR0OcRDhigz6a2fVozyHw6jBhXQc6LnYU+4kjQ3P1MmDv/nbDceHA3Z
shnq4mnY2hEqYV2Gvq/Fmsy0mRr8x+bcED5WFaW+nPjHjF2DMtOKLNWKp88nE3sANmDNIok30P3G
HM4Gg7yT3bB5xC69gfdQnlUBE5ERs5yf+aREJaj1CHHEx69kD7Rx01x6uXtdo0wo0jMcFkkgSFyM
YeMbFS/udmghksdN7fTPaVv3pcG6iCTGyPS0oJ4yIN6W/LwpUQB2HOajWkVCxQfArckSGkB8HKan
k4VEveAXKBXYRhn/scpXXND5/PagIJJyrD3CCvWIAhM/PZ30tdiByczqqYXJaeJEPt84h1v/domv
jD77a9y51FWhzPASlDT2oFU/zz3FCRs2aYsHLONg1vU4qA/fKfndzAmYE8ibTPwl3vjrRciqGE7l
tBf5azn2DrotoB5V4Kq9kjBS5ejJVLAwUz24avHi9WEH/eLzGi2rngfvLr8XilDAIvyGWbYhFoHW
l26fbG1XlA2S10JdSdViavkafeTpyxAcZJKBrek6+EEJNxd+5m9LPhkB6fNb7WzJ2M/WJAobrV7y
zjVg6UCs1PrF9s75j91pzOC2Q8W8JPzeINSn6jb+l+jIWku+RSAVtQjE4D8vKVWVHbNneQkznD1i
Sog8Pt3BLwrkdqTYuJl3j7Dbtb0rNsrK4GcnRY/dQpIgp9ugEbCNvG2t8b5TXQesXHsL/ahgT41/
mXljSVyjIAqwiTvUYSvZYR71x1xDxU6MgX8MuUP7B+R6Lt+P1vljJepMeF6jZcwRN15yAX2kYX1N
UtP4nGPds8ACQdrcI67ZSj8SuV2nzgM5pdEHHKkVki6G8VMP7X2tmLh3Gg1qW4CbtGPeIsXJTCKp
xnTQUkVSViSQnVUpdLG0WU2SvR2h8s15NJlp85uyn1BTFHlJ6khnDvJjsn/FCVq+Xm233vunVy24
qXrqy+UObJ6rB9yIaSfk5Yg0LjrFOd3U1ckS8JBXZE3n5Pw0YuDDu4YSXv4PNbmt2XdxqZWkP16U
YgbFf/zfCNqtsAAYCSKEP4VgqVl1j9PICIxDFBzML7AmV3n2fxpfSUw7ALr7MMmVVH8gCyZzqfRy
HwK5F43/0yJDcMU4T8SxJbrrxXyaxFXuWfLhp7dihTl7QirqVYIRFBqxzPb6IpOky5uLIVKA+YiT
VQ7kGONL8II3+3Se7PgplSXo4j7pcjamG1C+127+ctyVL1Jczai3+VNf+i+mCEvk7rYAMYDTJE+A
cSBGL6yPbLNtY5CEgN9icdW0wVtQBqZr1VwU4wL4hmIhaf+C5GqdiR1mRZpBKWeIMuMcFzFeqLzY
Zg0vP+sCzXAkHQ06A3dGBe+Az+lYvWKwhhn1o6wsH1kH+ak1Vi16Sy1Hp/Bb6yw5C0y/cm9TzZfJ
Kq/mRUtFr+vvLCW6wui+deF2zTjX7YFnntZz+6FlOBvN9uyHJftkJ5PvHYnZpFmtvAACEF3Dycp6
28tQyB3OYOHf5XNmaSKNQun7VY2zxvrzQGPIr8Vq/Rb1tqHLvb8nE/sCwOPcTqdkM9PkXndRnChm
zIavnZMT3OJYhtR7kJ5f+DXhd7QRAcs9Y/KuMa6uufUUBiMG/tCjJKTftb5sOHmrYaWqaiKGTq2/
Yht3tSdRWOQntomjJEjFIyVTIdGkKJbQ7J37It7cnSEEid0/kNROPPTG8DCSeFtDZ5W72uze9N1o
+bTD/JgL5DIQ6EOHdgg6E6KrgWZMOD8VDqvs7aDY1oSRSgCt1vvm5ndXeVtfoLilLn04yI0NY43E
1QXE+8y1Mxh54BhdmpOZvTsoR+6kYzcIyDNwt+OUB6pyFnLxh+52rIEeKkHxMj1bn7fo/9xABmVF
qwGykfTD0MLy/4m6RUrbHGb60ZHqZuWhCvJo6/FdGInEJituOJGu9EQ774jmzwQzdydrqfEHGSe7
egpYdQ4WNJ4U/55WpeqSOfKyGkyAIETHfTfRMAVcVsroiKfWswQJauVokcT0a3QSMp1Vv/9CBthZ
3UJ+32t6tM6MhsoVyOv9RsYrG7nE9s1Pq52ZkPJwmsJfvMCWgIlCNvQV0iUz2R+nJc+zU7dRqSex
7INNJdb3lzc9ZBY4qtPKK2RBDf3ruxo+iTwMbbdvVWX8WIv9XR/nPx4WbeXx4DrXlw+Hd3w6uQwU
fxjnHa4s/XMzwdzgeGQAws5kGtiDwpfdwgir37ob4qp9lTBarI3eHd3B9nN0iite2xY3Vl7XFoyj
Gfye1dOyEBNDBgVuRiDl0owjGdfISgf6wayptXX6d2mgyqQ9nk1fMkeYtEaFWwb+UAmsj/dTvLgm
vdSCuuK40xF7l+cBW+ASoRDNmqZzV77zZEQPtS5FWNZddUSXeFnqdCtAO2QHof5cmu2lPT8h71VR
qhT/Jocq+sIEf+h0gGOt861anJ+HnJicmJDs8FR0km3laa93Drf27xKa+foaUbBiEEKqaaLCkcu/
VBcbW9AxR9P8Skumggq/Q831lxzZL/lK7xsAwa/n1CG5QMVu9BY2miEdkh16M7tgre6BzM1eIFr0
6dWQBx3pmRe1y3OftVZ5cKop+nvznBzMIIUc0ivKJrg4Yo0q0LN9tVo6KuU0KGuzcRipDdvLRdpi
ZFmKLtuJ2YQ46KzvSIhW/wH+sI0C2M8OgNONhyOWZTD3htiwHKE3jqFTPmS9Msh2JaEvz1iqePKW
7FRnAB/hateftoiEoScJ8QJivzdqS57hkKUmmdkOVYp71xgSB7MQTwByvdHx8bqo0pjdPAh1AO6x
/idffNj//9nlfvfKKhLILSFTb4f66kx8FJ/F0wdoyzJnsArmNqqv2vZnWPevBbKZRCNc9rzAfb0a
ZcweIAsSGXzL+ufF3ZkatI7a8Rqq9orbi6gyFp41BaWo6vpk6oRJhPaycQKJXKFWtiRzWOvWiR6K
nXmXc0XeEpel6T3ffGEEzzWoM+EYXAmSIwlaeuB2r+zFzKPVG+fMVyPxf/amsT/7ezAMqTP2Ummm
IVO3bRzBrPCdFZFbVe9oMirvBOUjwSk9JPTrapcRHWOsA6jIljvTCiUOixyIXMPUAIJmV3dRVfAL
CWSOSBAIuB3qi3HKEyogpqmS4UOu+GA4SfGu+bwFac1kRYrdaJmnW3P6/49vEDSDiXPuIhEaRRRW
rcYJv+HCbtNnwQMfThtomhwBQC+OUo22Zh6U7TjIrUq04WU3Wb+xFtddw3GfM8W9kG5ZW6E1RGFa
On33LFH9zEA+hMsFT4yOsUbZAL7Yyj3c9xVQx2DTwiz6IooJJI4zvylTHaeo8VIujzNMum7diz42
hiqXdlw50BJRAo1ZZNgYTnYhXksQftqtWY48LYeyR0bdl3BnJ2PdjaWHvg4zDbw3eSI1wBKerlPN
6uLtfCp7sWF2x5yLKByJGus+k9YKjqxldTdVpZDay6rS/QV5VAT6D8Mm3IY7ClnI4THgwPLKrPoh
PnxRNDXywI3/6CRUV04oT+H07RA4StfFxPXmTYdA6ESgubhjIiD63zXEMhYS9EZLVWeoFcEoh5GU
qGN7CurIFNtZ4vul9+UXXqtbpWjTASvP6e/tOW5vpPZeNOICZPcMGye/DFqAg7I5/gLmiOK02Rh7
wDcECknsEYJ2fLGoKw6fMBF1IeTz3q8IoZaXqCwBOJFJWidBGfJu4znCUeZS9vTbpj7SK3faAAXO
NTfp1QI6BIam1h10Khzh3rMW7vSOvaJu9895nkugejJO4WX2kPZLzP6WMAbrGFbU8Um0UlX6IC3U
vpm9n1X/tjzWX7aIqWxRzRrvlKykH8xLgnpr7JlLvEkJH8DSlYk+XhaobqeTG7gJXpp/WllgLvlM
X1tSYkW8AmB9ySpnU9ZCmS3RDqN6exNELFB7QCMTDFvxei+1FiKSdmtUiJYlZerDn8Y/VzdUvoeE
/d42Y0Cge+FcYiynrM2wZtFBvUc6rWs4wqNV+9o3tsUOuwydO697Aan6QfV+GiS1MkXRKkP/tzj1
esuFtlBoRHjBpuDnkfv+5XHICwVu/xcKBcouXeGa4JnkpWwB9aw443TfWkzfA0xoqDVQ8Gxj5RX0
0MQwoGMfe+0qOngqpOzUBGJqXhUy8onHaBID6AAW9mjrWXqMjUA1//AsV2FF0t14m6pgKr8hqd3M
9d3iM1F7pIrgu0SX0KIGxPGxISv8A+B2xc2dLhiB6q3h63H65xDlVe7CJ7PXGIEz1Y6g7CuEBit4
GZxgBavHeOcE36JzHyB4gwN4ihoOkRIeGr3eV+IHsaPNcnBk37tVl67gmEClL9ZM/STChCn8qMvj
N7zKLGIzUg9OFdBkN/lakJXTnve43lEVogffCABvgnltzWHBvriwAKoI0TPv6bGcIm13Ymhcqzss
mDiQxbHelLLESHTXi7RYcvwgpQZ5P36arZHNr1TAg8fvLrVN+GRsXD1b6A0DREEu6oN2h4eLUwwA
0y2ylHox48Bih5OVedDB/jP7xCk/gXZXFbwO848Wg22BE5AEgUbAmsnk0hcbKl76cIHz6GarLhH4
yJPLw/AyY08bvn+sIpZLuVSeD0Kf/yoqsrhzy/RZZE27w7E+Z/f2vhyJP3TmIC0i2AqJ+9lK1F7K
e7NAMSWFz/+DHhx4PhLvtjcjYhrbhYFPNoM2GR8I6Vfn/6QkjypSB88f6hAxYKkcAxQsniYKdZHN
F6eTyTfPidhgUWbi7uS+rm5fojRngruvJKvChYe9f1ypywrsXqw7v2PMH3DXX2GOmULfoK6Iuj5O
CHS3kX1C2oPhtvcT9Gy/F+El5SjhyPOoaMN+7a5rPtiFBhk/Ms3uzhY+OmwabgEROVKoDsA1IVYu
0lgifayRk5Sl6KYbfM1IBnqId2xfoLhsGThpIzTitx8fz4BoGouPKHSf+qzxpFwnaH/Ci5UdwAr1
QFX9Yo8XntfjZx1S590CXjV97Dc3NkuSJKef9f+5a5jfa5LSs8Z1GkbeUwJ08FFKf3yQG0cYoCxr
x6iwdMmiWCsU2YoTnatAbZPUi8R29dUAi731BWbuianEOzzG8msRDLes01a7h/fGW82tbhV3kfrt
qLp/J87jdrnl1fcsUn7w7/mCE94I8rdgnM7QMw5Z9hk6YU1RUOhSg6Nv9jgw9DuPrmVzZpVmfStp
eW5RGYuZysysntd9an8NLqgiRw47zRHXhCpxGo6PQxOoMz7XsLcia9p+PmIWbsMTg1uuv40BI2NY
F3SHEu1gNV1tDCbzXlgZvxkJsFQl5RpF03SOy8G0b5BozKhnD4u3LJtXnZd0noGQGjdUQvbnsBQy
ow8ngSy5SKzirVnQt3QqdWIvAyB24uoR9HqFbdX5UmA2dKRqTAs+w8xGKg5b7omexRgUoeGRbq6n
7HG9cgUsoTVbQx5SAhjXBVdIz5GPtG/xT9AeNppUnQgd/9+GS8H2L9ftARzEcCupO220hvFlvU36
1HGENwPhcdK56E3/UE2J9XpfjSqls8DuKh+dem3fwepCjTabjl1JW4Uj9anK2JiD84wPTftiwYmo
vdHzZl1H4WTk1WrPj+OQSiPa3TwULMvpgepMLUG7KwCP4MWMXbsk2D6VgMDM1YXH8OBfaPX/54SZ
o4olWH+ZMIH0OVxLbNcli0OYbdTBk+fQ/Ldm0HoZVVTxyR2uNIZmbuKkRYmhj8oJqp3j2bLmi0KI
3OrLpaZxSsHmWxKj9AiPe8qaGiNBWdXjon9SxUtArdixXigm9j2xY1jnXlmLp4bso6PH/IL2uwbG
FiD0nYu849eFGF5TaV6fUesQ0Kk8fYn2qGTd7gXE2Nj9VREKvybZumbF6ERBS+lrnHcEslBl4grH
RQ8V2VFXwF5IVOyucsQ7LpMSBMSuoLIRNbZUM5Wwx6zks0DUcaJLvzyH1mM4nfvu63P42yp61lr5
f7b+3vfSsMToGk37Tc9ZV1cu+TloNShztYBwOkfjiE/1aA/rG5tKPFtEydyKVO7bRsL+cAAxf11U
5oaXId5HpPbsjfJ7Uut/LdMiIImxPRs/IytNu+XfM8RIn9MG+dNvUyCPGbIkaDmFU666nqFm/Z3Q
eH+GVL3bFzTB7yrb/5sap4T/LgibKlHZokQJRjPXRuzEytJQ52CTeDPjG6zJEiJBNWHhfLq5yHCy
8O/QdSU5r7BH16gY1+cxfdqLOTu3hOh+nFIihvsKWEqnR9drLcb7/8roZeYL8++K/vT2VLjoRVx9
U2QLmI7N3lk/IGT8Jjv2uW6juU+s2RnAAhH7omRZRMtNWL9rZ5RTgq6gfl7Eeq1pqk7DCgaI8l8a
8uXZUUk6RpmKKQl3cixDNF0HKWHbWAIUR2B1N73X1VNh/3xh+nz4GdvbQHpGKJ+WcS5OI4xqJhm4
hrIx1uELtlK2YrOq1D+iBhnfYApbq4ildatnF9ozgwN+zBAdFeiRH/T5rwSRy2sN5Zpk5Kc9osRt
zjlhPksvOEMlw9iNWJ2HaK81J5sxCifmyQPhuSQmVav4lusO1VGNw5WVZDCoYTcUnWz6Q+68N/U3
bmFASTsKLsOWPl3lZeubVN0WBsMj2iI920vj/s7EAhm+9nbOWVtG1247DZ5IocXQmTuTo7SoQ0Qv
7ScE2bKpImNUMAUl7ob4hop8kLG/b+JOIOvn+ldPPAGx7Nre44LdCWZ/CboRAAgzKev6v3VNV1Fi
5hlzGxVD3/INw2BWHisbMajApyHYMOmBKUIoB+K2Id4Z5u1t9sr3OCNnQ1Tyo41HUCAhClf4Rve9
PpLHlxtSXb1V1wtvQhFDHH+LRZxK1YxyhUqHJ8aO+uUHMt9QeVe1abbvgIgGtZq06VJYR6FFQVzc
lUj4dCghNj7LgAjLLklJMpsmzUE0z5xRM7OzX7XaKO14e5yiLu/a5mms7ADd4P37MIxptXb4SGw0
pXbTfWQyqbwePG62DCbWEpP3ds5pa2aRItpFBgePYB+Vk3n5qocK0O97rcjObzF7rN40CE04SI7D
NJlsv9rFsQe6dVzVjeljyOxkiZj7I+jfDsIl3z/6+4WpXHMyr7QgmD+NYMcZR2M1LJdla6ZCGX8d
/UtLYhMSDBComI0wnZU/7BREE8DrRIhX2vy8auIxLlaEp5Q02n6KWI9K4ZXlXDtL2h9KDzO0KUi7
D5oKdCioRopNkqMRmN5Nj/J7VVpnSZQZaD3/nxPmfhYblPRxIf9e4DL0s9Lk5lMNT2nxRiRcXbNQ
Ksx3K2/FLWBA0ZFdyNF2MzY79qpNb6jkHvKYed0ofNTWgMUY0iGFWBowkSkz2lwLxU/kf5II5yuC
Fe0yNrW72FYOsiU4uXWHT9DGbXVdsKP/Tyt38pBCLlHRIjC6AyBenGInoV5QSpGQPgm4A2DI5MH2
XqzP85r+NY1CrUwK/qarG4J7qrV/8XW0O3Cv0WKfPGq5cv6dethQEdrKWtRXtmMuMTV4QaBI1NGP
Xx+/uAMrkc6XJe3F4ajfoMFVRmGnwularsmVL6uJk9cvIeNeA9gfDpZQfi/73eKYg10XZpk4DCgV
bRirvAsCN7xuQ/21k8cetga8BDSbXfUD14Mn8HZS0GYIGtKDS6AjXk8Idnh0G+xhaVhR7hot1+K2
rcfA6ybHPa7gCjc+tN9VwqP3L+Bxq+LsUY8IzBTmus8n+qRrV5RfFKIjsHsDNDbAqveEL6jXCsOV
GMULjCEN12jBH5rJjJI10w7cxfQhky6utxXeJHkn7aPRxysxeYUosckJfZHSTadSnW3b8M7xi6aD
Ep2FHJMvXl/T5idiQFZze4obRdh1XE8ddtv2SI8al3KmtFs1QlOh4QOCSakO0bA720pggH57RMAO
avK4dY3uHVlVgtwU49tJKR+JNR3xt9nERDHQDf6uMIfc5zYSB7jSfzqb1BG4qfvVOZifPRWZTIuM
R47aalp1tp7uYoLkRt3id5NVUogTKrPCVaS/UxUvxfEbv20/PN2aBgfafMrEQv8REqDCcouh3zIH
xo1S7OeAzxVdTXFQU0SBoWtzJ8fnIGbVqNBej5zn40RKUjumpiAFw94VRIvJCv3Kpj3xdsc2TaQ6
jAvJcAHX4VK42SGUDXnU2ZRhknBhEKIgFU9ZPJm4VUMy/37TR1MhJJRyuMF1DJ0djdK/oPaks44s
rEs7gYTtPZXYe7P10lu/1SKg0Z8qWz1JqomJNUWSEYBDWckrvTr6h2X7HNHuwuG9GfDZyz0kxhoq
9rav/8ozAroZnw77TtCcPcMb8W32AfcEetOsdPQhBncJwiT5csukD7FkcbSfhS/k5JMPF95fp+61
GW3nriGq0w6BvjxyDoNQRydcW8rKCctV7BIcJpnJraWg2Mt6JPvsEVYFv3xgTdZDHv+z40Qxv86z
jMTjbbaZdaR9+LW4aSUfxjltp5qxzicqOY5I3PTWlAZU9p5hAd7/+YsxjhTAP8kCvDZinFGOZ+mH
wN0lbcbJ1KmWiTX/TjA5EFJ881IzuFIWHdbN4DmESZl+xawmgvcmA9IbGIjOD3Am6IlzV//NKRKP
HggDolmQLi9rSNXRwZ4ZXrEGxj7TJC1LKJLRoYRNhjqnI9m4fACbGjKM0ywDyWwp6UPEZxPb6yP2
SwNnIDPsot3fA9YRPq7IQg7x3XwFFlEJL4i8awKm5MqOR6MXSBLM38vuEEllE5R3roVNrMHPH9lU
IT26eFhazTMYKGwJJpYZuTdViErkYxmnq1D+F73FH4HMK0NR4C/dlxDwKsiOVxYJ/F44UT0CVsDq
Pbz70iH3O+VHfYIFPuwb2qsODdza2YTF9DtpvLO5LyyB+1upwd5X88iwZHYHcGygrlS8HPopQ2qe
PoeHd3PN8dMS3qbi6vVIpQeD05sK5++KWfg+xKKXutj7eV3AdHxO+lQoUsAhwaf+12IJNQ+8yUtS
GhFqlyc3pcPcsmpJd+HWPzaPq9cFdUeLJ7WD6o0QR0BTh8+kZXXyEDzWOlcDuXOEHwpVPbAmTF2I
s45zPc9IAXmPN0I9HAJtJN6rocCSqhrJkPNjzqEnjZwBun8UqyNRzjZnQzEXX0wTYrBwFqlx8HiS
Ase1zO2ZGz4irKUDXjc5oJNDOfpi9DTVf7qviguNFJnb/E4dHggNy9hsV2i01K71QK/XAwMVj+84
uh68kurSbqphufMI24a4/ZL37KkXvqCY1vuhSnTrfU97BP+/AEnoSbLmyzVibe4IBNZDIKmpw+oO
VkPN+dQ3JmTQ/gLXclAvoAAlmaWvOUzJ/ka4BfcoEtpO3DhCH6/wrw3ncV98tijFQrAirQkQPpe/
HjUj/o3i8GtCyRIqUSypEYprUi3iTnHTdw5uIVrI3uI2nezCFxhXZgOdMl1sUDHScMStr5/CCOcK
AUTkNhV3jnlS3XVhQ9rtUCRccru1Of06tuqRoj7zfqxFUVWwEFZ9oMakoDjToba/KTY2YfPaVm7q
TPF0T7lQiRIV5ccCwh5StiDMOL6AIr5OeKEKlJFFEENnsdZHb8NAX8bcegD3QQpkycclFuZEVUHk
8BACXHRxDyutI7b2nf+7IRYxPYwpudJkwDoz5tDFoAEb2tDPMpLMPb1SsYNV/uq8PHaLmWsaQdLu
CmohNDEcLjbEZZ45iJ8Ya7rknxI1wq0XatP0gLcNGIahWUxyjdIc6jx55mBiqfUR8zuQi/IjMgRP
VhS49dfQw2rfZVIgFlTKrIQjoxuIeXNZoRi3l/WifsvCQeRSjc6pEHfaeHCPySvTP2Fhg3ZG+I7X
YCJ7zRJXNFZlSo2tM1GLIIDAXDC77fBGeCFWaNWGJu822iOxxsceDpDYeD+aWUGuferg6vSTJYQR
obc90MubwixF7kM9qJl5eAs8ab616/+F6QE7J4EeMR1YUJTNSVni7kWQw2lVWwR/0+cyYmf9sUDu
OtAYz3fcRTEUaeiRHBRYK6IrWHddNoJuzY0rRia1fFb7zTb9YApbWOO3OzGzDPqEVhJ5Ctvl1LJf
dehit5SUL2SNVHaQQ3EB2XQuHAyT9aIqk7lu4Q2ephpYRV3wb6W6Af7/yDfh4LXbQv3hDxPrcIqR
Mqwz30nY98M6CpXpBc5dqCpfMo/xNsbl2WUqFqj9qASr1dwdI7/ftZRoLXZ6L8/WsLWZrVZMidlV
kEu48rNvsDKMllLM5M/5hwqcUghxVIwSGv1YUPkZHFhIAurIj+yLg3BtR/Hw1sCh1hFgTIrGeNsT
vh2lBGKmq5//OGFuxpDSK/pQfFJKiDs7iwuj+w9ugD3/Fve+ItuTwKAr60rJCFVSRMkKWr/0cLPK
TXwknR1dCyjX0UbAsTDzxXn2rhfrGG5e1tblztKE4/j8gPv9td3OGqG4OPHwLG5hgBcCDpAC2aiJ
ZNkMjtJowVKvtVMAhr/t25n5GKXpleolFzDwe8KE2pwAgRHQuIejajDhGr2EGowCNkOb6llCQnWj
6NgmDWoSYmT+0nbPU8MdkHdZpxfsN4oTwyOeTOO8ywhB7MRTjNjka15w/GFXcKCvhiuglVeZXf+V
d9jHQYOnM21G1kiTPVy+cmm86OgT7fy7fG6IuGMH/w3JKxjM2yT7CidvXyJJrvLrmGGlhM2/H+RY
O/Avmivgh7IT9+2uaQ+u6o7Em2PZjLNPgAiU3RhTa5KLMIF9koLDwggfaTiSqnhoOi0SUYnDBSxF
yKdM+IdeE9ON3YLuiJoVz/Y6XzCIfk4k8QAnm/Mw+z+buQG3n7XbrdgiE3tXLrBAtmmwK85Vi9MW
HMbMOufY1ZfI4gyTR/NSDIk4OF9nppgnxs6yjyGC8YdyPqcXC8EObunELtiORYVjvunK84Xia3Ip
49qxvQE7l+o0QlKHMWm0+oRt9hHxLLdGo9ZYEqGR8/tYYXGNWEDSakBdMUZPIGTL4Ya1Bpc7c546
e9dpMMpgnsdNDj49t2oxcrgrIcCL4e5HpRbggAMqDrh7kCh+s8z5vGGS3Fa9VcBsTHSIqUfOxokS
BR63Daq/tjh/y4LcehQ4+t9s38RXVvuF7TtZwjSsmogGZbJfoaWqfJzzdUB/GXIAeSsbTA6gMvIq
bFb5QKkcjc8qObcyJXcOlwfMZFLfbfQyFib7Y1OuYCYXwdqb3jnQiGPRlMurJIvg3VR6AvBRt5JU
GbS0cb8QJ6lFlCrMpR/WKkylp5uus7XncW8vcqmKyawew0Cu3W1kVxn/OVfFku/ZrwzmGXNJTqho
d3109w9JZCysyBh6mN5mWPocT7tjuEB+StAyP9FJHdvsmDN9u4lQF/UgN5JHN83iZohCFLRj8GC3
Fxslz+14JqRbLJUhJczeTuP+992qzhC/ir5GGt45/wuYCwQz4KCMMp8RvABTFg2DerzZusQmGPmj
RdV8OjQNLRLTRBnsaYeYZ4u5OF7TonaiMRq3O60/bUMkQ8EouJ8yA5GtZftaWrnG+dP/pW3hSpeZ
KqUOqZ59HPqS8hv69yYcpSW0KFaGKb8yB+Nc86658rzyQK44XyY+Ji/gY77tIXYYHNMWpXyAEErt
u5xK31hDQW1fDLTNGAsrdWaeXS++gWX4V9sKd2foOq8mgHwlxyor8LPwZQGsDMaIa7Krg8FVmIil
1Jyfia7A/28DfYKSqw5+D1gPhNwbZF6yligm3JliWKU0vusDdnRuW61Lscf8AzeMFB2vdumiPV3O
LV18Hl0TLHDnKzYTeYBRMf8YYoTu8fS6AvyjNX6MD0pd9ztmdBVbknLPEwbw/1xVaRooq16OzKgQ
jSn1STv7IEuwhu8oijlOy5ZTkbFZbptmhiGqzIN8yYcemv50n/g6oM2x5civE8QiXKo0lr3Np+G0
w4w15TliHgTq16tHvkTTxNys7bnwr1qthPdpFbb29XXf5RFQc4AygOC1MWt7/BcxeBOHNLZurxtD
BuQR2o7/HqemsNOncPITtWvOADLtR14WlEcvQJSziZAD5PfO8eZKZe6JZc3WD2tPKi+fOA1G0aRa
Fl7Y7wW3cnS0D5qqGp9WIfst8gnqEY3zfQTtaH+njZ/Ah0usXnKirQ9pXii/3N2eG+dVm3gkP+S8
fpW5GzDPZFEYhMknbNBqj8oXzmlOAjKqL03+bRstaslp3IoLCAN4J3XzrGiyAsnAf3lns+5Duy+p
cBCnlI/yjr6MDqG7P5IQv6QT2IPeUsMTp4z7kK+9PYOvT4FPLzxl44IBC3p7rgoVrn1vh11zyOyJ
sNsnKRyMb2+zz07Jh/SHUJM92N5rNM3suEdhYd0+cA3AS5+TtNRKvrbN686KxFciRn6M49OHL5kx
zEq7Aj8sZhtRp1Ui1U5KAnNKOorIzR5NFHb9vmeVEfDTF0JMfxqA7dlTnARvKM6yzc4cF5HrDhch
lJ5cFdFMpp3d8iFq1oZexzC/KunccbBihGVG+ve089vpkPTA4F5LQzjSkjwjHhL1EunTtAXVRhPW
/Cy39tIkuAb7uVynxdLCAdvnJVqgvwom2suHKxlx0I3XJtrsXvh0b1uOgaPvbnJH6Jddj1V6Npuk
kiBGBRO7AEbcjIFM5NQ3CgGrETa7V+WqD5c/4PdeidZBYLoTmptLuVzdKEZefF+W+LDhNMOXUXtq
fQdOmLy6Sqin1p+hYNfzz3ezOpDSx6ziPw1vhAllO6cnLF+bA+IrmpOYJGJ8AxeF4TETrszZeO+5
2Xht0FfFC8YaIdbM2fgYGbsBYr6lY48XZ71V8pbXI0zLjWMcBK/aaqpxDmqzbljDqHp+NujnSRI0
QQj+MpShzcXaBD8bpZI6fMZGm0vMjzSTg2vGn/4eyQ2dU7bOZJhYmBTiRiwrx3hzg0PKZ1ZCHnyp
oWRxvbqD7aLNVif4Vy/Nfm2tOOFd+FkBP5jTrcvTzz7Msz24BwnaIys/96Xm/oPvUDTMKPuAuF+h
vWiLHp5VtjhalZL//r9jm4dCzkQo/0cUgeJdAJ0/raCSTF/FVNJYECXe/KjnXVBZeBOFrd4GqEdA
GtBz6Kq27tT+PBzMzdPLYg+BMc+GAfSmcfOzmizqST23dIusFCJ6hrLipiAq8FeSe0wUwfkOLbcT
MsdBcEQRg74kecoRx2o6F0rmHEdsJtVpb2Hjm/ghSTh7ruShIh4GEKtDBqgnfkGscI/oPF6VaF2Y
PAgVEpiHRJz0J/t6jYSU9H454h5OBNw4P9NTBmygSgxQzazr2Lr3QLK6zYwSJ1kamVp+o9Qe+69o
AUTlFw7/TTf6Jh5Kg6buXivBQ0GDhDPmt7G8PHXK1q2COhlseQ/93cDNTjrpdXpyP7XDbI2PmukO
DjNgbBB5u/MkRVXYOU/GH/zd60FAJusyoHwZKsABSrAJtH7eRhXTIrMQ1S5RIsuGTo+DDNMQZwlV
gns0aSr/+du64Qmo/mP3/Dk345tDM1YF9RHShlmTRdg+Tpk+evlXaTHfN0kiihLD0newEbd6YtC1
SDZdRvbklit9YrMfwAr/zcpa+43pUz93lLSp84uvHRzCmMCF92n3tb8X5ley03OYRMSc9Mu+PIwP
P3SRWNZzAMQnzH9F2UM8r9E+oAOLM/IsH4agTXS7lAitx04xFRUz9ZCqp0om6VHIFn7UaH9qVTiK
cUzz5b3RTTyVcxoNHd/G74c/5W9b6SRx1NXEh6V7YQJhZa/WGNEN/w3eep3Ijo+sah7AJpN7yiG2
gZbjXWGlDjpPhIGsakSUZ/G00xPKl0knZy7xgtRX57XNKi307Lh6+qaCINz98SgEJvCpxciN//7v
YEYkTdo1N5yFO5gO32XMScmyWj2InHz+HbC3JuLKjZEi3mI8LiBANnexepFreA/t1sx33a2vV+XD
bPBhH760IwWincxb6KrdwzZ93e7zzTxf4Mypmx8BiFLTWNiP9ybAk2BGV9wZ+UUjV4IkF7kzBLGc
dq8DVhnfj3E11e9GcYG+DifZ2eZpSFon0KVMduf55lJlFWgCe+5tDmqF9+sPCwCOgyHblhFLeq/O
/YkcbF8SgxVb/hgJSEz9VfhP+Kh0/+9/QRVbAGxszD8N6Yl6l6TSpPevmsGk0Fwj1sux0WhNlH96
C4QvbA7aeirxcTeKP18OXXo3hxjGSxZB9fLEtZh8qev5lecprsCgZj5jkurjvYmdNBRxNAhVOu8H
OmFbmc2IcTvCT+RvbGMLh1NMpZsUZ8qYnTSySZGPSClksKP5cl8KsKrDcibpWrf3nq2ttEruYJf7
qJJAR43ea2IQso/nFjhXMhNiIvs1XJt4+13DnRRhj9odzQtQROyKG8AxbFUwgkZsLgxYizpcv0+F
blZtM4sHmSvc1Y2PPXTW20blb5oycM6D7jXG03NijL4g2u/eCuZaaAA/WPW4x0xY0/3GFzwV5OB5
sH+5jRh4W0NGzDeYiv7FdAbT6jcZ1YKOgBmOWEbwomUiRsfs/eW5IeuEtjw0d2cVr+8loyteiW6V
5zfbAVZbX63HJWhHXmTQcJRRT6cJKr1CXADwUJXWuG5YydMiFLkjD8AzO8P0vR//5Bb4fOYnGb+7
1HF2beQ8hFGpFyL14vHwWkyKxckS70BuVUVwvTUaQH+TeW5a2G8TJ0+Ff3khk6GH9Z+s3+0wKG7e
ttaGZ4bUJr/ClIUHzKaRZVCF3BQGJm4uwBWAgwJ+naFj/rlz0oPVZsMoAM6ShIiKwEwb+go88uTN
HBtDLAsp+aj9U2krTcnWq3TNhFRpH5wE62kyc3ITFcuvssl2Mb855K+H+ET15A+FV6lkBll46h+g
7bbU+i6Ftat6n5VUaQnWZUAtDEUngD1umYEuFMghlmlcs4X7hMe3X1LGcObR016P8enEqyMMbKJT
9bkFsyw3Z0xPe/DN+ODMFD3YqerG/kx3nOy6Qa6OldOQSe8/z/8I5CZNqBC1StgzFI9v5+PElDcq
31I4rwjkFF0uowgk6gki7x9Onqdq8mPM54CQfT205kfCz9B3NNG640zG3MvZAx+ZDBYjNU1veU0x
UqA19wKeIrZo9ie7a8hNFeY7+ek0pDNZc+X/+l40LM060H8rj9H/AeY/pdsH4KKiGi+sExwHhRPz
MC9DfPnTe0W1u149s0g+ksG4a4G64EWC7eqmDhYRJ8D/i3nUddWIDsDe/gB0flZjlKZHzh1aePNn
OP4zvOrDDPPscN6swiswD8YXeOKCgPUjBdEOfWMiklPYvLIRWIO06M6zruJ4O6Fh21d0t9w+HGdn
f2vbcJVTsa2bUZVDwlQ66JFtmjlTKcXIA+xZVjoPLMud5l+hvY0PBpHkePpDBbLrxKfYS4Zt2FCG
V9kAeid7iQWnzKU2pNluK16eGHt0G6fNP5XUh4878SG5IHClwiy5krcw1GbL7EVDwji/wh1H+zMc
XB7K629lp44J2H9QrS3idfe4jb0uSsdicCJgcEg4/HqaHNv3pz895sIML0abPvghcfBU9yfzQtwz
Elw7YtpfE7oP+zHUkNCCfPSp6ulbo8TZV+icqXMjIih/YlMHlai7GDZFQpDCKjrMUoNVjL+y1B3b
341/UaGfWHXGd85xKaa2ji+Jrk5WJYwTrajWxaYt0NyZPld6Lnx7EHSF3s1+Qp0rBX1EW50uHbqH
EjlwH5C4xidWURSJwpvTl90sAQA3OF4Ekmm2tXobaT2Eo12Xa1bSk2TtsqnXJxWoAoy6Mv3gVh53
OxQmxupQfyM/3PESBE8Zlm9Rux2jCgFBcWth9KbPKp94GH/P5gHz8zvtwoc3L2T0QL0NLeULlimO
OLmOg3kgcetcw/Vc0C37OWkKo8SXG+aLd/7VEHONZ1kqcf9sWiwtnxoo4FC1s0G9hmfgzD4hX+rv
nLLllTQBlUxRAUJ06l3K0kb0vnhGIQpY8uQFa+Hpmc1mwsbg8uCRLj0+G1OsTWwvhDrXv2Q6yVE0
WNerbUhlOgrDbaX7FKCCsstDYt1ncrEPdx7s10a8cHYUHbAIRrB3Sa0OJ7LDuT2YGR3A6f4tdw+L
8LpX0gHEq97sTFsqFwTG5ACWlmLfSV/C8/KLsmuIA3UyX8nFebzAnKUH0k7pvlq7AsHXvNh4wHwz
5nTRw6kkHXzc6AZsYCzW/nnDHXHBVFM2b4DbxIUsfzd1ks2Hb/DOvLE02bYsVfA1RdcQSkisjvrw
LlqlhX9fnvBkxBB7TVZIjhnuDOEfLzkIxmF3jXdYsOXDCH8gfmu3YhzWynDHJY1BgVC1YjcA8jEr
Xk3rFy/pTit7YDjoiA6lur2CX0pFIgk44slmprMw8BPJJSR7pc8XaTHSthdrHf1rvazgKZh+TQDN
DJmN/JPppe7hmFCHLhD2f9+fKuf+vjZQy9f4QVdaqnOGfvVMm8MRku881a0soGx/tfRrg0Ecf4ZQ
Ccef6H2pfEOhuS5JCLN3UOMXN9S5qGXwzOFiJYM7Rib3H8zGRjnRubWEa5TklKr0HpB0LQ/Z2YFr
wo5H1ZuP/TEe/LuDBsM+kAJ29w7OilhjRRlsIORSosJH83pCkSAmPxRPa6tZoLZAMrP3GpvIOs59
mCBMyzPcMBIkz0/4ULG6EEExDPj9S77Zj1fdvi680QxKhSLNWTkii74s+3AqwoQmhdty8IbEnfzW
mPJqm6vJJrGhZjbWoLZyPzIAg0VAsZDcAydXCEj8rOaszwQUFdMonKD6ZRlGIx/p5atqHvt+2G3v
sckCLNmXfN+YU2lHkbVpk0UE/naRmZfT8tnQwgARD136mB62IWy+doRLIFUAfFrAsB5KyTuJGIc8
eXj1JCOdOwZv0n/VqKvcXeGoTq5P3IvcXgMDO0hxMlF+1AVVmre0oRy8F8B00LbD5r8Xh0Fx3uZv
FO7KTcQ8/6FCT1QbQqP16mDUm35YD06takffOYcHD41NW7/OTIJ9cmsfDhjNqp2xVJWId0+6qVNl
QDqdpA4704exjzVqJ4oQgt0aeEBtSi6XT6anruwNYxwncvhXt9VAEs4Bq8qa+GPJTBo6nNuA+PxA
VWJ/wQUEJTCeVLXNEvB2hr4k28mxD1IY2WuXao7U2JAbmlyQeB1ct67oU5mJVo4NvmLmMI8N5o6h
VQ9DWRkl5oblXTY5+DLlDU6JyykiRqYEMUOGyi6n8krSBlPrDPddHY7BYkNBj+ZxgaQglW2i6Cy1
LYtjIe9K/Tk231kx2XcOMQW85GcfMN0SbcM6VL/nDKJkLP1kXbSXEhTNzybt38i7j7GveXwaCR7H
wdU05HiNTBf4gUTt4yPKIIXh7TQJhGoIhB9ve+gJkF+tup6aVr5Z6g2ZhhBT8N8hnjMBLmMAM1OE
d0wheVdF/X6CXAAsJJYUAnJLccsHRqTVj6eFafFTPHiUzuAqmYE7/twFb6dzk7kUsSIenZq8nPY6
tQBJb6k3tBMzaEw1098NUQVclKOGEIeAvHLL/2Dk1vcVWK7Rmf0GL+mDnOwSa54Cj0B1DT0XmAH4
5JUBRsozp20v4HRYPuPVn5Cx5T+FIKuP67endU44SPm9B4tKFLlFWed++A9b4cjla/0vJ2Ww2jwy
TvFrRDmVBSVTU0sGJ3BSB10bybY47Orv32zXdcLhhJ3GTOM7+Nt9MEIWcS+cg3PgifbhLMxq0OC2
PzVB72Y+1qgVBi8oB7c31sI10cENWZpe8+bxMt/5BNsokRp+ml1sJ4Oj/9J5Y5W5CY1FnJm7oRHa
oj3tGjTmH4LLpaCnyIkSAkYfo54ZRMqTLTvmMqO+INd5aI9b20SiLhhH0JMCg/3Smp8EmCRop6EV
RWSwV11Yu2o50YtRpIGkARl8zhSoIBaGwR3FRv4N7R1KUljfnqwk4yeoQmK0CQd+iLE2vpR8CQ/O
w/eCbj3jHV8YKkoDcFvvm1JRP0MooJuOUq/NxmrU9Gpze+rDwL7ComSqrYDKpPXRSVI+9XfeVVtW
MO9BmEoYG0v2Mq2LOArakF5xNVTSw3O+WVT3Q3BZq4Yd3NQOHsqLCsyOqnZNVdo0jCY8IoiD1O6z
xaCDShiWookhYtO/DSa/jqGi6dokubFhCW/8VFipmnhGhSvgYeeVLNgAF/n7+HJBB+VFSPDh009K
B4dl6P38DJmRLCYP7hR12ki4tP+xVNCWWf5CpUZ1t+nUPls2Ym4sEDjebm1Osu2b5V2ShZj6Z6Yo
abXssmPuXgXLHbKnHvS20fr+wh2eNyreOt6tuuB2GpHvKP0URphPM9HrBf85e6ErKEXrs2AhgJve
up0bNAXjihgANCSqT+8JS1Ok61e4TJ7hm8qpq8Nu9UW+xGGMRLLTvTLomPPtSmWEIZ6BoFX3V0TX
S8QwiyBCWk7rP8tgqEeFo8j+bVjb/W1E4JPyy5Yy35Xu8jxiEB3JlD9tEWHZm1W7pxXnGius8IxC
9k9Dh5xqun8j9EdHWG5UE6HQQCs7XQTdRvEifQ5EOogEPSstLpZtUPcNnA9U4onYXRWva7LqWGle
lDsUjuO6ScpdrWVLew0XlE3VTaMo9yts5cjMrayeWWHaQL6V0mOw2BiIsku1lKJim6uIzmj533aS
2FHCZw3rkznMVzNMzx4w4DukO96JuUo7ymL+0DbXeddwRX7P3X5W8cPf0tJNVK8d5TakHJfi3alp
TmF1iN53TUrNkr2qlC7LDunYzwUGViS8ryXcd9KLvbO+T8R0gmv5DUB1iUr0WD4H4aZeoNCBmUfy
AvC18MSDHYfuqXVGWAmr4kAMCiqt9p96PpDnxn/vPIJXtcthZ5vqCfsU8IHfeiwAuGlk6OERNeY6
DuhPslYkWOZ1rea64MAGbv/gF/E87jP8KTfSSg6ueet8UD4aqkp+HGaPOX9kkYTDBkrjAL39HHle
gKp8ASSH9VqFYV3pNLMh7HUn4RbLBSt20CRxUAJ0vs8RczbEEPMNCydvxu6y9KrphA+5s03rT1wN
pWAfzLniu9bHonBmbJXg5rUIqPun0VKb7M5BzEp84qM8m2mL94WErrIKJc7/HoXzlFTunCYaq7DJ
ZqXpa8+Osr0kxOdGSA5HHGjFQ+W3tbxfrRi9ZbE2YUGS2Q5sm2yPMfdm1KndZkP+D7rRbgMEgAmu
ZFgBqJOZZd6Da3kHKaCrCGdB0eCsKSFsN9FpT9GEsCCPmLfPhGjWw/3KQwJDpXBZu4Se6/VGBQ18
hGMaSXCEJbmxQ9G9XC+PX281mzYp7eVEV+m8XaT+g1NNv9aPHx4Q4qgCgKNMZrBziKMNdVdQfm9e
opffuojv2HIADaEzJuWFHNxYov5OUnupBpgfX0hzqteApnzeqeWemYRL2prZpaPpbRp10ChCQ2ns
O6giPZF4fPjonS4ZlSsSN4t8k9KKuIvQYGekkShHmOi3kKBzgrBq8QjoDZcAsZe7DmcEUs7xKOo0
8s2ZDbr/+NIFqiOBY8qAz3GSeNkqWphjZqHzLZa90JIY4nbr1kTDawYDoTfOPJT4cD/mdIKvrwFU
tO5jAlRDbLzZb5fQur9+8SE/U1uuYHbN5Phx+Cy8hNzUWrjshQXFZD47gDv9UXasEuid7BM3sK+8
1rN45LqytB/LCi/EmDA2+vMhx3xcuqPHd5+44DFeVgEjxTBcHwGnesBJl9U5EY7xdVmhovajnXno
iHBewdnULo7JNKHTuoQ/MNAhOve8/if5FyQG7FDid+04WavIQp5T7EOpghMAHKxmL0Lh4tklGUnC
d1el7X0QsKxKB+FEYj2Nd6MncwfrpIRoOMpf3ODT9388LvW1CXtuLdSBrkLQRV+57/5pokfex/mq
hlNo9r29BpDpj58HZTeF7WXGo67vViVEZfZCdNWHP1uLiZK04H0FRT9P4+fSZwra5qQwbyd80Qyi
Ksi8miFCD4xg+porj95zglUs3zD57bpOT0nzJuGnE1WCVTymeQd7KJVoATaNOlpT8GO891MWHpnc
Wm1ZxSrd3XfvYtfnfnJBeXoL5WZ1o8tqAgC07/Zjz9b3sk5hnsFkQwEbaYLvfT18EwsrVGO6oorx
IvWmg6EGjBIsgnps/jYwlq0WI2eTjrv7FaLZBKIXxm3Oc/PMV0IfjrrGtM5z2/1QseBSwVF+fuXw
vOyKXNZer8g0hy3uZkO21pKr0PVmIJQkonRUDNcxy79m9N9SKn2DksajsQhYpNLtJP61grouV2+4
UuMu3Gg9c1UwhFei6WK/aioxQByqSWb+RMnqx4jM3v86A1KeiWB12fyK7itS2SSnFCJSjBEFfzWO
UA8gk0kG5ZSRtcpMSoFzOtUJQJkAQyfYL8zyRS8Qz66Iz6iXZAFLt+hO/PUzSdk+rL8XbfVq6IJN
8DEITyXKv5SDUaPVlqCdpknZAPGMejkpupBjMsrfafR9fmZu4vcrjf+KBNQ17IssHa4eNBp1WXSs
n7g6AahdKEeK7l4gici++ifaszVtJm0mRgD7ttivgsYsNqaiGwOD31ERC5KQ3J1TXdbiBRNGb80V
/JNG6fV7elSEmTlM3w5UcP1UKfRmpP6t2G9d36dZBdDFYX6vOSqoRjO07AtKdHJPr1RJI6vhezK+
Vg1LXBEcGhMIzX15oVGxHZ7VPxdRcEBLOtOlPbQPN/TIlomPbaW+Xjpb9RtglGb7UAR+5tAJqayq
aAk2nGUOs9Pl56BBVUYgipm9KkGE33bjyz9nqgnv4ewMKr59ibgRF2y8e72bC/GPqdz1oKCcdnIY
J4xg34NMs4KRxvV5GvYUZqloK6Q/qqo9rlt5pZ3UiEPuYFCbSEFr1RBYu83SrP9i8qZRC+VI8saD
IMYAXZDNHYKtKnTCiljyCYUvO5RJffXcKgxuWLTK2YlXVfsY0jPjrTSoKWRqKf11YbyBJ3nmAoxl
fMz2hp5tLE5Qx2PmskMgXGvYiDzj7ozRKLQa01VaNaOBCoxDqzbuR8sZMHVytMoqy2UV7pYhavF8
vhWGDbirudaosPMvwJrQAc+Wx5srnmkuOIuAGTYi3gZdZwUZbVUoN4w5hadBFcVXmeDU2GYDNibs
N6VfPdQKhFVZTmEcHBYBZMzwyFIUt8B4MXm1eMI0wD4p80BMoI4XVnOZIJr2ZoXc2+pXXPKjooRy
bFEDlqCGmdfgoc9b6DNaxAXDUTP4lYqcYsms+SdVoK4NCnU8JKkgMkd+PfvMb3mAFm7LdZd3VbxS
hxUMaRkpC9Xi9kJNux4WfNQzJnjDV3HpNeknByi0Z4G1CauHScwv2F7GtV+aE087ngL2aFtPMsaJ
2KpZ+LfWSP6cgrxdDwwNxZ6gRD96USALrf0pWDpm8skam10ymTWWk0m5rG060HUxLlWNMxYFap/T
LgzzrSNflXvOZfZRnMwPI21bXjl0BYbH73SLx26YvZh7Wl4xGihePndPqBUHiZALfxOLU6jmBSC1
kKhCtPFKi6idnBzRxE1rR6HWLO31Rr2nbacD3jIlLPeNpSy400fJiXaEcqiYEAzR7H+E/zSGDEwn
iLufWoeoLAkttMuxhGT+bovKJ9ydtpJCCwXgQpCEzYJfOyAtWrvi5tWU0L9fXhOASOpF5+w9YMwx
wLoEpLbnB4JGgqkp54pMvfdthpJFwWxaC/wT8ysBggGj4NGX4kyNvjzD5CcWjTUD2Svj49/9tNTG
XFWLuOQu6hXAjDlCEVNneUEAzizdasw5Az3ty/1a5mu0NJRoec8Dx8PEH8iVZ3Iv+IQHq1SKA2OH
SfOuByPbIAKmd9tYbphSeSHNxFz5M2Bq4mXeGQwEPUTk9gRmwJsOdzSlwASMnYh3EU6JuJoezjpC
nCUhMDpnqm9VFUL+yhvT1MNprs7KLS3GFMAOd7mr/KsqAJBEWny6Gycpk2MqyPem5auhxVk2mVLm
1gFQS5QeXMkrlw3jtJi47+uYQnlDwt2VZGt7bNMdHopqXOh/1rY2RGDPSqRdE6r7xPy3Nz0eyFty
SP7TVf1CqDguQJ7oJDaosSyW9JCgbE4HEz1W2p0DytOMTud5584G1LokM8rgeMuOja8+Ub2osNrm
iwxDuNf8DpU+9itfZ2B0HBkcTlvtiDjptEbq1vj40IQUUP5PmyeolG43l/DGfn1Q37XJooBGYI9k
n0WLFz8vbR+X9NRzOfSATgXE+mH93HG6h+VvDhYzSSFzVKIehxv+mT3Gj9lwKGJyahD95Oi748Lj
UzQNtWf/nJffrSi5aNPC+xppYb8JOUTp1PxgJJdATkBqxRlHt2sRXhKF/iyktuYDtX9lKe+/Tq8P
Vx2+6TWjfp7vkJHnn80If2+2RtQMkasoILs5fuAnsTLUnpOmnJTnvio9KR0DfKftW5kMCrIDG13n
SS98Bv9N+JWO7MeMx9WAqbzWfgX8N+EqYXZNRqfPdPzbnNn88pxy26lLm9P4QaNLL4AwB+8z73Ny
IzSOUQ93M1dvpgsn1mTv8yilmJwi6wEz2hwxcKU2Q8ZFHsRKYVvXxosYd9xK7T7k+aRpX38XzKrY
uOTKKTFU7DaBnDa4jXEPzTTZ7L9mbx2FvQUnh85FaAldkoeodZkFpbk7VY6CU6Bohf1rlubFcKAs
xc50aA1fDPsFzS+7SojkY7PhCG+8MOWJirp4PPUyvDp/ga/GsfA5/hTNG6Jxri7RyTT2dhnirnFj
cHawpjAASF8ViH3MsLwsnijUtknjNnYcH2WOsBU8EwPvRxJwQCyyuRAu0DAj2RT+tMpNSJw07yVQ
+sUMOgM8C0iv/V6c/eRDQkMqGxozrpX1NiNtjKJUDhv12U1IDOi6uAy3W0f8Q2d5/PuCmwhUTU/o
7eQnHiCJXgAyyPX81Kim5rNg5Qkvh9Qlw50s6yby7kcuFM87Qn90xzUHv9A1/yXf1FbZCYIJihsK
1q676fe9ihZjj1Za1vvAY0paXKtPBpvpCDLBwqIzfUoxMhXTl9HHEiJ7kp+wXSoUHN0xnIoZ6DJ/
0dPmzilOrwOv3cWyEs59eZ9pPdQvgvf4NgaLur/SfgcscTCpaA9a0TuC8d4VgH/Qpk1NuHL38+k+
O2gkpgdBJvCyiCqTSbjpd+9XfkLbypE2lxyv8uf+689y5m58o0ARgY1pzt4Qt3wE4Vbg6MBnqlny
5SfNs5Id0DnELymulcDwD3MH/nZN5a5E6xoMwkT4dLrU+uZT58syuaaZi+4guxi1zhhDoPie3OWZ
lBLEgWXyhkP7F30LTQGwQiEPwareu2clAKIByGVD73z+dGjkSFPQNG7RXFGGTDGMWFutcT/b/vWK
i94oRnA8gGyoOvx5OUf92m08VJTIS1LowjiO6NFXkpnZMDVfp+0Hig5PQ4gWfJH5AfO5jpK7TrVP
FkJVpj/NoufMoWP4sdb8XOpTCTwr+YsoVNfihatMcvwnUwLC6GWqSOboObUvZvfOqMH7Biqw3+yl
1f04q9PEnG5OFeBsS7D3csUqcObaZY7WkS04+6hdJuMU0PzjwOvl2KSY797aBHrUPG/RCr9pNB2S
FgSL3hNIiGfAuR+WWEYUt3u5PVxA0aAJz3zVRhiDI3Cj7QONUXOjA+zGx/QTGAQbwPplWqRCymOJ
HKN+YVFmQRrqmHzu9MtfKt8Az0OeqTulxu+StGAVPlhHHz4N3HP5fxZJR6kSPS0ECSKcGTY9acwO
Q3xMKXIL9gmhiy/seX6MN6bFOjDgx2Kk4VU6SLmFbJe/A7O5DRJcxCzSCGCWcE3O7JonnJqd8sHs
MfVG4jqO7r1PCxPRAQNcpBLdGiImWQqb/8vQw7NUYPUvxp4NjyqLHPIsHbj3qNDisqyNqg7BRi/F
vAtzWlhm5zU7v4rDfxHYbdsknlVrIALxCHE5fCnbRYVA+O2koxn7qoFtNvsB9OxXNJMd2c3/j/ie
3Tnqh9g7hnT0GOkQhbzqrKYx7XLGv1qic2swMZ5+lOyiSMEV3djA0cKizx3xYjR0d+I5ZpJWpFPn
fIr1WXGbNYCDjKk9+z3hCSw+aGRkg9VdIru8I4Se41g8GFRXr8nA7c0H27nLd6AfpMqAz/ETsGI6
xORzPOmHos+HYv57qxLs8Qcij3xxDH4KarU738di+QnEP++j9TonIuZTa8c5r/mdAl6J3/PCuGHE
FNwo2Wv6Tq/ehJLdaxubp1MjOjBrkJSdXcSNF29aCwLlmAjO5KDvFKiqtJhqzwnonv2tIkYBh8M0
NgRuyhPWj4UZ4nVsSm1ntbpwLDEw0mbzLmDTfppb2g883Yemm6bzKfOjK9Pwl9pNYRmLtme8IXzt
xVA0/4FZbCtjSOq7AqF9liMaQLs5aGELTJ/MjaWEgpnBeJMhCvqEp2F+PYmNIpdjMevG/99Ppnjc
y8tq6Tlo0z19XnIMblCeSxwIdhGXVfvD3PifbI0M00cabeE2LQ0a1sySFMt1x0hqumSLCd3/qvQk
OYRDIGPzAq36CizfqHridUgpC3jCxS+bkM3EaVxBo9WYrBOXoCm2lD3Jf/dUd3jUM+UpJujhc80i
SPszlSYD2UOGSHY9KAptm9+ioWztFAjHiLOJK/MlZ6F+/LvvE7Cw9zggkMjJH0WgE9JZl8PGoj7l
U6rXSLwZsBGHgxDL1RvcCeNtXcNHy54Q6pe/DP63B4aRWOQFcJu1C28glTAkUJVv96mGsr8dDsl9
wSrrOuGR+LiZmYGdBmivj5M+5XJiI1tz4VR9QRHE/qqKkXYEbqHKFyGtbWd1NUgVC4Tb1Kx35GCc
CqpBoXcrpz+sA74qmU9cN+6k0Eg3REm4g9MLXwAeQoEX02ER9pSVpSYYedRiv0kTR24LnzwnuGok
uii85mDNQaKil2PCsRvEc8s0OXmdPhZSYBzfLUR0jjjOhHDU3uT/PiGZ5LcEJ3prYgyq2JQ6bCd3
cKcCX/5jYxYCa9kaPgn7jjGJM6eZR2U4Up8piWrRzgNt2b4XNlM/FcZL7KF4SfYpCGTW7DiWJPBX
4V6SMHFfzKG0lLbTl4prnmE7m2wsri4m8wPoKbwyPLqzF29mhRrqpFGeB9gyOtPaestfhe76FRk/
fMeNZyglp0RfgMVG6cXSHzcrpAmt6no6wA2pMO6tO6gVwCfWxCjGbeMuu2CCTTdBrMvhPQ9XrlUs
tgsGO5rQK3ggZ7NQSS4K3ud0hy2Jk6I6DKFmdQRed1CxwSNd9ynD+M+8LqtqUu+IR5jhko9PZ+Ym
aMSe2Qz2KxyLlqpQb343C0xqsJyAYdIhWX3Za/5wuLBoxWnWmMNxRGuvTKrS/2QPnQ3wEieKy2wv
8/Kc9VKBUMmqdu/G1K+dmgmgLYNnRXJL7TV0efKsvh2JhTTnLCHvr2pe0s/gE6iOA1El3QRckKYD
j0uwPk84diAb/gqfJE2XZsiJ2cTcSpA6BVj5KL3+qFpa/qEccPOeVyb0pX/4QR/6mJTODNHihcKU
6+F5WLXZmzjmYbXuqiFanqHHsjKS+YL+T7IaSR0tARfxkYAJ2cDHMGgSWpkd0wlfQFEeB48FApia
Y+WdZms1ch0H9IBrBVkBCi1MN2g764HdHWNgWJ4V9BW6MEW/qKBlE/hIa7C9XE5PDEBMGZr66UxP
RTTAS8SV9eP+EPRoiYypE1bkDcy5/+xOrC3Ppi3CvVyUF++38qvq5E0kST+z7v/RgS9v/cJgAlOW
WJBMRKdxIXbPPxl9nLVztBaTzzfdCTN5LUQpbd4Z5I95s5zgM7kn4yIBtIVL7ooA565ncOIyQEkN
TRo5NArtrUGyL65EX0vRi5ewCtXYmgwmPW+T4/qjHHGkYWffJXIiVdRerx3q6Kxv8Mmk+eL5t0ei
YFkeCgdcPIYtYPZwlVqRDJfPAUK/Zez0HEilzpOTpTrYkNtcu+P4TBB2cAckrWl0JtWvXbeDRbZ4
0xdx862U6thJLPPCSJerc1D1xIFaPdCPoo374WBKMTIXZ8KiwJ4IdyVFE9PFGBW5fuX7bpH7wC18
9ACJ48FzOHjLBscb0zjg+j94T6bouOAYcvb1KbcZViRLQKq4x7hRU+Kar+CIvPZRRlK6jd3P6wKG
/xZIjmChsNCE1rVGfag2aLOoaXtPf105lc51SBLSJCCsRBh+YYMm1pejgJeLX0ALwo/g2Lq6AUNS
8paT6fMz/GYeoQOAaZ7rNIO794HH3g+Iw4yTKFksIpI1KeBQvJf8CogW+KE1f46V5QdZQt+4tfHZ
3TaxSfAGQnpeHg5p1MA0knEqUxF6cCNUeRM+P4KJtkjv4QY09CdCGEz7HLTEPcg6DXFn3cWwjGob
gFn2TL5eT7UbMSQK4kEJ9OVcjw50y0/EfNudBVZRwrLJLOBj8OjNSJQKKedaBMFYSOgVXvZiv2Ec
N8g2bFkxxCo52A5qwnRWUJKI4pcQaeP0Qd2yKrS22NKZjrNSrrRbZWDeUhe5Fu+ZPfFN60/85O5H
O3ZNoY81TnSXe0DNjOmCMycpJQPkFlYEVEnjcJrI1toFpLtw5/MMSkR0m8byuIml27vzJAPAabte
VMPWrb3MrR7QHhDZfhDVsDk1job3YE6i69XhS2dJIuE+NZomznctKZPaY9oFvjk7WccsCuUdFSWB
vrV44+C3os7A1i1ivpmgsv0mjmgmTPDDbzH2uwZHHVLVoZtALw74JX68yqZsL2y1RAkOLxqcjX+Q
+LEMSmUUtY0+/B2k6qrnovkKZBvhvQbT4NNa1f/otSK8tAPZ8nhrHjb3mYhCTCDwterOaKwvBOEj
Ws0WNr5/bDPCrt+pDSshbYyqoTsfD3l8mda6kQaBNP5H/x2OvToAdZLFe5eLzL5SVh9wNldtlm0k
2fK3aYwgkf9kHIjIvE1JZVKh2meeGXB6/Z/rq3dK1k0hFJsRYYNekNtIgPDIY8moVhOt3b1lz7Kt
uci35K4j/JHoUwhryU/oa2wPc/VRp8tITQVC7ziOyXGt7pLJMBxCgTb0HXnabLnG9yJo2WTYVW33
9DAqDko0V8GHrBbs4c4tt1jMUSZedEf4hbOhp6bavZ3B/1kb53skS6douALUQZBZA1XsyHXhVjAc
22A4kB3P79/uGYtHk26L5T3ZkXBzYf4HDGVB+Xd9wxz2XUtb7q0ADJnnMiiBmI9tGUfsHlD7dPsk
wlsYCP0IM42ix4ZnL2pIG/sEsEpa920Ajfr/AIzvkqLYGo+jgI3oit+CLKKaM0wzetT57Pb8DYMK
ziY70FbcitoeWvgq1VT/rWQo6m8WE4CNXcFA0Ib2a93g/6Ot7YIBblLV+DxTE/lZuUTA1UNK1Gu7
3XzQFmd6V99VF9dUV+QB0trZlSyr0crA73ag0ex+uTskqQVVl2+oaWQ1OmXNANbPWk2nIn6GGXAi
ZEPpr1Ssmshc7nEfdaatVcWnuA/NkgmOUDjldX6tOSHmLEzYtW80uxmQtZXSH/qU7NaG2AnJ5lJ/
tFkoXBqYRidgSohq4aos/wO16bTa3anGnUiqRdsoLBLXIqvsZWFOcBObgtzDxwkPxzf36fwQuVI4
lChmlIneBds8QQ6uu0CSb6lhubgDEw/3Kczj6N3Yb/Sb73VWdqP+Kyc9iN24zHtpV9hod/wrGL2S
ZEcCMBPw1sHdNRmTGmXs96o/SH9R4p4ZGpWGUKG0zbAx/mqkpc99UFXm8CgUJUqX8Os7En/YlNNS
HZ8pJ2Rj84y91C1sWv8g7iIIwBhgOyPyB3wAHIchpdgTVggKLrsCJ5/l2ieJ/88EESMFawpKZzkz
prxqiRZtI/4pdWhJxjlL7xmpqu+uFYmdI8eK54oQJvB4hMXfPYFCgcM4vttcDo0YUm18S6ChW9QF
JSjvdrtjKBu8lxf9qJIy0mIISJtW3030MlzHI43+Gl8HygQzDuvQB51AwJ/2F1YF7VJuWpfkP1Ni
YZNy3BXCHMweHCK/fnGDox95FEeMuZv3Kdyr750790TCo8b2PU7zr/VW+ACTaqyU6sxnbx4XOmI9
XFIndQcYwEIeZ9mXfc+jf7YoKc6K1qhiAmCOIUh0LsIsN+a+S1juJhEpLwv2pUI+mhF6PysXdQM1
jmIKJ9rLPLAPCJ+u7qUKdPCF35AbeEwTlqi4/7RimwYaxlSJr1PrqVzL/1N3ktXZJ7Z4ti8kBndX
fXWL5BZbmRQprcILDdP+uKRPA86XUQFL8AkLDPi7R6OOTQGcrbY6YQiju8OhuuEfk1O+J4PuSKN7
yZrf0BJShaGhFJWv6ohcdNn3CKyd9s6yxYpz8ACMZsP77ukPVWF6Z35cCyJt87BIfG+fCjEgTM0Q
RxQ+pGicb9imgmHPODPskevy4bIvIFSgyPbr9N9S62HngnpbWp95QGGaltUoQfAqqzWjXBegzJ4x
+wQ743/ecVmFTo98vuaK0nuzcZhhHrzm29V2/2tfFjij6ZrdvIyrcuXu0AVkoDw8WElgPkfB5EVu
jqQczREnW9Tr8Zo353KdYYvGZqWtWnHogL4aOnmx3Okl0PjEMS0RFDSaveIRo1ErpHEUuvtpPFGl
Q07cvrVYy6J6iQ51m69oyRQyv6xFWqZ9Xvxpe0bwkSAdYzF+rzPwU7ZaT2nOsOQI8gEaDbW3Ghvj
RIXBBl4SC9369+FQFnp1Fa1E4g1rkVstgUOfxGMjsyuWmDSiaDd5cdaRDqcgQjrlSdJ4yUa43mEI
e/koB3HyWlpIkg86GIGJEdarY3hmcAG267MLecX5xebB15m38BNwF+VhpbiqjzFCQJe84uNSuSNk
ZF68sEXCYjFDKek6fVJwuN133Oqd6a8HJheG2q5+zNQVyPUr++fxn8I7bYhqyLAKV+5ERDmIf4OA
lGHQ0rsK+NgIovkqINWN16JawPpA+dsUID2qAaR2u4YonNqaq0MVVSChEq1NrrFgh1ZcYJx18F1d
beh+tOKbRCqVv3jQCxXDEpc6Ez4At7HEmlkWtZ8AESv0qdY3ZSCa3Kp20DAtOVvhU1wFFaq5xxKj
g6FD5aIpgx/0jU74ivc01QfwRWXUJWuhxhWsZu4DW9lQa1ZtWYIlUv+GnjumLRa4kUfP35c28t6q
g+6HP9njP4VwouoAX6AikYiNh1KQk3FKknZQ7+5IAvrK+s5HEvBxXIFr8TLlCFCe2mQLSJ43oh32
xd26CKv3wkE1SjPzQc0SKJiRQ8ZYNA/BWK3dwZKGIzgeBPYyQzcaqk6t0WQ+huFrxuBYER2Zo+MC
AopNtN1lfEJSM02xRFGU/UJ1EbielJ2Ryq3caXYWl8sEPqu2HclfAVxs/cTHX/QLf5wDctl3smUv
FDfiu8OQLmSnPbsdFWRPc4U+eHb5oURo5pKWgT+c2EsGuBys/lBCFUexcY71X70FWBpKXQGBvsuj
sBCViBqvRvlJ0+4VjoHnf78mOqTHWl9PR5U7hZv4quFZWq+6cXUwzKBi6uaUkGfwF0qlZ0gLnoIq
+P/OZ2wT6HkHaVMav44htnGDKxq0M24yJAX1J/sNqATCLSJOLZ2ocvpfMKy1EukzJmpcsv+EJ5oK
hlqeZOa8xPaTWVTyk1C4KxjzKLgb360kuzCJiQ4bOHby9MEPEN13eHAStJ5QfraiI7PjYU+Z/yw2
vp5/jynwi3t2FtHP5VaydlB5RIUXYbSthQJ4aVZXQrLyebZlaQxBs0mVecb6+OUj/Lj+EpJSVKg8
FaGXDlz+t7Xm0BLjc8dsiSuCdyeFEXzTGaPE4fNoe4HwTNh2m719r3bMRfAkaLuyTiLhG6+x+cEA
VXqU6DFwHAXbyfzbCoM7fSRHHdLn2CL+S1pDFkBKVXgL3kSf9DPDEf1azvLqbKt3RSerItweUWyK
gv+W2suqAHUmn4mSRC4Q8OTQZ5o6YhipsaVAjSCUPPyPMmyR6TpKbgdHne0Cfiu5bgxXhH8TPM+g
BcrnUgck+YyyB5TPtIPl5FJdxgUi6XUZOwC8MwwLg4HznnCCk4d0obny3K1+1b6lHJszV6TvMk8e
XTZkZwkYQD0UtPNEucXQN5jlyEy+Q12OlOKX9SsewlCBNvyzhAwG/ogTspbkYCJ8Vuy1EB33X9pc
IntLnfTlAxBdKqS6V85bbaF5PWg+ZwHT/eVe9pi8tJNsElv68eAnct78Q97yQCXVO9Wisk1Zj85E
IFRtzKCm/uVEqNQpwy4v2nYJ8tqUCY4sCQ8/tHF7bOEI1J7nvEmDA0gAOzjty964qq0pESqcWlJc
mzS0p7sU/Loj2mkCDqIY3JIC9Z20evY5fXMVLHFyQ67m6e3cvDR4RqxFF+i8Vl3NTKvc2wN4Eh4G
9ipQgv/84Yu4PTr0V4UNM/zMTO/4pj3d1coTnBlT89KerdQdHeQVb3JIOjJnJ/xuKzZS0vnIhpfl
sQOPYzpjFbdkd4Ut88RYCUBwlQ95Nc/hbVKMZSdU0lwcJwpLVQS+VIXYgOaQOXkHu3gXGEVClAki
GiNv3bU+iw38EGg5lvqiwnHFSltWdGHpxU6pcYGYPpJIXRfI/itx4d7vGkDFA8JEMkFyvXI+0GgE
YgT0xgG2PaM4OL+Hcr8TCmKljQI2sGGiMios+L+NkV2iAvJbKHBZNQgFqBgIyeRGGVmGhHhNg+iZ
5o/XiWN5suV4beUAagwcmoxCm2Cv97E9kNfAhCZ/+U+3J98qIOYkn+mKEZmMNQwVh07zmWBwm4vK
51JPA/Bydu8Xwde0nvS0GFEEWZ1psp3hXZPdvQT60jqgQl42xBz0ZgIEbR8DMy5Cq/1nDHsfBR5v
mCrP6rgaboDU2KBKHfVl0hErtj1iq1fJu1k5qH+BAPwmmkqF7uA+dfl2UcTu/qS/enr34fDgljJA
AZdQoyQgxHPCsjc62f385ExAXYIOts2HDY5T51y0hybz93kHwiB5ahL3HPbacvXAaZPP9HWo14zp
/EjGXhKcYqj8eAlfbLwXN6sIKU3UsvWVRY+zedcQG848P1dE2vvmApYq491BQJTENBTEl6oyp325
6L5VtNjqz1p+DorIcEoWl7bsEmPeGaEME36CahvpV8RuJ43/6BJ5F7VMtBQneFOSsZklGajJuBzh
gx/iaGTmrvNpkXmWPeXNXafbPFhQ0ivpotKTZJt5XFCnc4H3kWc6tBJSd3he0GEBk+2VgheVON8F
bhtSXrV2p/50wJmdvwNSr/ZQFSBocGd7JlwHwSZoKUjA5oBKrno2iuie5lP0+vsEF7IHMWGG0kxq
NodEGTonL1bg1/2BfYpCpgx7Q3sMyM4FiTnViEj/mUPCsSkY1IAqJOXP/HTvbH1lb1qqoDpuKvCK
HgrLIX8lVTPTUlEcrm+jiONG3AD06nzOQ3HcxgY5vPSW6lfRbV0NDsbPFeWYOgJfRXEg4dXs8j6E
rVMo8u38ZHh0GdJq/l5NRInHFxbiY++eVHPEXKBpbx6EhErAtrHbFjafs5VCi3428B3WfrMHagYJ
OhL6ng0lLFw2J8c6TR9h+1sxRlCPRZ3fvG/HQ109pK+kRpdvvzJTdx6AcJOHeUIsVW/lQsgc2Fkd
D8xuXkzvblPXeo8cFedJdiGK9FGa8uY57PHZisfaRR8UViz14Zy2Xrq1hBtxnaq30Hf1dRAKXP1p
0WbA8NZ7mBkjOR/ofM2kgfKbDNIf3rWH44W+k6TxU6ELzJtcrqS871FD6AVQa9dK2ldRFgXEPhu5
+KgRjBjwm1bpSN6v6nOqGswr+neM8wxsTNA/k0Adve2m6grKb+2f/4azhl2TUB2XjV/qjck315Qb
yRhE3tTFwC6CZ13veEPyZQUkH7XBAtSrgBwVHSut80IdfyyHXK6T4KqCAbhkp24btAy6jeWQLc8v
mMN/emoK3qykZWxd+tv+RpfgpUSGMDmcrlZm//x7+KrAjh9fwyPJtAzd7J75SA6eOt33Nx10JV6e
5uU6sBSIu/71ivr3Eo3iyREERbAnykoazePIJ9kxzb36cYoO1nRWROOV17wzemvYA3yu6YP2C8V5
DwvxI5Mp9rHYfFjKjyrsVmjDJCU8nkKPFOb5j+ue+PzDlKTzxzDUHtULcKGY8IymE+TgFHXkyEPL
DwL9ymXZV4KUtIMD8rpWIw90FbJbasH+7iZVUYYW7VsxnjIIi2pB1/M+fyPfCZfqF/DQKzQ3yC4I
ipHgF0uWM7UBcsAhvSlnYxa8DOiQZVBD4OAUDxiYCE5CI+W9dw0K4QNP4Cq7NR4VpPEW5aW0gk7u
jU46NvkxEkCkWF45Bo7bPoIpWcLc20iR9vZYOGmvD01fBN4osZYIyRZYY0L0n//yKv9Zk+IV5poO
O4BuKpD8pwt2mYSg2aIjXvivIlTDZ/bQ1IPFooETRzaEI5jqVIDIcwhYT48IDLAizzxv4ird3FsJ
zi6TeANmSD5WSnAetvay0+tYmqV/cd6VdxyTMIayBogvWXNDIq0WBEofeXWU9B/q8bGJEEH91PJu
0z0N3Yfh8DHVfQTryNbCEKZvljpOI4OwwCdUAeNtks4LTk8WZpUhIhO+5Qd32Ilihkl89aSH/97x
Mvaec6Pb2mZ7PrlY1jrxOJH4pf0JFavJ/l15DTXZHjEmaNeSO1VZ34ul74BnQtAeSvx+lTlDjsjl
i72Ii2kmiThdMw38pJpOEbaVpOHCiCpdJu5pfqYI6gbe9sHBfsNFtgOOF01bv0Y0K8Dr37PXo9O5
qvdIJ/dP0xrirTVAPxS1lyyX2w8n130MR/hKr6Cyjls3VR19HcRvXfoCna7fmBGiaXxvsd1+5b22
1T//AZxjEaxqmPmAM/a8iKrzGLdKd6s5VXGiJkpK6r2Y9TI4Ki/8X3JNB4985l+r5B2xURkPGeNj
jmn7HxdL5Jc68OBevsrqzWeeL1yCFEtBRNY3nvtWizBenz97MrPbfYj8d1PtNSk/vXvQz+K+MWbk
x4ZqYNf75uCTPcGAHmwHQrW2ar9KNsxmRCyycTsvWkiclMmGbiOh0mSMk1PgmRyO0DYcPt9UEVzU
ByBE1+D6IaWa+G7Rs6mI+DI/mX6SraBkKWJbZd4F5+loDa5MqtbVvagZ4y/cXvi69RxWXTKxgTia
Z5FG3DUsDXsTWpuMtVlbHsTwDMthczWYj5bfRxbOuNIcJSeD6mSPRNsVhvH2+c/ljcnAfOXuhW9w
hMmpBX92L4HK3xOw3QTHHlMz6emrAhKGEiPLU9xXOK2S/8tnnI4ksGf0NUpZH+BBiPhHkQnL8XuU
OXTrCYkev9KfgIIQvLNofBdQnB9tV0dilLuSTzZjfEH5NHFYfj+W32pEtdULSkZiYIlnRZjoVB0l
HA/iT84CnOaUD6hto+LowUirOGu4rwr/wQXqs7VnJaZtLnvxbTc1Xd/L9E++GUhCKDactcyT8Ovq
UtBpHsO0Bw+71ZCJhI35VpvgIQ9GYqcx5g+TOl8X05FvvYZx+tEKUibtQa16yp/8NwwPfvdtD+UJ
1xCfXr1yy6RIJMqAlf5JXmMvB/AUddp4FVNU7l/GCJ3wwuZmh8BgyClSvy/2ScmIoDNhvAgCEZeR
czNzppI1+JDGzXO+8ql2N9sXIS1+0EIl3IMWi8nQTkdBcGDMn4Qr/T+ufcZCdf7bCN2Phg0L05h1
gbQop8TDWHp6e80i33JbpsEzmjubxJkSHAgleUPGFSerd96/eHLk62z+5QEtFNAEBxT1ALLwgNRB
ed9R5kZPHP68qa07Qx6+f1bFomKmEHJtBvrZUkv6Mkal/4gwCnhHoYNELkvlZ/3kmV7R5qo96KEF
Gao6URzsUIs28t+Iz5ubSDpFpZiSHhHwdM8NHo5Cqke9gxxINL6EaC5iHSFC0vMKE59HIh7Yc4mz
kEMdJAnGuy/yqPsLjnNtZlf5OfsPyw17KzJ4zyxao6tEt4DbeqNMsQgPHr06cjPZWO2LvjnjGtF3
Bpy4SRfkTEs9jXGZC7bhOut/op8n7TAtE1zsXCUB+FVuiQpe01nkgePm96wZMrDN2JTOMjXpeqsB
R0VZqhkYZUbOLpFH0PvpUxxAhDB6VRaap6aN4/MKTE3Yv24Mr1QAczdBMwH/Ylypoq05TPeIPMhU
O/eWda0RgOGl3tsEOAue3gycAQ4mtNRZAhAZUNHvFgjchzcPQIWmtDcz+rIC3kun8D/5jByri+i7
dmoCANJX+b5Vwl19vmQfi7Cwb+NsYU+1iEzG4x3pA2fCxj7C18IOfYxXCQFiX2A9Ucp2GmH3NHVA
HN9Pir3QpKWkIbKRvpu5YmCWAVJSRTqQ6f7xBHkI/MhsrwRH5rG9JNYRixxKl1Bx1osDSo2Vsmy9
YQK5KRLFVb3go0wIfrmvchPxlwdybW+5jhI9x9PIjaUbzeorteWrJGmDF1CVeF0RkiN+IlFaHbpt
JBR6Fcqdk4Z/AiE48YMJeyMhEwpVcPA3lZsWh9SKLaUhtYAYGUIO4R9NY6uyVhMj613J9we9jqjc
98PTPHdepKrplur/a1B2TECCszpHs5WdeEXglcKq++0TOYz0Wxg13DxZEv/wgUwJd92vrizSaHpY
Uf6jWXkyhSBxulkp91jlzWhoxki+J94eSiyQospVa73tg0k+3DSO8/Ssc5Ezh9MgY+h53cvhlRZX
l/k1Pfqx692V6MO338f9NqDKF7KTwuwgK+W07EUC9U3BZW024YF1Y0TadnGoMLKC3zrLCdrPfWFE
knTDu5F2hkeij6v43Wplb+jH78F1IFFv2g8+1BxJHgIZBdVOpkrCy8k6oeJyeRno3QOYDRK4atvR
+/0XeTSpYtZ+9vzF9Lj+vZx+TDaFpdigvNu447vdOxsF4g6oAgYEeJEcuo3osuKQ9iSQTUPqb6M6
ZJFISccyYU95D80YkJl42Wzq6Ojy65hQKVvDYzxrcgtLKXLmQ5KuHm95XFtvuJlY/1BaN+MeP6gb
OjULGjmAJkHLA8tj8cYYyFIteFH+zYMgVuc78i/z7LXEdfu1K6fxf5IQPkj/iLQ1l5ZzwC7Hx34P
c0Q9QF2BGgmdAeTjwyG2NGwPHqQCBtcxgy5gdzvgWTeVz9bLsbxatMzlFxP7B6dUtzdViHbqJHz0
v+cVp9BeqkZIOQOedMrAe31PoLgxJYdJblmQ2kDuePVX0lblDEglXu1nXz+DJETedORS9Zz4xugK
H+H0qb3TzlcFuRQnyrPMOn70rQMsztwOuv/D+xA8UQJEnaX1P++xmuA8e12k11BdqAaVeUE/pB/7
TBIdkjhTX39D1XiGcO5HVk+at7/WuJ2Q/r2lZd73wkPSDPZ7xRNckjCOaEqkF+B+bJMThU9nkn8l
5XTTGG3dED8lRgJIiIksUpJLuk4RFavfuQCYbvzvG3yzcq8MCeNIWoiRoaIYrhC4jf8dKIcV+YJl
dj35oJJ3b2r5H0zBYbK58oRf87bt7bW9qa4XiDWwjQFAIq6/WTiunZ8RmN7fTe25YG3YSdnxWWtL
fm7gwx7bvMNQKp/13e8I9T/UZAg+9Mhdk2v2WkYpTwHWIVWdhocavauBe5pCFVvb4tZGPpbdHnsV
tv7CquOcIQrjVWI86cUAzNyrE4+G/f6FR3l+hyxNGWaAPglndU0LVKBTOv3BpCnkwE4c+1glh1OJ
hkhY+YvYK10W2ywZWu1CFT2R1Pf6cnAQJHHQ8kugMLn/J6hOVcbyIYtIdRg4ypexy6X4IjTu0Gqq
Mi5aC8QvqG7IX/IzQXgfpIRkn+7Hb/D/WMMA8uaBUdutz3AmJelLiyqDFVxwzczc2OlWYvMSlCBn
P0PrnZgV/wvKGCoXewbFxrdlyNuN9WSnE9Zfl5X4Ce/K2Yanu5UqocmKc5VawinEbsdIFHCnw5ES
9V4muXGhtKQf6TGJf4MvBGzj6P0OhcpsE120dKnRA+KmVobFcpMbd3Li/PCpIifWYfCar56W69t9
WDbhHN0GSIBgJ6eRqK8hl4ExOIBjYAaug58bw4rqoxpWLnrh5hv5I4gp1Kgrez15oJg9gW0G82l7
0wg5Ml1KMNFweFhjYtaznQQiQJpf3vC4sbbb36W68WonEAv0cz5a/t+nOApMr2TVZqFDSUPbtlvI
huWHEcsjJeIkNPlfsyQXMqAvAYXheFs3HPkxHYpGnswUmzTQOe9qPtChOBUAR++kiK5QnT6pSe9q
FnUPryVL2oo5VXn4FS+hgCPQNaZHVE4oik5pib6BZRGFpc/ZLWT14UFl3S/Yrd/Zp1qX203bLMZ7
atK2zcuZtFD2ZGUES6P1duwSN7tA3flLHRUHmhfmNiFPIv/VkGHiWZ8hdNLcsFlAZUkuiggVAsiO
ZLxdUvXxgr5GfIEg4ov4WbA2dExbhQ90FKZy8caUAMefhjxArs38jGyV1FfYkfarzrKImDG1xhj/
1tsOv0dOVTllAzlVOQYcJZUbDdCroJIT6StdbRs4QTyiZ76fUuB7lXiA+fXlYGoQlxYIxr88fCXK
DXBpx8eAt0KM/CY/r2Rm2sxAxCh+W1uHwyG65px6oLxFBaTeipymd+81qNRSuqUYONVzlSjW/RKJ
IjYbGYzkA99L9d7pFaUzadT/5AFxB8NqH5/An+OXPI/EhQuXi3YWUWe2e4ySfbfsucWsfOS2Gl8W
WNvi4GGxCXr/ImkKeq1j/A0JWF0CI4NA2lzlHD1jJoTJO0/RAnesBEl8X4tvia5yVJ8n4KX3ZwO4
H+CIuXDvJD//tvnUpI1r333iEFbeBCPY0w+J5me93Jtj6ZBZqy2o4wjGQpkmMHbkwwkfN4TjodDn
S9UufX6SX2momZx8uRFmIGkCMP1ag8qPr0syTF7IYTU2Z2o79j6wfSTDISdVT0tYtjWyTX7NTZ5R
J4GPqpCPTAaYQrNJ9RzO/kiyuaAv11vzi1o8L5X+d6EJcG/6/NhXpkPs8yQCB0cj8WMHpBkQdGY0
/FbafsUEfi0joLqAYG7MvhwAdpQrfBd0WXG/Ue1KXoW1YVvbjYyml5ConqtPuYoHFXQQE+KTq3yL
Q+FXw0l4kVlu2gk3Dc6RqT1EVuvxoX9NnC1HOyE0kjU69QyS5G7f0qSXOwp9Z3ugodZzMozyrHZL
N2HtdUGZbnnimDPhO+SQB8+0usclnWzdyNlgycLSTakT5AKy3x+jhNudKe64ZT95Q4DtLBKdrGFj
rsp38H879lBxM89pXjFLaSoKBfj08DN9jolsJMXI1a/3mv8sHsuNrQEXg7d1EFzYhjxPek5K6/jN
738Ckn4t07WnXx9u6431aVj+tBOlxP/nmb1hFDW44IGmq4/Y5z3UGC9u7SUM3uckXiq3qmlLryjh
qJiDa2bWZyQby2c3ZsKNelrl8AMoOV/SNC/MlC37P1qGNv5KFOQL6L//xlXj7FWbFNEO4j0iXw2w
BBMQUgIvpTQkUDFp1swzBg4UX5gZVi660g75Ss15Jo+GOnrxi5jo7UGvZFncjrcB2r0NgxMmV9Ie
iEc7jXBn64uqHPN1RZpnL77pB0QNgFgGaodCGyuUZpDGUR3j0q+WvPpH2hXgQqMjEQjMZXW1HnRu
Db6oFRgP1R/HUSj7Zy+GOniuOaT6fvcEDKk+lgS3nMgm/PN8wieVuvYtHasOaJBNOI0KNlVgJp7/
ibXD3x49LmI/2VH95r8/U4LSK0wZzGqudgAzurBpyvQOM3I6heEfFPa7sUtbdBddi1S5Hvv4KtDU
HwHJWl2h8vJbDEVq8eLjCbA0s5rIwj8xJ9Cbh1Fs4ARdk2GPrZZldeys+/QQp4LxlaBbBv3fd5gh
aJaWgO0yiolgO9jYVgyaY55ka9qI+sq41XYLNl1XNkuLrnaKiEvuQL9Vzux6le+9fEwu2+P3PaHM
13WYRXkx98Kjccmj412wRtcQnPYwcCWvvjuHYmi5RipMo6Gdwtxg+t7RNb8N/6mnuwOWQalpRdbL
BLMhBBQPhcjzAScl6oEL3AgO3xIjubfdzDnQy0tOjaom70wVdScBIdtXOr9cm2CusxJGtJEbpb5G
hrH7DJbnk1hHgcc4+oah4XbMvsMtwyr9UCAr39ZWGUiKokaFP+dN1gQYfRj/FeMKLAOD/yxqebza
s487t9K1+hsRDavlOeKr8mpWwJZPI6to7BKXk9DQPfsXayn6yJ7uTjgOjm+Pd3aNcG/ozG2LaV9P
dGTDVfoWL2sOm7+isMfVfNuq2Dz/l8QfrEJZEscZgujUHZuXdLUIvz0w6KlsoSipC7SF/KqtIIDg
Gs4PyynJMe3u9ON7RUkF0YkiYcm0+JAu70405Lspq4N2OIBbHBAcnhCGuONAgA/1x2rJcMXFV4Ev
xISXVMA/3wxSGbx/w3BIUvEOO44aiJZk1RVxo6rixeoPUMWDf8lL0rToqJBgBtsyHRFAQ9GpFugM
nqqLVa3FsHm/xKx0KMRKEBGBoHwu139JP4X0xfhGoq5cZt+PabWki66ooPJ3QPYexUraNDeDhXk5
2HHO6vIT9a+vVnk+EMTGwO4NL4A1Fk/7YG4LJrHK5R5dG8S+yrGxx5vy+Yir3C28YvDnDGlPa3I+
8tsAAOrMGppSGus+ZKp3YrKennP5xCquaR1JUAu0tfUQMCaHfvgpxouY+UEAywHE68rwbpIXhubw
/i0FD8IfuC97luf6m91Enpr30uW9AoGttSYxUM0lDGg66qwXxE8NxQFwSVhkwMp4BvlflPGmgTt9
9pAa9dUr/l6VQDfKY1YzJdvl2XOqWyDDsw5xd03fX6nhQi8LBeHzMN66QwgZ/kRrzuhKFOetcxWi
9677UZkyWIZCDfRo7zEs2Eq4QGqUm3P2fCzN2JBaBdjXBPNBKAinnCCRLhdIDBjHxxzdaccLzOc8
2O/184rNlxD4tuFV53WA2+beFRmaacsGm/Qp5TaOCdPKNBOUFILfIPUehRc+aJjRlBOjEmChGf1O
vR60CvnzzF9CGNYYsQ70+ic5JQnzQPQnRCkgsPoh1pxNXOmU2T/q0yeUrFUxloFz6da1ZdUNbiZ4
zuZEASkSKx969nAO6TJ2RtcTaCIwaqL2v7w7z/W1KoRpTM/W9MglbU/VAnNWXOQ9Ju86okLpYF+E
EDxewl5Emh0d1BY5Uv2+aLwAS6KtJXCq9WzsvPJKPo6tJ3JYInLGFmv2OfMI/LY8c9ghyvEuHx7l
tLdqKSGZuT6jPMuCIOMGGkRqO+xP5JCNHvY4Iqco9jSTAmFhPmXuWtbrdAhBQV6sH3IdfTFeIoL2
vOxSQyML9GNvec4MGteShDfeF/wyrVthoIxvnbTcc0TJIWcuSW5SJW6wU1pT1tmoacxzK51r6hl8
txsI4E5h1qjWVhuMKTlFFOXQfM004mZmPGZ5R6JxoMDcFHECsLK41o2mTYuFad2aUBO/dMlorclW
6Rhi5B9fzrIhoQ2sWT0Ib0nE1T2iaNaZufvQzak/aIjQ2LcAA9G9mHhEKXHj4G0x/JX7cmcAZEqL
Qp9IhVBGf7GZ8OdlGjW0262xt+Qc206y70Hafs/fTBi4JHPH3SThal045XEsefzekMxkn386aswv
r/WcxC3X1TyV5bH+dKkLlMD1XGeFlmNTB4UDjwLQNLBfS17ZkbwS7dOpyKwiR7chcl+XsqtQGoZ2
03vtnG/IoG9Snviysx2jUSN+IK2Hn4nAOKmBHSgRJExE+P6FgEZigQzkWqYJJHX9ENkPOhS4mrlt
088Ey84tZxWWudRjOxLUHGySDf8GULLDfmJZNwvu+Q9kmoFtdcqcmaeDirhHAikqzsauw+VMOTyG
+gB1Mm7HGvpx91huLoO0xNFzHXgIzsQj8uzJhCVu5tDUnV8PryakF61OytLz9F1goumu21ZX5OOx
QWAIAXLR4SCrLdqk+0mRXsIlzRKGWWNddlZZyxjCbQfkkucfwAwsz+OYUnef0hWCxnMLbQxxvDSH
9EZCJ+El8zOYK4PYTVz2e1K92QNob6WFj8nzWMRfa+fCQkJkUZoHN5RDzvN9IgCJks+oVl5tL9DQ
UZQ9Z+SUIjiiom/hjDp03j2F5GTf5vSnGwNjc4i2P55iuvc9C1HFqe+Kq5TKCP1XKNIXh/cynGKL
Nv9tZzt9tv0e3/49Xl39vQt9zO1Z/LVSA6hw7FXOHcxXEbh9C0khk7iNW7GUJFmDxArJqrC4etHD
piG6h+olsh7hCxbt7ZEqGa3uoGfenEfhxndbPNzTlybMeOG+LZH7gzBgNm6/U7j66Wd4gP5vQG7K
VR6CtWERQpuEgoCMf1KaES1lk8OCsOidBpm/2M7cW/YmffL3hnxssBNS2izI7L03lrwuV6obguA2
y3mh0glSXlewKgHL6FCPS29JXD//FDQ8edtj9F8xzc1XM2UZTluICfG5Ax9Jbf56LkErJHtjYHJB
rhnSi4pBW6okIwfDpkK7k4I0ELYX6d+uEgETXmWTjrYsS0+WOJi+UfB0BCg19X3ce3MqXNWLQ3zb
7siFqsUVDu5ovy5bTQKW/3USN9VQ1VwcvYk0x+TlKXHtZZ2uyeVU5zqdzwd4wL8BjVBt6E/VlVly
rjFLxz5H58NxFv7IEClCY37NL/g94HlGeNeAamKULWh5h1iG5XXaNZ/yGHUReBfJj2LEcd2kyKAA
sHXkLm0xhwnyOJJ0YvNkxl8FFIVcrxUQ5UIAbCfA+ONEseVjsIMWaShMziqLFflohojSEZq38pg7
/X9mdvMG4mYLEW7jGrEJL/1w02NASQVov4hh5gTVdzbcNKB8ik7x1VZjp820M/M/hroYnoab1DlM
2bAmsdxn6cBaYN8+mfB/ek0+tDp4XnC9KmIkBJ+3uLn0FVlICanC1rvn/xjgEmZ84VZ57xWXTQhx
kHAEtald5LXPKBSkZqFXq/bhOITdHR6vF56BWYeyZ9ErY6AJ0dAVmPFdCxdZJMqjDb4AGNMEYGgP
zhzgxTW2fWmTnRA2UbHMSezEgztllGgNxdXkHXQYMWO3PM7XPPPcKko6ZX8KksTJV2JpOUKddUJz
DVbvfnna/eV0g7BgQCORaKldlNL8ZwE9vYF14/uzEz2ken8xQosNy6YchKiQhI6EkLK8M8gw92ab
71gyTHO0HEQLGdSjlDMIgxKnl+Al+A+xi/bVSEZkd1AwkdjN1zuv8jOYPirHbNnExzCBGn7tce58
wFompLtdNcvZFnxlFDl2kMyFzeQ8q1Iw7CEikEyg+KaLCTKoStLtcS6tVNT4FapeoVPk+O9RZw/T
K6PyY3dG2+Mtr1Z8uieFnIfbTLzQymS7lsqbnHIgun4tIB3kckX0qUMUsY6aFa0yI7B9geua8aL2
TCXFMffnN0lhxyZ3vLCcmpYpcNma7pT7JCBxdeAPHnXyLJEodNz7/TQY+a3uYHIMoUsIbu6feHB7
REZtbY5o+U8YGpOCMtlQBFvrhCumCDlyvERKAdpQc2pjIOyDc2Ds7qK5gqbwsasYXRT3+dLCZl5D
qj44XyhWRLrWsZjCzm2TSBA46izA7FVp4WHc3m43ayfaD7CqtT5m+vRLQobjLo/0eyHk61Qh9ofB
uohOoUFOkKEfqDQXdXQ/oK5iQjtC1/TxvLfrqem2E3SAFmpwTBMqEF8WdKL5S6GdDpRP8uW3ktUH
54sPLFjMukofmb18PdeN3Qj1s8WArLSacppH90y2N5yn4hlJdJSu//Z/kxfSMndO9sQxyLdDaj4L
TQJB9E2kKJZ2/MoIJHRwhwV/r9sDJHLoaEGXOLhBF6AfexoftiMUUkNyrdJl7sO/vllMDmWwHBJj
IfvI+Oc5cNsC0sZ/3CUUiowUkoqErPVk/ArUOi2NZjv+eZORMfWAApVHKVhGWpMChGUeWqPjoO+U
Ft5rCyD9tHtjOFkQwv1iu6zs5Yt1cvc856yfeFoy8lt+ztQ3oPC+/8n44dT2LTIwIG+2LBTMT+tX
VEx1uukw3vmPlKC7QlExqp4ZgwMAtKSQg0m/8HUQZvSYTnQ6fnnHp2xrONuTSBUw5q7spevcXAU2
DyeJ0pV0ZZws3yhl8gzS4bDQPk3JORhW/0T4uaqa9rYSQyYupJ7+Rz7kxOwHn97vtswtNeH7K1UM
MLxnOxlm9TIu39kf/7wU/1PCt9TN3no2wcRoM3rf5Z4MvyoJ3mwjJRmU9U4OjCFaO1EvsvOQsutz
VKNceARfSnFrZX3ioSWHEzn81DmIqB26Ft0Cs01MpFgxuqWZUG/o9VDR7fO3zRrpcm2rXL5n05S4
3nnf9WK0MzPTZ4KbBgvGiwLkK37qxigmjr/D9ezZ2PFIVXsiUZ0eQIMcR7w9GC127+IvX2vhnA3l
BY+rAbPsDwg0iJfvRNnld/4JcafwGwxFSa9PHJ21pQsQWx4ZhcbiPqCQ18gudns8OL7caQP6vJ1G
6ls4bZBP3UzeH3cK+MOeeQNEd6KlSUHwmAD/Xq0UOwM/xf3GgsgUFDt1cB/tGXp4hpmLxJjQ+saq
AVoM/WsWDSmU2s7CkmfPNxaGXoAW3RRo1+5q4ug08V/pNUga4IsBMujJiIVKAnP8mxPmN8s3H9W7
T8xBRDji5dIKe3JJB7tnzNh0i1+no16bvtPGkB/U7MSHcrpM1VgWGNsHnPI4lk0rj+IRHaFX0Nre
g9PbX6i2IiYkrcsa7ZMGKyZupm5MG7cc6R34N4HOADus2hfGFLa7doJOXPPW9UrL4V3Jpb8CaBUc
1Dfe8F4SWYmcZODd8o0acg+zJ3ev0jcWr8CfQlbz045BPVheoAH7Ro/DzLJsa0ROU/KDSYe/gIJr
RRb1LE0cRCA8Gqpv1yIVpzvgJjCIO4E9iOnoRG4b2J6kpgu4iOVKhTWFhfhYmEmZZdDkQV1dMkFb
cS1OCjYLuDJl185nm0a8SSdxc4TpvVK7sEdDTGJ1S7Q/zPmxb+QFrWtbgAPODBvawQb4xOa6E1S9
NUZgRtCiVD0K8jZjcSHgxbMfOyY7dB/SSe+llKeKpzLUVeyPM/BU4I8mWEWa6AF9aUHAeuZy5wnu
9gF+oDW03u2MebQbt8cg26fhruZF5OpAugqwIyThVKclFuGLeIM3l2zONBywGaKbh+q4tDt29lq7
TVBMjoH7wMkBkYqgNxNJw0tjSsOB1y0Go9yxej+j3akvJAXsYwnvAkg6KmvFB4SWr9nfp3ujNKJ/
VVVpwdtU8M9cCaasO4kWfAB9sH5i74RbmQ3Py1JPsBZx6ZMFg+VnG3uojLX0cCtYortGsO9hQxUi
BbVp/1Jp/1vDWRAKAprN4gQ6AJHftAxRkUXHIG2kxo2KaWD3f5UaZIeJkbSDIA1BlipTKvz3E3f2
tLtes2uxItg9/GOqEcZka4GMFUyfbNAFa5zpP1szMmP0SqXdXReY8ehF1Re5hYbn+/v5WzOVJzkt
QbziNmplYFf6T5TyMJnnHBzRN77sBA13Acaw7Flc22m5sSa5JUqHJRDfsurwwbMB8k+JHM3QhFXn
zM+/DZVi1scxcFHgRh32+citqIj+zWPT3/RRF0qM5DJDq/VTiWbCb4V5LI5UlA3M51kUsBirZ2wb
Wu2kxlRQBxcneRSqWSCuZ67BfJEJEMItW6UU09dxR1x0/b2vsFBFgg9oZIx5m6Jbs/T5LRzlKBHh
Zq/SpRoL0/9f8S6lOpRFsmig3dXJayn8B8/ISILtmhLVSHlN8FO4iMXf+XYcTRDtlqE8+f+kiseO
uGDzHvT8gU2dL/6frxNhStOf+ITm5yyp4JGVCuBEnxeNqmlDD/9uXQIxA1LyR+4iPhxoKx0wkX32
EmzGhbD+e7Y5GkVrvujPuf1HuD/BnM2dHUn5/bVWS5kzSPS45YnuPO9rrw864FuLCVHLGM3SIbOM
VzvjZwZszJQoMDXC3K0YrOKyDQEohX4w6od0RBlR3xcTLwf5cVvleamqq41KxqOhyeCU+15qmNIB
Iqs3bhJFQQrz9gQYhln5f6pcMJWHgxsZUrcukcOoy5d8boTYjbD0sJOZX6/6x5/dhUe99U8tgLzj
bXT5E2CVA5//9u9nXVkzcjZM9FHY7aDqor+fwdVQ/ctGZO95ogy98dtxGQe4yxxezUtooCFNmq+k
88q9+8/GiK95O7emB4/F9bWTBPokf5T45iVjeqkbPhPilqdYTW+Ro+5ubAqKp++lxd78yQR2y5HR
TJoNmYbd0cbtq4ysGmXKOM+09LucZ8Cwx0+aa1TZqLlWAN6E9+J49DFXolFoes+E6VN0gUm2svyt
BQIt5f/iDiEexRxr2uZ3hLZhwuNsNhi0H2O3yt7gypyFEZMJYtfLrQ8rMO62dWAiiW0Lerom2WPu
uqBMHbSgwj6ujH2ESIFDYdZtCnAdJDrnG/w0smdyv457COQiSrJCDTy3i5ZLS4D7MXQFLORce2Ro
+yFXMZXAd+P7R3am/iYd5XsgUi35WxO1ldvh51I9jpRGkK8y/yi1pgVAd0ZG2UbmRyhGb8PZ1Ad+
g9gc+q0r4lPtbMpzk57pTUsPpp98kBQp+4Iv/9iT3haAQRQKO7ivsU+kCS6zvhbNDPaKAwtcsFGv
fdB7lbq5rQ+kv92GLjULoqvstCQprL4OCnsgkHkpijqLRx4v9XBhpFo1UMJuog2ik+IRImRHTkt4
8RH8mIFBaB7gT/ET0jvKmMMJN5exnBETpYQzp1b16xEI3I+aDRo+9QFBj2Tzu6qqfCcpJj1fazF2
Wzt3r4GyHYtEaOBHct49WtyWjBWzu6dt3D+Cbx8bkEryQAJbbaQVftG/8WdblPLnOLt212Nxp/fV
LZl8HOjyeA24I6/GEP7hE7ShuevDWfPMkhTWHO55KzYbRdjHDmnluhegwp0zHJSWAjYyXFjWV8oi
0Mr+jGjaYCFgtSVbcmtrLmjCXacIT4kbl8Z0r81j6rwy7KtK+Rqj6sdwiCAQpkdUQ7XPVBi9dsnv
n0hB6VfSY690bHwdFi3ZvezuunaAFHol6wqj2y5mIdF74yZbaGsVy8V3ineLdYUToJrfSamuJ4vJ
vvAR7ZbaQiFAtDpeFvhpW96/FNeIhEcttekNq9NULqMDOLRPMxl34BkdDCwA72SzuKv4LsU4jRMi
G0CrfRwJtr9m8sTS31e2PplQL8gwDsGrwMyimmng25vbbzCAgS36Jv9VfXgygKGZjAIqFy9Bqp0V
ufdDHENmhf+SE+YSVk/f+js39UWIsHsAdgQ1AB2vz2ld+AVYJFnKpvodO1L+ORIfg/OcVGNpTeJq
BIRuPox2euKoKT8U/K4kzGkA09iP6nf702K66DRuJ1O4tR8u+OyxSmUP/y/cKON1Lf5GJKKZM9oY
xSwuqFZZkBsRJG5Ojk42X10JmMkp/JVCsTaYjRBZCKfqoW/rV4Ujxx+0GRxoYA/GgteV3VkcuUvL
PBtQEoDvfWDHZONbOJAGaTnEM6v5yuHIlI7HkOt955gxSDvHaQj/hls+6ayO5hQcrSjcVmFwFl50
40v+DcRJXT33i2lDr13HWKhJGb+2Q02ghpYLQHT2iNNzKeWVdS89zZZd2AsQz8c5dOE6e8ZPaBo9
RN7rQp0PoCS5sDtBKFt56v7ySh2GhosYW6W1cHkx5qAGmm8c/VmgfF6eAwWq+EJ3etjzPwweK3nP
F8ehazRkZTP3Ut34WL/cK/eKkba4X9TTivyFpjZdT4y2Zejz/7xViaRQRWfmzfnuTmLIJsVz+6eE
hLwDyh7Dkaa2HjU6o1XGzzyK5Ibiul0Q2t7TXwfpSTSeOg7p1G8kP0hS4JY264yzY6A0n/SqY3sD
DxLhR/8AEBHDRdwhcX9aPqzUDfhNQSRflP1mtvS2NG/OkN3trWdIS4Zh04kXvH309AjQ4FJ0ox/k
l9ubYHbQL92L5uMljfuLt67y36gsAJ+onfI0BeXSLKklLeCq8LQ7dEUazzcPJ3jfBUz01ekybHeh
LFdfCBCHzGYPSYLnAHxHPZo766rPAVIEwrAkbWMCjcdB66ZAfcSar1S1zG9UFbCY0u5fECsxJ0+2
nQ0A4uZcNTqiR6aK8cMnbO1S9fSIhRClJMkV/glePScNJ8VOxwQcsW4spyxOEo1bpjC8tFZLjIGD
R70t1Asp6SR6JqH8nJmYq3Y0dOyAiwdXSb6Pg5txWln/VuzawgPR+WbqMb5mx3a8FhSA3I8fPRl7
nuRG6/qMiy6XwT89T4pjRGDU2k9VRKpPyapVLbxwC3nSlrLXuTUsStg3zZalKJ0qwO0CpLGqNac1
0jAcSPhphybtWrDEBAyQ+LRQdlnKhzxNT6l9Y4XsKXjjCWQtBYTJ+l2LPj1vSZQA+l1adJ9AaaNF
qiAl5E/vqETkXENHk+ew40Y8pZmICYcX/10znFmndyGqII2ZvKvLUrpJxo/ieMBf8XCqTp3VuBzJ
z+BvtYXPxT1fVrC3TslhX8Eq3t17mjcxMZwzcN8uYikdtprzwdh5nJ7kGnZx2p2cUiV7EXh8QXfa
lcctBv8JAcADSeeWimLSC8LYILucEGPn3/BRKwFBt8d0dwEbwBtF2zUQgtjCDu4Ge9TABjZxgd2b
AqLGJT+suBwFH01ESUdjGCyWoBDpld8KjKw+K7oFl+R4nTOs3EtuczzdX92gLCaOsg5y+7jbpxTm
dud4HFKLzTfsa6621mmu7KLSk8TA/nVSRW1uey1Fa40demAJ2hs/3zS5De2MfOqFtb/TnDr5YJN4
7grTUiJ4V67Df1as3ffpXd7V9UHfbAxLJXv4KHXcQt5t20p2B/OBmyU2RpCnJfh8FH6a8UUheiCm
wzJHK0EvQsVUZy+0UWu2o9OwG1tvBLOetU98m9kFeuidDjqiuq70XNCScxrwWndverbcAH7WrBXL
Lj2hqR0L4M3JxLa7Zi51c0m6Gq/u7xLhwbfZzJSzLynf4bV7zDaaWIGPTG4jqsg91btQOsxfV7bn
PgSspc8wYUYeQKNVomli562R9mZsaB6RPFeTmPmEH4qre3mfoYEqyij7jiQnVgAGxKmLbc8QHo76
X0ayeEUVTrJIuWqyWmMdT09jkGY4+HWS4BRJTJhyvhJywKWlZbj8piTp2eBOR2+4AitvYtxjHLgp
gspobQPK+xOcyzNDY7XpwN67+5DF8S3ag+dRJ8gmegB4gMfVzGuoRSF033GzkeQ7UiHcQqauaQHm
l/nGfYmoavdkIWX63QFPs2mlH122sM9wddw6PEEf803vRZwr2ZIjMWO/ZxO0mZBMDX4MCG4FMOgW
H46Ul2qCObopWGcQhjv5CYz/znvH4D5xPsgzxuYP1DtwktRKlmIorZa4N6mhvsf/1TdPs+tOtUsQ
eOYbiYWDi3Hi/LyZFaCQ61kb4FD4c7NhMx3a7ZJnqvKYSRkS9pFk1hqX4nSZkDvA/l4/9uvVjtdi
Md6+eYElLfGUh9IxxlwDO3ISAZFSKBb4s9/Sd8YTthb9uoy6heoMdWxdpXXCv3sMtcXGsOvcCJtA
/5r/hYfVd2vMAtOHi51rdNoOALzHGe8rqu/ihgFUCuOjwpZiBXoVHh+fenpND7l04zsW6CJoo2sN
rJU7cZCHtTuNa6BG6Q2g2IOsgrwRZxGCvkBEo84q8c0c3XB7yIme5KaGxZHgWIpvlxmLEwYcgrMs
Raf7rXjzwiegTwd+UDyC0XfINCjBLCrEzPEzwbyWxNqWPBUh0hJjuy2oIg/ox4TpXHFR8ZiOGcBX
YLhoJ0R5qPOzBZYdx3VEPa9VAqZ8n8q/HywBfDwywIlRtddgL+TC1Mq4ULNLUy9XrrFDfAWjw+Av
5j3Y57YA84Nok3rX8oLTCuEz6ig8kQG9rIq7z6N6QCJolf8o/GoNxIM5hz7J2bsNog/x0Rna9d7M
FKfjxIEhgGu7NcA/cJQK8QXgewsPJXZ8YqEihEuSGnJhTwLYHEtxQvnRCy7zxffq8dgBDzCZLgpE
RMg989KDQVDKSVoTNp3PuIEDSNKke6OiF7DSmgf7uZStB5/+TcNlFdmsbAUQK+++CHg0m9IK97US
wRl26vNBhytqXpilyckUhlJtG4h283E1UaIzzZwtGJMR9el3HFJ7aMqnBw+/2tbVHegU97l5+PF7
YNfznon9RnnGijLw6cx4UtNjaoqckfRUVmlcUnWwUGYSZh8YCHN+U/D0Za0IMRcNypGVXfpP+EKm
Cdov+vLyqDyZAbgYQFw+Th4gKEKbdfPc/945Zl1+YuKrps6Za0puoBzJqKM8+EU0kBj/qJyGJrmA
EZcw6uLKBdyd3+E5iDyTnv5V5nryXAaKnB/u/hE8QIKkAm96m+V30rpMoTkRCn+lxiXnz6n8Mgc+
Ca+eqQcwwPPC0zAmGE3QeatInmr9lBE8Mk6S5LxVv6gRUGkXyjt93QC2tc+0yx0iUgKXyyh/vper
LjIEPBj6F17TqV6gLp6TBV9lJz/nb7GDn3rJ0v+gnl9gg0IMPxchfqLCUNxhRiDn4/p/kfxJVCdU
ZtVjSQtshPlu8HiUEzcELtiKEYNFNwQg/yjJ56SvEMRmvF0zFrfOHnyzwsMbS9T1wjKy8nIRwXdX
LHJJbx+EIKRkCId5dsLn5d9eNmK1ZKVeg4IFgzxwclb7q7XHk8jUjBnXGgrlR9CteKaWXuR30fXK
YAaOCecAWEQMZToYXw/2/DtJFHW5LwYUDFttlHsWiPxNpjD70F2zMTRj18wWjq9VXI2hu3bmgy8w
BqZpSR33se3+z/P5zWA9t/BgcKZv3tbLEbvhXRmVzUr7EHoKNyVakeu3ON87AsvW7irvq7vIdslD
s4YGsKONtbtiNfZVbnipAHFns18y1uGYT7yzILMvYrf66Xd2SNNlNgEIiZkRe/XnuDgzuUAi1o/q
9omI0Tq3YtgLtuW0qtR0z5JJCcBhC+jQU+esKqpa7oy7mFNZxm4PNzRI1ausa0BjEBCt2mgqj+Jk
XXPWydmHRk4fhzv7Wu/1Oc94lBiR/KKJc61FktlM9m37usEc1dMD1YwOjs1keSbATLoXXPMODZtQ
+eslGpuDYpVzqydF1sT+nVE+QClsNS0ZBfnq6jtavzPF/pAHnZrK9GKolY7HnVo/aDYj5ShKp8yv
JXdJrRGKSODA2qpbX8YucsIDBEqwK0Xs8HKOyyF9NZ9ESdHkiVkDHGzfc5qirPyFAZJ8mvUmuKHC
vic0AVMsVGVdmbTeWuqEQU4n+XjSgaG/Sz10/SqCxvzeOXZgGS+H3gfoKTdZKVn1p3M+8vw0AiuD
+dUqBrW9ubk4bvZ42kHxFojhnmcN28ahV3Gm2XKYW1k/vrArHt/Y/yfQHfrAVniG9VFET935yoP2
OsTyRyadBOUFMeKhS8AiZgqAnAFDC3x48N0k/5OfZPW6OPRXefTYbBmWpgrytotjJcaSA06DOpkH
JZbnuGh4XMCMouSlCsBGNHB/UnF8IKvmLdrbp65V5d0tulk8CwTFYZd9brFVBzScAZ7ve80g8we6
ofZsRubEr2wy76MDRb/Pph7VAMfHeGACgYm14u6+wqaGoX/ZGRm/BLLCUpFAifCzJ6/Y+Jgk2amb
xkVmlG16kQ0wdHe69GZ5u8C+sPIx7iE8hM9xCNxSpFcBYMAxbRgDiYEOUXacZzPtkkdOH/kAGCV3
Jf70K4yI/TctPHe8HE8R6IUBIF0iFD2+QwjZrAD9J9Z9iVFBXRpjLtVD4o8hPYHQ1kkJLNRgfFxh
TRLABjsz8CRVNuCHOTZpfAtF9FU+tdK0tyWuKrC3t7if8oqnXLQQVaG+ldI894JL7adnANmjPbT+
YH/5eyh7Cb/1H2yiWJLO9g3LLU0u22kKNQE0d1eHNxPkFqvWe3UJwoWo6GfA7gyHLA6dBj08oa28
/OuTvLU27/egUabCtuUrmpRv6IDaFVRtPUpozG7VHgcegrzc9FP9FzXB7dO6gBiQJ8bE/vT4M0PK
PSqE05XbcAXM9t8i1e+Alrn7oZDzy21L1iTWL2i7esWTjZJeSQ1SU2UarXGgIYe7y/dwkgHlZd9u
sinCLVb0GoeitVKX+Zc0uNu2FCc4g66FAqSFl3PQzFkDqLRasTs8XXclQFcC9c6eDxC0pi4Gpjty
MGHTbzSCsp0Xrw6bjSWmT6biiRSwMn0N9O+kN+Vds2ZZeqNHPs3UsyYR9jsjolvxxZWrMqe9hLV8
nGhZk+KsaJP7rD9bxeSNiNXZN8aHER3+S9UiPRULERGbvk65pnpFHAFkqN9+hu9nU//tPJE3AVio
OJ1LHglhD9C7OXNa6DKkpYzPkKIfkVwe/2YKAsMrZSAPYZ43MQZGbwqFBzOWj2+/R6VQVR4avmoN
PoW/sX3rkPJUemily2jZjLXFH7NzicA58v9BY5zOcykxT5wkxUEncNuDBxZdIEgZwTfeXjcKXCav
TOdA5VM/upM/IwNQUKgr/hg5mdH1ZORHMfEx3ewQ4KRhL48Fpk77zQ0VufnlWIXjnHZ6PmY7nR7F
dJtpFmkWTNdxH6TqZDWIkFErR3rrHtJOEDyayoSgX+W4H7Ipq2lOLrgVjAJsTgWTY+1pmO+vvl3B
Klo+K2cxkOVXySkFEggrnnriFJORCNbrS8V27Al7X844rnSAcGBQw0DXFR+uD9CkiIoaexiR7Da+
CPZI47K7SIDAMzRhg+UpkjWF62gJcCCZ9OGPsTHChE8thon+8rejHotTEEvGfP4YArXGFe/zr7yH
ujKG9rSANvItzvckfp+8d5YAbdJpBD3xFU/Z2lJUyJxDlEA4j1gb9ak0p/ONsBs10rzThfpoEZCb
vlutrBeTeqlmoXA5cW3DRMvtkVpz/k4TOniIKGbyGnf+dlA6NRwUVJHrLHHLbuhfhDhJBU3zY8ER
79+XUyz+xXEUOb36QqXV6gIxe9Mes9TscX36k+nPBLKPTaExL+gutHCfcpT19Egl+x3CmkO+CkfL
03K58JS0fVrP9dP3EOT1O0VistQ63OCgTSdaUJt1mVdpAYqmXwXZhF9OL0iLwKlZvZyYIJ/cCSND
mkghaYpQAX0XfpzePIq0EzSzt/zsHtoJ9X7cN5bR2Rjh0WJvusv8lv6HfxQi8SW1FWJeefmD9js7
7dhtTem8lGNcy0K9rLZ1D3Tl/Y+2EM90VIJ2jWDmFng3nPZdy4JR436St+hGWHbTemMMff1spMQZ
TtUbbnHhXKlqkkxW96YBvLZPMaXkgrEelgRtPX/Vew1x+CsSFUPS4lF6AnQsAyiKjVcS7MqGMXsh
AKETX+hWPNLQjt5zJ3OCwrHvf2GtF0rgsp6pQvbNrdlQ+ZapMW9jz41brwzQTKER/wiCcGHI8cSX
GrrRFX7EgOniL7VcsJG/KC9nqA0C4LLltXigYBZzP10gGj80K7qiQpM/2Qt/72RTADdXIKjyme1C
nV3rvu/nrGRi1fZJsCntFGSpCrzu2ERsfOYdQDZn1t4pQbf0WfOcvRqrAaaxElj5tC9IfS7GGGr3
ffARCC3WiSccc5ZR0U86ajJjcqOjP53DwuP3iZL+EuvsL1kgfRrFy0o75BGGMEkPWODoGUsUqaiL
Yei0ILBGXGQUEPj1w2gijeH30aeVQGPn9kcHycNkik5e0l0kfwfkZG2vGCx8cvO4hhOVj5oGjHP5
5Xt7skdAUsKQU4DmPbC/tnx3ditV6eddvt45UjZtdDnACTPuPOgjYVwb0AZHAOYEP+7LcjI0Y6nj
kc2ruhVKDA1Kz3NF8JuoCMEU0z1rdDBlaUUuit5+zFkJZlNItBqYAWaVegK9xIlJNk87yzyDqD+I
9rrYXRkzXQdNdUFgECtngH9nBEG2VZXATK5CXGNNpC6Qku8y9JgAgJDMWu1miXW5O7nYWLp5ku5V
bTHe2fVxKDe1L22Ko9RfkkEeXloXJydEkQ/o6Yk5CkjWamAQ8iFwklEba210GTmSOsIJtTva3EnS
9Ldgh9RE6I8rhh198s8S5B6XN5nvpn34VAD44qetpXWN0M9P8c0dWbIDMo382ZKwhIlOFpFsxRBb
SBp4ZVpvApw1eTSvmMky+9LR/CyxRRNxIqjRoR73uROlUyWzy2/UGhKo3A3kwzj78HezYit/oJoJ
6mZEVgrdOB6WnnocSVQfQ18AdSlMPiGYZZKI47AUpnHuXlLm2xs7HaMKqDsffM+wqP9HBc4EJUbr
DF8DrXmfHfY/KUYlt7MSdDZLmxnVTR9Phueop9QysesgeMK85ROdp+Nk0ZFH9xrt5oo8Ya9a5RIc
I3xLdnpIv8xBhjsstkIf6zqAMK0x+c05LeN3dwvGZGXRyqlgyR+7OimyPVzOOGnm+PsfTAbNZaBZ
/a5brnAa/RzL9DvBlTHFp63g/58awBt9gXWI/LyiinxM4gqF9yl65YwAhSqIRp3uqq5s+gfSbgYf
6ipcJJ+dLAtgkwl+7MmBFdC1SY7Pn1N1Nq1/4LSC+bNllmgt5JsS+Tq5nKeQnSaNm0+vkJGPZpTP
I1hETiAqBjKKu2k5soCAn8JH0Dzbf37rbp5H5++SD7QLtq6DXS//MLAqN17Gap/qRZC7xTsPA+NV
JIOkk1YRCFL8tkTIrHK2vJQZp2yC8+gRUyqE+IhwF9Bcz+QyYtefVBb3qvm33ozjAb6VKnleBeiS
gGaGo3aYvz1EamIj7huO13bhY/39wV02PnF9hjjG1xVRtnXaP4jSwzZSEBdJ1M8WrDh/nOyXSfOI
y02puNYt5SW6rml+f6Sp6++QASZU/W/fIrJoKeqFySP7eHzfUHrrDLgkmJWLhLrTxqOmKtAcV/xj
BIstYBq1Fj+1FKZdTi5UIs5UWLt0D6BB6vBBl1PrQP6oOsdGiz4c2sXRnBmyRnUrWG0kc7l651KH
owjm0uLhdRnnofJSqspAgdWzvqgi4afZLQiS0ym1hv2Q/7ZipfYUiavvxCtPz0Pgjsb1VMj0imhE
aNbyEVUMiRuwtOcmFvI03f5UuNOj2ArXW+ttPqXQhoxMEuLC3y89FUUTgeZpLw/SKPoR1H3t0tKp
9Ihpz1K3zYpVOvilD+ulhGp4H7LSefHh1WMwd9hSYRv+Nd07/+RFfk70EWr2VvtZKPwuBeRfQRdo
mZl/x97cNQyBLNAqJhq8Wt+VA6zuobJ75Mf9+9ayTjvlkNp6X+zO9WjGoVNPvM7ptdgGBW4S3QRq
xOCUvFK4NBYOCwpECwGHAl8dTbxu93IVI5IXUTxapngvUZumrTBfRw5A0ZqS7W1kH5Q6oAUcTIrn
GJdUKQfqWOntnLvt33Agczp/vUTeMk9sgB4HY81ujT4ifVkL4Tho/RwG9uvLSGL4Rs0Wh6FIPqcW
b7p2Rr71ASvfY4aNB7ZdHzCReXbE2XsWuukPLSya0346ASAp2N9t7iowyHGdTpoQhlpeWuiYtlro
M2OTfl/p3Lx8zcMX648OwtjaseF5s4LDM/uBNQhMFSj+BFHnf7vKM610ONBVqQx9bUsteILGqxrQ
YleooyX9oxr/R0WkaVbu+oDC3+TLpqhgEkGbKuGQUSDieSBDPFVD9yaZdShlPZKEc7xK978BPQDZ
GQkUBq/LfuEqtm3ggoYrmfCFgRn4/m9z6WiSWWH4UOP/2Mp/XbE8PThYKHUxAjkoDkXMZRD9tJf/
qLG/m8MW4jNcObxLR4/LNPZsWiwWUgpby9Hxi78P9wRI2O+mQoWUEnaNPFYr8iBA2IMoIw5uT4wB
0rm0wDYFC5Cjn7gliRMzRfhJY+ne3ATFWR+N/mo+cvLTl0xUxmDipD6tW6+aRraAalz1RqzkyC6d
IX7s25noAs88z6zVWfbBuQFTKg9+8IwUXMp4rKgjZmRhYvvMGemgum8VWL89OFxso6RgMgNl7RSv
3SCFdVv0+3UNhvzG9QToy1aJNKTIOZP/qJboHC+comey8Wx0HETW67YlsNgZJo2U2ozvw8HnK5Fk
+A4OvZLu01oNtM98GJ0M3TSyc32TeMeDrOS+Q+IYzWb9XKfyBBcJx6D6NJEdnPgTnN5ySlAOhfQS
WsJP37cctfk4kfGVwZ7GVlZn9WO1+e8yynqj7sjzTMqi8rjkqKKAorWKW9sxiJveVd0MCOGoeLQD
0dsMBXmqihhhNVLf9Wsn8QX612qn2tBWPJiq6EIGLnqZdbKae7NEOPIpNrf9vpChAvCJVlWu+et4
xrgajhyB8HI7Kuep3lssCib03rR0hsfTnTf4ieUZsArj2+x+Meer6URLZr5wIYmvLb+gGk2huNdm
XC/g50ssHRFjSGma5gL04gP048zaLxLDfiqeMcd0hb5L7opNhZCRR2obOH/pilh006pVanhP65i7
vqMch3q3ed0OSfqJ38e8l0hIAWMkB38yuZ18fJEjxZ//1IzB26oyNYtqE0+55kpQaHb67eFNblt+
50YTk6VCd8a8OO3daykGN/hE1IzvVRGkmljFHf1pJPa0Kns6aMsJRkSNEgch7nJhzZ0ZWE3Gql9N
kBXcULFO7QoFC3dHUHukuG4KHQV7DF2PHaijZk94RONHLTEhaoGl8COL8biXN37WpZEfOriWXdSA
xhhZ5642EEdtyDnn9nZxoGw4KIIrYNiGiK8nbGQ6QLmOuVnhtG9zNNj17BxId86XrlIvgCub4/Sm
W68TYFNZmta4OPBNDgMm6VpPnGBN17IV4pWvZX/b/WkDvPuPAiYXHWGkkK1o6vL84G0OcmW9YEwQ
E15F+DehQF1J5mM7ye4PsxT3xwWetx8X6yzrWiuWihyzUmRNo3bB5odta82BDV03ijVGcdjVeEzc
oi3bEwO/ignUOMcakisSepPNZ7stz2LRzBFWSxjRCtj48JZF55HqU0wbVs0jtBOcQUutfBo3EQiu
p6mq6dciNZCDFF56+lUpa+agxsVKSPC/uJzhlLeoWdjYNRLYSg2Pbw2LXca+EfFgMQNMfO64PA87
g9kH7zE5QndMW0W43RuqHBYljbP9IrnAX/v97vw/9jHoKiKsdmZJ1Va2apg3noDLAjxNMHI19YTN
72TSJQu3n2T6YzF+8QuqtzOOQBO/gVRBdi00QtHHzihzAp5HCGUtkHLptIubZzDXRbDbj1qZ91/U
5G+Jol7c+zm7p5ipQ9GzvhPrUBnQFbtuV1fJzEt+YO8NRHN3uzh9xi/eCeHclnLHk9TwonrjptKq
cPNY2o4EX7aT5gd6k07llGDyO5foF5mwzm53Q5eEEpk320pEzHLlnC+DEv2DYXC/0VcoQFlQFEzN
Hmb2tXQk7/BkTBEQIB4ftu5qrkNM3nGDhyfByokfOuUhx/f8RS+zUlSoUyw6nzPTt5fKiJ/Y9Nhh
CY8SsDg29CphutOV0cRMQF0KSCeJ8+QLNRNg5lOboof8RvENLYzz3g7KBiwXxDyyEETi3Cw1NknE
naVTxlSakJ+Q867youKC0PGuBfVe5O4/sNAL+GP9ivS15omv5iBGzM8L3ZkEMJRMEEWeUDTEqaWj
2QSsSqhUsbYMLLurF5X28cT/Mybq3dGFDFaUs2m/EKkUqNkEyYgth/lzWo43OrVb72zafnZrfETw
O5GVnXH0SEBqZgjnEfYSw/j3IxyKnODCMR6jdHvJwiiaLj4jGVCxi2WP3htMNXFWe5yL9RCmTx/x
OU5fYyv8MNsELCv8N/fJp0Zjy3NGMoYNx+if9npBTwaXD0zmo5IGG8nYnMYmLgCEHOzaYuD5oyIE
K8VRaU/Jvh96F4ZS/vvIoDgsPCCvUyGDp2tjY6aUltpZYTreH/JO4x1C31WW78LYmjxp/ChXUqA8
xyjasUkarKwe5ElEhDDRUetrbzxvAqPMPK430InIx+VpZbS6xbiSahMOOMarXr/l6lUlVhBQ9tau
D9d7hmBg3J0MzJUKZi7v3WLkcBArQDFHtShOmvnl5MwQjPNR8OeOZcuuZJkZpy80MT9VyGplLIMI
nF2oO130BF44CPlN7QmdZCsCf37YM4jc1Ky7w3ysVoCNDim8fpgKkZ29X8Vh4cHoYQExhvn8pHJt
WZJeLlN7BggVRS6Hl5xwCiZpddGJUmwMkanGc512qdRNjB/A89ol0U2HQ1ybx824I6y1mTRDNDRw
ToTtD3ZyS8n/DvgZIGQGV+GydF3H8O1oEyN/RixXqyC3yiD7G30QD4sJtE+E+/qNirs5H1xW/s8M
KYbklD1Nb3x+1jKEm+xYaTX9Y25vZb15Hg5iZOu9zrf++kJYzuD6HE2p8fOqtlhtr8f713LOuIcy
A27sFIBzYDJ4ASBzBBl4Ugo6rKaZ+EnQQls0gSzTu1Etdcsq09IXwvcBPrWWU34tKVY1DC27/ykv
T4IWa0UtGLuVG+qsfGX7PJ3hm2gjLGVl6wlKPPT53nDPNMClSaUePGSnJuxM/cs9s5NLwF3ijYra
J8iD8SDCakICU1rqS2DVidzNZRZYShA9FScyCYfqoNgw57nLyEXB2zETYi7/6H1ILRGf+KGYEgHJ
/nkAB9pNIeNu4e1ZbM7/eMnMTXaaRJ0M+IN1tRyFSnTaqUeDgnTTqDVnFpIoZLcGl7JZ3tWn+eme
IEVW+t3xrE42honxoark4eH34lQtMl0GBnn8d2eIyuHg6gv6H6ytqd8oJvE8cZt/+cEMhht6W6FO
EpESS7mszVHwVXzPzrS8yMGpEJdREQrKY9o5ZncJwFfdFXz/LB31W7rpFGewMKCARuXf/Xy2rp5u
eC/S2LoYpmblVJpeB5iW/pzfH810ZrxNpQKZbAAaNyriLKe2A9X7Vxtq5GU08YRz4g7SfAb2/oZG
H23jBa87xHsyV2ogURRvL6j8q8GR342tL8f1Tzad0kIfI/mxpLn74xh79vnW3UEM9prjHs6QnIdr
d4d7+r2kPSzsA/zsyqNLqBqDHbVICLIWe29JT1wfwN3ZNFhDMFTwRyWTWD8ECeFU83EHZ6I7XDMg
C6/MGVA+2T9z8KfyvqEvGAU6xJx9Y+ltZikUzsFMSSVg9X7PPq95jPneFL1PZh9eKDQdCXowIOH9
tguib3Gdrpj9dOej48RDCdhygAO8NJUIF/tF/55Yl5Xv+iyXlSEHO1ObWm37EchpLErsXnbZ0PGb
lwPhTshplHukLpfWRyEHk/XZHLM9JtWa7CH0k1Phs1RhNKmebksVGlN/cgEDlRwHR7UXLcNicCRE
qXiUmzLDS82ipbOaQz31W7aSkVfUnPNZZlIXElqpA8ENbk0jFMmfDf8bLV3YFstjvbgCO1IyCl1g
mGT2rpO2nhRcLaMp+e8QhLymG6iPHo04wxnfo2KoTSvEm8OhdgRlbP6yZRrg/rwi4Ci0SXoy5oRs
oqCBLGs3CsbS6Wrb3ZLN85A01NNwSidtvq/7YUmtFaANmnwuffkjzJH6okU/S/guvVaQopXQwAlA
SrluiEaEiCCEry8DdVgpUFf8udk3UGq0Nv4JatEmVPHGcKWXekbCothU/Avz6++lPnJuGW9jxMzX
Nsa1Y/zmjN6UWCKkC/kAnkmeVkRz5B4P64cMXLBOR4G5RIeKp0S7xNLCqdHPQ+bG6cXpssou3l12
IQc8pbiuR39RGi1J8kVJIDuEnY6TiebTSIdqZLb+2d60Boiz+FlrgU1j+gQcZzSVXTR6mFeU59vl
gFXVFbK9UYwxA5xvaYoP61ROs47jnXXtYnzt2qYkRu2joM2m57tfVRvwSKTg2CID8R9/Ndv7gSVy
fJBY7X+BAjPcc5cXCj48+kQ+tAe1iFS+sFB09Uc9HSn3EO/lGr6FslrI263suS3bvGsG66Y1Spa/
/eMWZi/UP+Na5jM/cal7yDP9sWjvUPdnrDggxF7NeieiC+Jk2wG+hfjd3sTnseKXHuQJVb4OPb1Y
Hmr9p46LQmxgPOvusLI2e5ezzyMCQTTbZJwCHDk2N5/Jgm8YEi3uoNs8lnVyojhm94/4U0lhJR4s
r2hCaa5kOWktACcoBNVdlmf85oGzqVsaDPMVFIQ88fBcfW6pjie2MagPUElLPqNh5gYEzucQR0+e
6G/NEm/lbc/gI1a7gS8PKxybr6uah+1WIgG6aZkpGsD1uAYisCVJhAFgcA7fhTIb96cU1icRhB2X
GDHql7yl3QTKq8xplHe78vTd51aSrtujDqnNg15rT4sva0G+EbXoFLLdkV9+zU71KHEv1dkp1tyD
h0cYvNWzcXmG45pVyawnIaAIIVweL5knAiiVhWeR29t8i7EmPtaIXcADE9u5DSZU4sUTWI4Y/sok
HsauQ6m640RmyC7191gA6BgQ6NqeybBvjCvfB2TmcqB9LSvrF5lxZVkr+ErzbPHIdhAnUAKLOh3s
kIzx8x+eLQdbE9ZSXczsHRORiguP3SG01viGWnocBAcSpeGu9ZG5kePn0v/xMS9teKFtGo2V+JRk
AFm94UlrXqFhK9jY7HJjK4yEBQvrz6KSLZThwKBGp08U4p4y1i2FT9zJTLrlAufTwEZ92pK/BbEr
M1Mmr3Fy1M9GLz5VhYCtSOMFpI2Wc5EXt19OkSu1EiNG1QdO5RY0bYPkh/Wgi9Xvl4oBOYCRpBmW
BvdrXC3jkCiNqCZXfQiMAMPdJonkZy71Mcp+fm51NQWz09mbzTNZWb/8RCmkFmJOs60ZeDXmkFVl
LLb/lGko2JBOBNyuG+FXtq2ug37Z2ZUSVTyeaGG8NbgxfiSGmbrYnUCqe/G+MyeNpevdf0Z0Mdm9
lCVvx9fJEBXIfm8oy2Jv7j+4xc3kurm9gBALYzwvKpAL6CwkR7LisvBLRCH/Pjc/LVwBIG1V/vDN
WDMidbfmf66liKPga14/1mydRR+4GQ26V5lQEa/AL5qNRPalt+DpaMUyYCgEtBlx1g/ADbHcuDXt
kbqAA4zUpCS50pwBnZR4ZRmEAM/2HfNxpiuFMNdF28fbbmqu/aJsdSaAIvP0/HjIft/C39HTD3Y8
83HG3wFAotlrjlCoggVMTyotSFiFLAorDMn2zAXks5e7TZUfR7urCJHsw56nL2KBD396EK9Nog0k
M1c+u4+6Emz+DzFKQJYcDqKYkQUjAybfURt+k913765cJ+ftIGDL6y5wUjfZv+enHcebYJTTpNgk
sgI660n5lWbSOiLtVx98EUehZ2G3z+3oxzlLF4Bgly58+i//D9cLrs30tpuzjzHqot5zgJXnqcqy
FXTIex4OXlaijRxi5SHnyluoa0MPVqckp/tWucB9OtY4XgYT23SPKFORVRKw0T19+eb4BUFmcISk
jaX7JSPIof8yIEA92m9yiMKN/L8iCr35zaATrkShqIkUeeKU8O8LZtaZl3qgY1m5VztlqgwmKCpC
5U+S+/01wNCEBAZj60IMBYGOQ/EPI2sffDexIlTCI+btnGwILfps7pK6s6Td7e33zlRojbKyg6Qh
QUmwgd0+nOXB0U0IOiyA06ywo/GYZZVj0MnFLh7+qp0ZTF0Ep4fllKGHlvbElDWwHnmeluNRKPTa
lyImrQdLCInGiiO+lzAYiKWKw0nZMShyDRBT1ou3VnKP1uWvvdlmzh10UnA9nNpkK0FHs4Kgxi0j
JFKgqaIJvTamBwFGDNzssnq/mtIinEbEciaEqs+nWwKG9VqMClBfJj0cQeTDPSna3txi8ithWcp1
RqH3dDmj/ZNyLeBcRlLL7FI0UMHaUOyCKfJeAuxSaj4whVq7H/trPl5BFArchsn1PTMfe0kj53qT
a4/w2JY/Q69yoi/ay3ZOkraUdjOWJO1AT6sKEn5zaLc09OqG5IppK6+WUFhBi/UYf+6xhIrw6XSi
/WXkhR2p14ArcrPUoK2KaKDYWEUi1dGl39SZin0yeWQjDRXytad5hNZ0lUqFNw4cf46PA57/pjVu
knLP8dj077tcYMooBweErZ6+UtblA4HX2rxYo4Z3VrMel9Cbw4mEk+Hg9QyaT10XDtt4ReZakNfY
10vuJ/7JhLxFPjNdmzQhe4pjf8sZ8Q5tADrpa6/2ZNG3OSiE2lMQGARGPceiz6XGAVYSxUwFb2L/
4qXKwwkpkuttFO3fnaJszCPBCKM15QMbQ6Adw6AHqAFjVroRFQC2D+O3OLTAVuYZXg4UXWJhia89
lWaQQCXwEIiY5z+CKWyE/XcsVLaPuyOFL+WYhKmh8GYM7CnTjcIstlRmPuWCr/toWdc4tnDAXPIe
26tO5y5kax5fz1r09eAKl612Ny1MEz78pHfSrMx2g/ajIAAK7vfE2jyAqh/FPOB2JVhfpkkj8FsT
a6p3ge+1PM/ZZPcEhmoL6OHuSYcnFLyig5qo3xHrDVKKY5gbRWO7AnSRY+r2tdqcHGZ1dzj5O7g5
AlsokxUifu1lQ8D0M3k5OK4AJ3SN0Y9u2dF9bPoB5cuIdAmGjN6WDmNyjX8AwT4/EonFKqA/cQx7
VpRif+D3wANPdon+mfO4sV2K9XvW6edXWeOFlSRzrVxCTTm56ZOqgOAATo0PFJBEcOgG6pvK34jq
0Vj7FrPCcK23k2Q7DSYK9h9OshR5P8ZBuyUp4p7/m6dUopv0azV73zxB5fIqVi4r/rA2qRK4dFgR
6fv0q9LMa3geix9xA3mg3P6amgeeZoSlCqFYL3fbLFIOg78BtxVuV+IlyC+cF4/99GHTx1JCzaLP
lYFHCyT+lQU8rYOXlQj0/FH0gPchQWftj8FYDXfAqiSEwCmg1u3oXsADzECtiZc9QKeqAA/GwYpz
nA4tRrRGe0X9hNi0cWtDpF/Gg8H5NcbTgG2aAC67VyQyqHiHKzm49xZiq5YbHGsxQYJ7YgnEUwrF
GQnjWoFxzo8AHDTCnjMDaTie2leMPLegdGQZ5SIpVSFfH2hmUQ1fID7ZHr0nsWYhv7yq6YXKLoE9
nMyRfbThdE9wDfotjTL77om7SOt8ARnxbDif459DfwbYq0/CRDUXGDT+BQ2h6yT2SIEDETCA1Hmn
Ck0MczzrUxZy+Pk20TY6/DMDuefNCb//eam/i27VCq+rnvptYn50MJQeTqErP8LVF/4GVEeyMUIu
yvZ1z5wWU90FCm60Ep1gosAcIrDRbOi3SrI8ruDMYggdt3yWzDiHH3RcDxpxJM2jm/xw23A0/RYF
TIkyU2PVqa0mva7X1gYe0qdQ0Y/6Y92PPJ2/b9Koa0nS9hlN+NJrOTlDioD6cK1zVcwPBq9S3mIN
fHcpo2OUmNxKIQFw3NU01IRmRZtrachif0SLhI0El5ejkBDFfhTLzEfke4r7bSLlgVjj/NSYtO9n
mP2zpvjuch+zTLqWKc3KDccY25VXHTjx5GVY2/gbpOj5Mtg1sk0RT4GaE/7TiEy53wDlIxk8jHhT
SMWNU3L9L9LFIQC2CJAh2FrQ3eK6E1sR3vuTVA1dX6A+64PeMCsmHmNITDcQBBqm0HBAIIqUTP1U
KuYVlG10iE1C2mAb+Ql1eRBezrbIdWi1/QTHQoyf93IBlcSn0NmZcE/0tlRkNcZOVwlLjB1sxGTr
hVeMpAGp1aEZEZdUMKB2EfQ4scy4Kx2P5LCE5feIkr5FYNQrP55Yq9Simnzdy0kwcfzbxtNuP5XT
o2bf530SFxQGtfRaIlbPQ7IOiE4NGWy+SLow3UDNXHwOmdJGmHDetUPhzBOCVgZC/SwRCAcogbgp
+iYCctWM1VsSQdwW7Xij7h2HUqK+0QY3z/9+VQMtcyY+JEkHFpP1Z0emRsHt5FsdUfDZ849LBko2
Zb4F0aORe4NgzTHHYpweaOZikQRwxu7nmGw0QloPLkYnwYeyYW4+W/2KQQi0LR5aCnfoaYgGt7FD
aRl42Clu4yHj8NnYaufeO0JQn4k/lluD0Bs5LNE+N5SZ7TsLCdKMfFh0ctlgEkF/yykbz/PHq13I
Xq4Gro2tDvnHu9ETVQ61dPbzuUx6SponTUMCejpqE1CrSQ2v3UKv+wU9NnfVG4uN8psWYV73JGhP
gO+ORQQ+LXlS9EWZjaTcwylfkf9d0Kll5NZjyWNqGZb1HKPeVXDDKBNztZB9oAQUEQPHLhESvgmF
XimooWf8QHQDZ/ZVAkKQ46E0xE1nLSL7PYbGOqzeJcht5dRAcF40lj43oXGly9Ms09uzZRtI6RT7
bbVbSOmo+kCYFXl4MQHKCoInSX2F7ZeNJ0GQFLA+Q9Prl78i24JkkwtAvG7bMulHdQ1j/xljdIPu
y6ZwPCOg0zwk/sMyD9aM6Akwiud9HLrGq4TT5ukPMLQPuH3e8KuBq5Ju5NOu6k5c62XlcJXXAKHz
WC1xMzBOl0FFHMJ+d+Wdg7WPoCkddqJE+4GxL5fpqhlFLaD2fTB4VTrR/Fxj0dXk6DMqRYfnywbX
Hyax3rGxVtH1j4OmXmvjN/GfdQ3dct2s3qGNgB2u/V+p7OaaqggQtMOJnsY93i4aZgMV97M5AlEt
1Q++pzIdtip7L+tBjgutHpdV4lpm39CgCv4dwK1iWIqg0zj/8A9+nLBfC6Ad6XMiX8fmK1D2/OuC
QQqQ1MuJwNCBXjySlL3A5dWQ5rzevecJpz4DRQV3RcEBbf3b/pFi4TJExCLbw+PqnOMljkhGLFeD
lBJ0VO6D2uTPwUgya1xwNS/6VH2Kn8Vdv3sFWsIhMCiKImr+6h8ZWnUxLb0WAgXkTYA9u0hXhAHg
cMgB7JwgSp1ZB9XNqSYEJbZxaEvQBQhq6yLkJy0lJEmpsvJNDXcde8WlEZh5B/Z6VAvPCE4To3gs
Mn/twlTSfN7OAII9fxOKXoypMn+frAgVqV+RKkIuzROo4b8YqXTTGKpp1/cjYyXcIn1YSJY7cM95
7b/zO6d9x7TrFq2g6hYMM+YAx9eM+Qwp9WFxMGCUtgfQywcsn1PlIlScL9alXZhV1gJnFd07DKa3
cSE3gfG0aJ2OIPCEE3iCW9vh8a97JNFHvJrLRFCVOB2Yj/ikSy497V0YRb9/2Oj3IHIBh9Rbh+uW
iyH77rILIMpTzxG1Vmf1PQLuhCNrys7ikVb3rcJHlg+u4geAKH6BSI0F781dsbafTGiLXCNqO7qd
Hz8iQetaaB9BDc1EBMud3pTPppgaglVYK2oJwi5x+5Yocfpdif4CpzRf3SttSHGf4zoLtx/1A0pd
vvhcWsMNIQRUPHxANMO2x4v1qTSfa/lzxN6Xct0SE/l1WSjrCjvzke0yY4bAJaAp1HX3uZlHyLu9
fyJF/zxET8X++9z8L24m0Smv8u15jC5UhZRXp3QuW6i8ubL+p1cZfZ1dCz6Mo7lMYAGkaXmiwzcc
OYkqrEyN7jdqyO59GexZGbqkowC/PFQt/9XD6ox7ikQtCsd5Y/yoh+xNpaXhC7eKkOP9b0jlqqcq
U2n/VoCI0tSDkMEFDKYdcC+ywcZg8FD2+MJRgaZ4vVxmUdLO5wgaC2VmvbWIvWgCmfRaPy7OMwDl
Dw07Ab5AftVuO9HgWC/SaxSr8obvkLa5Q7wJRtia1xGM3NF+5LLp838nuV7OkQvjLQJD8vurbYYW
5uP36iR4U+RmC4s2/aS8RDgou8r5y/ccq6QiQR687kPx3eC8TVDO18PikGWmsaWLtG9HL89HVG7y
uh1x0EjOynM1klAgLl9Ksi9/ix8QxKR32oq2VBq1zM1Ls5ircvVD/JJ8IU6F1vAJvDf4Wjmf3Myq
s/GLGihVdPtTFT/e3FRYuqPgpxT3AU21Imd7HY2nmt1/svmf1XzF1u5amAoWenxhzzRrUhPVgl7d
M5Hpaj0DXDinmHsXbov+xI59Qbh7uE69fDM4dSPJdT5jTuo0fQDTkNblVWLAZOlcz6vMJOkJFNz5
dh1jx52ujlumX+R5oBDDoqyiUJLeaWS0weyQ96XVIRiqRIWL7L2q0/zz+iicXbPBLt4z0CUAYJiK
eiwc9FxQnsCYDm0Up3KsxMsxPM9Do9hWF80XJXObXOBEzJ2+cqLJyP1UCNSVEJxYJOw7RbTQcUI/
MDzAw5NZ6iNR5Z8kywyP/ZyjFhFLXejsib4X9/5781qRJG+B8uSE5WUfzxdpkgqPBJzL9vpoo1WU
Du185ZGFVMg8gyhTeXq1IgsN+cCiUwWPSjUgqXqeKlH+VyqcZw8COjvC0++LDqa5WjfzwCjkLjdb
wYXoWQSf5zK1IPi0+dHQRT4xU1B3uRUxKKenOZEIKqp7NchKQTCt+hxvwfLwnvLi4nTAkJCGUEff
JCE7l8XOiID0TN6VCVLKCG/1bDENOcZW5eDP8MC7gSg4n3RJeguJajQoEjfrAZirHu1ib6rnrCjX
bavkklpc6YtrmkF7lBT8A1vN9ZfXH50LBIrOKz1WVdLNCKIcpGNfZm2wq21fjP97RnbBNfGozk1M
YXCSYtoEHN1iR1XNndIZ/aIZGBICSHRo5HLGz7tCok4sjXdlme1WSLNn7fIkd5sbDmTa8A4IoOfC
3AEX9wwhYMoV7DMEB4kfyiNus1KvOr7VDPm+YfGfbzcRq7kUC6a3qdckwg1NiNf3Q6HB3QVhaP16
u8pnc+1ZPBKdo4cgPQoLEmzSxu/2b5QSsL7pAwbDQ/7u6wzyuJmOVwByV9euNXrIsS2YtqvSZQ5+
kpkBCi3jOQNtaa2kvPPapwX6GzMVTuuJoJLOdveKyzJrPvX153D23p51ZCaOGGz8S8C/C+fXQI2O
X0QEnxgqClxq51UopsC6xR5IBpI/Yxx0myePGPOxeDmFBKZ3b6KyfAV/lhM5UXazgs+Sgfzi4ae7
CflY1PGW8lsNQnU1GYzvLgEbohfJVoMvNmIEaKixmUKKyV/Q+gPEh8h8D6GJMxXBG2napXny+77x
MwsTGt+xlDoURX0k9exOsryN/H8jM7oS29gOhiNPbXRdeweL8VgsgpZTjUNPFRcxGA+2cjECWGer
fYDANnDM7IQfO1NUtREGswp1w9Mzx764nO0PHNj5fo5Y+OeQFRY89oXipO+kYNgBWTGIPgOhCXJH
mH90vPHGTu5msKoSS9w9DjpikQGoQg0co3Fi80GjFKbCpjsR04B8CeJckXNhhvS8nKn1CNUA8E70
vcrcV5NrpUaqMihd3MTHPLJTlpP6EZHy/W6j1S+nb/abFgVGpWrhM7JD14qhDs1xsycNbHoqxnEq
ui6Xaj6YuH8sDCzUXlMlmiJyg0XjwX/+11XacgBo+ijJItaH9YTuXEt8H8KzZSA9Vx+4SxO8UZoR
qHsqgRdS7PpB/f29cL9Eym4vRvW4rcTev5QJ1Qfk2blWDrTg3yNsVJfephECfXDgCA8TIuWgOjP0
2B9D4iFFQtAI9uNzKpqPRIj+za2BNSlKf0BMFZleZD0f0+z7JRJ6a5QHODAZRLQeTRpOyGWGL5Ah
cKo1hCVQPQoM1DfWRpFg/yTD4pXGBq7XpTcpIgNSgr3VG4FR9xjX8C/UFJrOIpVhn4L0cSPLPAQX
Tix2IR1hUCBLe0CeOmzP6YExxFVyZ9UPFfqozspl4KXbfFGv3lbMgMXjK572KDMU/cLVvJuMPdFw
OoAtY/t16uBkOIIf/0pWhIR2P0eMbA2YS/AF9k4O9aRP7/b7Ov6qNgyh04kuCx+qrvPQRaYvTvqi
PkteZeZeG5Rsu9qekWHbhXCYup/R3JekBJVUblDp9ub2Yk/NBebKYqOxXMB5sm9Z/p9orbgFsciS
BhwPr57bT/+ZHHjbWoDywqcMIrA8sCfnudLofMw5Emj5B487ScCNurtjvlwKA4S1M3kHtZ7PGV3A
d1cycmGkgQFr3nyxTYsyRIovzBT+GRMy1L7NJEclW7T7DDNegVegXLJ3ZA9nQ4aUnsWTI+1cVXrr
lOzBBiZIgucsvrUjPHetV37sOKK/5O9nADZizPG0DNUvWB7QRpFivXYdcyonljBr6DNwjDKCwdDB
vhyfhqS/EcQdHu42do6VhpryWhS2+SkkMm9FSSijT1AT+f0PtRyjxw9+9RbklqpRt58VhvZcev3S
fWONtLSVMit4NWCOv8lPp8cVOLRV9yYCISM3N6hQpKkJaeMTbB7sE/1avB6sF5BoCX+vvJe/Iyk/
QX0uI9/fWELw7bht0N7ZFhfWAMw15pYAyKEpynpO/cZCDUXzgC5klqdmQgTM5CQogQTBlfk643ut
Q5/jKnNVXgBsyxQceJrrNgIJFFDrItl3haUjX4aOBja7olEYWiR1n9V3mtzzrvUawMndjavCQhIn
FY3X7fW0jtq8MDgm8eIsD9rhI0I549YbQPFbIEnjfZG5Jf1YBelDlBQy9AtqpFSkhM2i1zM2/gfs
o4lsQMVVqP3EOYKyzukASSkZkUiFQXT8yJd9hCmg7YUkncPMoqJHbC+ZA5ETT4tGyMd8h1p8P0lD
TIQ9JYzJq8lvpr8BYWvvjQNTdlX/FzYHzGdtVALc7X5rAXZiL1AIeZ9aWl0k/z460pdeCtbWtW51
ISrnZCapb2YygLQ4AVrH4LGVt34RPet3gdFdx/cFTREkNL6tCZBuOgwPd/loZcPyEEeAk0Ui5pd8
nFgfCWGeHE5pfEdqhS3+e1+ALEesA7YAiN0YPas4nl6lqFmU+qNtBaPMTq8grSDr7Yir3FwUu3co
TkqXcpFQXqhI28KY4iHIJco4OAk6+4SyjXYx3/S2gf/PBEUlDsT46pLmRLMVyQcZ4FEcVKWlcjYQ
G4mE+i/OuKDNcaVk+fncuH1pcofciX71PjpkCJPlxJLtfV1Ds4OuwekmWu3IqUXdz3MzXxWCGRtY
i+zJQDLgrDqyrH493A3J+CFGkKZJ0qhxZKyw5YjMUX2GaDZsEjHvChgxM1C9EYDIKNHOf6kia7JX
m+adpVWOOnq7DduzfLelBN/tWBtMv9fABhGnQCyyyTnxsP2+Aa40aDv21NSMLNLc4XjnzDgNiNl5
StJRtLt/oP+TECbstsfH2mrTH2Zvy9GA40ovMvO1w7xd5KWYstBCIYHRs8gPlhUJZO62uwBW49iA
yMfqTfWFvUoILXqK9Sl+3AzmpNFsKlu+SG7JgjUT73wh6wAavuB9+wJJVZobD/aDtzva6cBom27S
+VVpe8haqg4jg0nc5WXgDe//hFkma+KpZZm1PAJUBP61bnxMUFqdko9ZsC1IXzk4M6qY/tMgu2kb
GVZRrnAxCtZrEAIFEZXIBdGMeAgXq/xA+E/5SOs57Fh8xjAjo+ZRI5c1a/t9yGxQOfV+gVwsUTAr
LhnfeNxzRtOm+LTN5S3JEvb85vhNSt/OcVGHlCQJ0rsUpXCPF5HXDaZG4JnI2aprUOMGlX6WmIiX
9wMZ32G0zmJs6Z5UoSMQcqydSZ7IT75ICardryx5dKqu/FyPZwKXMp5oFABvYNKC1vIuDhq2Vyw0
BRYu/liHE5HpfmlWU0jFYM/onO42+d4RlZGyE8skRjzUnNqqi0WiYp8iIndzCV97Zpr3mgjccbKM
8QwW93KsVf7+4KdWpUtZh//+X1iVybCPi6VTJgdFfuEEemsESoVbhJulHfNre9NJHb8vd+bU8X5/
P0k0BGplmEeK2jgWmCDLKJPfA4Zo3Y5ih7Ic+UBhqs9g5kpEwbojK6eRVdNT9uCrjdkusm5Q9mFC
Y/RvSm1ABL7fHsVfOdoIboM3ooOQ934PikZsc6iPol1ZkfrZntA2cc7+2gWRH44YQwljYTtz2IFt
emGHiC6Vk6OKnwGhmlIssEceSKNBdI5otyLNJa66JUl7GwcIQTmVAEQGSZS+4XOdk/NpIJqBmk29
lYmmwPVbs7Ze4Byh1ozVrXYyHGRQW4EDMK/rWk9RobmM3Xg/ZhPSsj9/GWNuG61TYOlA5qUCNwix
wAXGaMpNUmMMPv42AbB7bORZqY+GpTglAb4Q/HDoshsenkF7CPedC0WN8SXMajO3lsg9yVKKmM2g
ffw6zKgZc5gTR5vxu0QAP1f8/UvYEb7xw7TQ9iJo3kttUmlYhA4BQoIytZWaSsvYrwov0BhyjslL
fGeolreCVXCBphmfUso0ODKPPNEdoRsUVFRwyxCxIcQHPrxBxvwURD9ZvCSq+PQ1juueGOtJMl9q
0qbDCx1JqVSRqs6qnJUC/ePkP7NDD7v+OHPhWAquEOIpLz7TLkPtmEyiKHBNnkjX3sTtZHkpS7Wz
5+IUpdfgfSDzYwCRERqeQLgdM/yotV/D3CeGMB3XDI72gkHlG5Fq0CEKkrymBnWOMrhZhYbIy/NO
mL7JjTQCatdLsyGTgqp+MDYLycPf6NwSG4G9cTBEKRfhUd0dloEk1ZOgLDgzSIiouj4BHygayTKw
jaSTs9Z/LxhJc978hI3DwP2woVOlGmfh5YuDSSbFcP/10VBu26gKbyAJJ5hNaxCdddMAg1/BgNFu
h4hATkaUpepX9nQWIoh5FsvYX6ts+CGRP3p9/n78rEktrcArhspxLeqUnx5ATJ8j9AEHLWCIPUeh
SK5IWAp8N66Q4oEdp1ybdekd05S+cSX6zC9c+71W+n1k2fAh8rBQEftvsanML7DId3UM5afWZuFu
FjBZGk/2UNgEIXZ9HJnA8gfvpHTvjMkKOSC8IVynK6CWtXGBIODP6hRn+mXDnnGPCKt5zsYJovDQ
8T7UhElSbpKNwPxtxhBDLQdBIb0VJEmb9V/Lnd7FiWn5pci6OvQUw2SEPwBUWxXS9SYBA+X0Kwhd
JDjY84ZYQEEPN+NS5vVUKCD/cvKUFjB7RiGXxVOLAP0FdwRCClJnBcGUJ78XTte98tYzPaa31uLA
To0K51FPQtOI+jI7fzfFsVkTYgWjz/1QYWChthFj66BiG1uIOQ8y/2J6p/DSOAqVQm9nglVLhA0L
mTN6WveBkGHOhKgVug32DNfKuktwR24EWKWdUYYHYkW8MAQ3kKpZwEjKM25L++M3/KVgxM72n/Q+
R96caYtwPEbwvWUfyufze2NqO5SsXcQv3pZGVKoQKzOMX9sCaFejnDmL5JPa/oFH5rlXPRaMrx9L
tomq9mBiI28GgwPvtVytBSAWBOpg2GdwsUldssGJlxX4i3LCEn7SInV4fcuIF8HnncgYcaFFziBt
WbUtlObGAO3sfhSMEOZPZ9IQjotutcpEA/4P8mSjAZXQr/qNoi0zQP7TeiRiCBULyWHQcTjaR5/w
3dOthX3BCSvlw9yGJTggSQ5HWCwnvksRZ7t6Qb/K3lWsM8hLeiaouLUj2QjXpkfzJhlE041LNBZ7
tv/Rbsv4E+lHL07Ma4GyOZr7Y+AKfxnk6cx0kswaHDjIV0jP3R67ShLzJRTIruupUV1wNRkjSfCe
q4jnwQWqocvYV/jjXTucZVNykRZO4NXmN0Qkysaik1Anr+7WlUA9iYVaF97TZNyjDdJPl8Bhkx4a
8+chFs1rSpBxqs4WoBqTUeqscu59yPExsJEA0lSBOsYUv8u/RBClktAsmK7t4mHk9poTSyN0riX2
feXTe80TkS1eELYNn+u7vvAaE4edDTJS1BluXC/tSzepsjoWen3GAR+e0P34vbyHzHOrTrDhaRS7
pr6F++f/nM5/Q8cQPbupLrWGLKD1/JdnAChoUFiJo+2vgQQHvfyS6rlJH0kTLhRF/Z9n2+VjCbsf
5wU+0k1CXJ4ZwNyjtv5Li59VIEva8hyx9o1GVTdU/L4igfOB+YBzNo5NaARCQXQ/8atGqs5ifk0K
P/GEkfzo5avA+5Hgk2jElZRyyodf5azVrAOS1QebHyTPTjgvqpesvZIF/Y/lJtDfs9NIm7T+a+5L
NaNrbTB2AfRjCDxORAMGi7O5vA1AI2H1nDQfgfBNo9z8qSoiqE3iZ5Rp4lqtcretZVrkCAjfcWeU
+DkF4Jmjhq0N38THILeC3/e4Isig8WWmXneSeeI01AtvKBTc+E2ASNScZ65ai+QYRdOb96dcR4V8
zkofWIK9bKoHq/k19LjWkYJuT+XgK15qaYi5Ic/XCAjcHbHfc0+brGGYuMXX/ooKVTaujZWebMgE
RBlW9FKlCBO2lqpLJ1hq7idnBdowed/p2BXYLDFgsQDzpP8h0RSH2sqEaussaqTrkAOA+FruZpdw
dnOM6qiYncz1HnosvyJp2bvF57SRBxFZYB1GqL+gSbeO5yglE8R2MP60xuK3S5dKxZIdpFASvEDB
ijnURRKe38/U732qKRP4FbE/wCcYQ4/3j4M/qTYifF+Uy2q/nVqZluidnty/WpUO5LiP3wqN2gA3
W7A3L2DIe0/c1fRpSkKX4P/j3VMx3RtKKwMS82BUqTTETe7flv/qs3a9irJ48DBF/kd73XazbxN3
Tg+9WKKD6ZODURYTSH5xHqudcufMy9sPor6XzhfGo6J1kmrKqFGEsmv0ftwlG2acoOibDR1UwyJi
6b45Ett7101EF/vTQTIWkSSYKLZCBcMCSnJMedd5Zx7ODaIYSZALmBPgDpeM8uk/BcxgKIBLrv2V
VIkhJOy2CmK9MaAPfUK9p9HOxtAm1KcVlc69HdL+e2rgbYIrwrkVCnJXm/uIvAGG0Celtcgi7H5b
XwQ8jVr6DYOEuH6y00bTSxqfLaUXIxY8qLiJDWe7+1NVB4oiQHjueDH9OS0uIW1mfMzgfmEXRiJa
BWTRXeank2PKsGeNlR0izwbMfgP0pS0qsbdLKKAGXhHpbOHVuvoHwvfFr7JYD7yam4n/gwQLuwOX
HhwuH9fZQNv5KOkhX/p74D0wgzvTDII3E4pMBtVay66kNFPGlPqVo8ypRw2JcntyE5SoqoD0KnkK
EX+wMf3tCLj1+hM0pC7UcPvQOL1RXC8/pG1j3h5v8Ehetp1jvFaZXz0F+cK6R8g8Zxyie5avFtLf
Vf51wnrDobtuUVeadcbpzlvk7iy7uitTBmN4Rys3R/09Zqjug1iel+72hQiFg2jMApNsvbTKICZo
U6eNMXjJcA89nk/woavxGHUKsg4xJpkPoYrsKc5aK6DXdJPovrk1tsQMPsSaBs2gsXlC/zRE7Wu0
LJkwQ8YF7D2k6dZpuCqGA4o4UmpZAgeTD0jAinviAVIhOwctuNaTo+UJv1e+KxKtOe2aK45CWqG9
a/b9LJj5mnXKY23HqtWy6VAJMmrJjzfQuwFv6R8iZbSRfHx9K1L/n0W8UoicyzZxUarWvJr/MPHG
QttX+t24mxfipUBT0gZ8sidC9k4DyJ5GgRzmUYdEZv3iI9pLKNkJkK1Q5Ufz2RgEzFXdOLHm/2NY
zSl27J1Sd1Amm354r0BSpH9eEn/aWbJp9y0wyeUJRbr/q6oZRM8pjbZHa4dG3uz7xkuX4GiCZaFi
//21ojPSvPnh3kQmTZZQiHGucH9o6UlbgEqqU0Cz8AqicmuJroXCEceSheXjxhhmf/Wmf7ElanmH
mEHDPVl9aTGFpwI1d10htfdfy5uPASDdxWGCiqXNGGqCltS9swgW+uDk0fjPVGlYBhbV0SyT0ld0
LXZ9hEVfzguAsd0L0ceH6RBO1ZMB/FLUAkMCPgn6MnYsmCHQ2ZoKg7RdQKZtNcKMEIoe5FgjKi6A
hJ1IHyaAFSLrMFANlEEZsEsqbOYo847Eutpx2kbmz5tUhH2V0JV0BheZUN+tVeulVKMKJu0CRWzJ
u6M7ueQeFJb98NopPqUYaCrCffaKrrA8wHhaczftx5uk0ymhYe20FyzOp0MQMtNXjhnrOIarRLaq
fZNKQuFgZfnEh5IjH/NKIHttlgVqNBCypQ+g4cN9OYuoGjD4+cbztcqM9SJBeup+WWjHJyDmcf9H
M/Vtxe0eWKnr4cEjRS/XvVuk6pYWe/CYzEsF5LGo7XE/Are6cNQbkcvTEzIVCTZ+O9YNcc8NsFo9
PBXGVL4ElHyDHZBomLOnN/QxWrVymPnIH85TPJLQgdl47Cj2JUw6ee8xJF4+wclDQZblPxqrrkiO
/lrRGk3rvybLBr9HlSn6t0IOaYA5s2KYUBxnzo/ylqeP7HiU6RdWE5kYwxn9IBvgX/ilTrFRXPgV
Hp0PR2y04jl6lhTm+cpv43Ky73ie3W5SNPxOySmyeRHqs6tyUXkQvmBdoU6943dsfRKi/2gVjhmj
BVsQERatr11YAYxMYqzaAhMYHbkmvlPcVAdoXkDIR3wY+5KKNyOm/JZSAhe7t913x5EEdJ7ZPRf0
dsZJ6ju7q5kyo4PKmDgmbP837KD8/C7VF7AEv9OlQGFzpNai6soGofbVoirVw3gyh1MetD9asJ0n
tdvi71faC7ricFE6shWrTVlwWzpU7OzKYaoGUF/MjjydTsJe/VwuaL33sHp46G/9daO9TAmFioB4
YBU3pAwOTCtOEAlj1BVZATKTJUOrQAyDoFU5/czOWUmK8ylbMDVRunrqhSEcW9ZE6jghqU3RGXPk
O+zb4qX8ujwVLjh8lGY3zwrvXhT75P2iYuVdo3kXux1yK97iFLtgn4t0HkfjfJm1tQNMNDjnH7h8
4ZJk9jyjwfqSuTW6r11Q0xhcxD0qLkjjQdZppSOzrZNTyc13dVVfclUTEuvRguq2B/NeYPMxgjRh
ErcmG8cjp+iIvaB7zdhFhfNKmeMgCOy1xX/ywDnKBJeJmFqWpmBxs55sgOFTFQtaTojvHCQaobvN
4Q8PzwW08vLlqgG+gXWhknpvI1yEgXk64cBbrkh2c0xRiOVUBQ5wC1+ZRwKo9VVoeoziyw9vXnxj
quoCy0lShIqhsBREzP+F7fxDrkPp9Y/Ggux+OTX9/YUwY8K24xYg7xqbnhvM3vY9oKBM1RYIX7s/
TH8oqudzQHOGEojOTek2hnm4kCJ3AvahwXYINdm/0eK85XgxIh5D+RvwEFxs2k6698qGotKpMRXU
GcGXHBh11hOXfqJwgDTzihkjqNeI1C70txJ773lWn0Xc6WFF+N4FgHd4N80E43lxhyBCRF8gjkex
15fSFWXYpWHvk6UeKGS0U4WxsgGloKXlHVLVxYugHE6d6tZaorn0IK5SSvTUdIfjtu9nOfzsLjRA
/rxC9qQ39xcWcKkbZssvGfRhgeAHpJbS0Tn+Yhw8bGIbqA7A3uzS9NLxKtaLinshkoCfutcy6wsA
IQ8k1sKp2ypzx2wllWh6qvRQYtPlzSR+hQkWuP3M5ZmUdeeu9z8YcYSsDvLIVGPirXFQ7k6xtK5E
2+FcYGbKE1uPw23bf6q3hvU/ZISLEiPmpOYe/QQxws5QHbM31AycMDiQjWUZrE/wPlOGx+Ok+oM7
I2CbQ/K4rSYdom+WZLzXfQqrZlGVvjOFWogizqEda4Q8oD1gUwAgazeOWNsa/Wh1tWKBEh+nULLz
HWmUdTd/+qZ+mY9CFpUJCY/h6yQMyvutDy9MUFtU1Mnc+dxpyPcaUZQ3q0jMNpzkxXK3dagvTy31
n2XPI1BNvrk17RDzAjyGq0SwFU4Iql32k0xckt1i4MhKppNrPAjLT+QMiVuD/Tuvd+WaAbsgTeDa
7k4EIVt6f5PZa3vCO1ckXrgCIw4C8DKl+/cweY6BmO0N5hvca6AVP+nSQJ0FKGHIpBZmgOBttNSN
jkLbn9FWA445H1af0dfV2KNi7PFCk2ySxJYN1e9YoM0mL9XxCYKj9LvBLcrEKkeRf5uF61vIOSDn
s+EjqcXNXpUUy+ZQtkMog0YMFM7sr5ikFhc0J66sZReRBNx0dYIhqMdTSYuYsS2kHjUIQB5478Iq
DTEfHaSzye7I88t1eEtWnGGuqSnGorOREhtTwSjeW+i4guFCqaFURSQuojPscwtDVV/hzqc9DQj0
w+F033VhfYl7dk9x93c2uaFk73qFdJ8JWNiBFZDOIfJwZ5QUqRYG5hmVqt+yD/gDTIk3xdiKm3jd
byWBYnMlgxT+/Nrs02PdZqXIgAMVwiRSnNP7gWfO9En2eG9W8WPZsuJ6lyjPYIhFouGie/fQgtbu
N1tDURs1dBMkx3LhdHYycvbMSCFduoEjFfqs3gNbqUaHtlxnUKY6S+KQ+yEiIJZb/Y6A3vQdlEB7
TfLtXvOOuTIOaPkGkBl9kwj/TiZplRUxDP4rOsNy6XwK82ZR9Ll1iFcYq0mgcTh2+GoX1hf+gRm7
WqiMRo6B5CWzDI7Ui92SLy3UnvtjOUuRaogaF8aBQVCik4Azsy4B6Lq+mANJU6HUl8BQpYLT0DAQ
1E3StpIIWDWo69Nnc7LFUyX9afCspQc+7zgAizkASTOH8lcl/cWfekQzQRF+BYVcNZQHteqZcbLM
/kA/66X2KdXJhwBA+FhJ4WNHwZ6Cv0qmB3UurMvL1/CVYMmXzorVZdnYXfLSpl9vz0NpkNc7AzA7
/SCcmMLgzl9uyOSCoHRaIQjamI6mo/PdnJmNlcwaoZiZxMP48NQJZ4oNLs17k6/7bnun48S5Cy0r
pVEwHAiDiRvVQfaWETxFEOVfR1l57q+Kvlec4Pxc73vFwQIppekiTW7X2pBP8EnbyZI5t427iSCl
usqXpFcQ7Dyj77oFJK3U3DUp4yVxZVZgepkdJBGEzI2665QWGkd9jDx/YPyxZPuyEeO9xL5/evyr
OgSjpgCIOpipCL/xO8Nqyea1c9v2s3apmUm+VRsZLx1K42X955rUxy0i+z6ZDb4Ro49WvKumgfIX
PgUarhxqr6qvA3VPY9MKBliKpGunRHhoyvZqRNLTBGPhfLIaWLuSfDU+WxC+Yf8U9Wj4E0XkD3Zy
Q8ePu+ZV5DcbTkJhfXZbWcXED77R1NE1EN3TtvmKPiLPpk0dwWtuCEl6Y9pFDhzgH64RciDWnjO7
U+neRcql07+A4ekMdzqjgz+Q5f1Lxh1mxQYy8T6iBIYwsbRQmdu+uJD1P2xTE112rAE4b4qBTaWs
ezuNq3hKKy6IJWayZSjJhMiE3jkLqr79HzVP9ur1LUgunRuJJKXxUuPQ2Vz0fcmCl5qtuFM+9u2J
R5v9WSOzzg+YdZJIRidCXbVv4H+JHx8/DsB7Ysfd2TRWv7Jimyq/1SmuRiERSp0qAtqlB/Ue6Zp7
YP2nDxFOQ0lkWq1sjLE3bqVZ0ppt9v8SylTTqcx/a9+DRY8HRGuz2ZUEexVZVnrLUBrIM2ji5tH5
2/8RV48MbHHFCX51U/RAOrevD89Lm4+heyscnYlyvnmmV1Rc8oOskfdH0RpH1rneovDbAOnQatsT
8p7McaqAZV/7Bn/Wy/XZ8N/tG59VVJA2fQyLW3Er7yRjn/cFrfN8vzCQG27evOOI3ipp5HRih8iR
be8rk9W8ZddEkkQ7mcDExKyYWiDj1m8qpAuX4iMljGeC5paUAaqk2KWFeeNeLVmWX9ozXkrpBcto
Bel3idyOW90cmWXqfRPKYO3otxDh0Kmb/OZyG4XVdixfqepfgc8KHE4IwlC+4QdFwkQfKnkZxMNl
K6WPyJX/ooDPJnvDszlytpvOlVjcuT/6zcFRHZuipbF/SvfSKPNmWTyB1ZBeg8Sc7GH2+i0SrDDq
Bt0pfVofod+cxpLvy5YIZbHebVBi3eXGncRLPhZi87EM1AOvJf0SvBeOBU2R2kFebFa6RDA7M8rM
ZtmRKTuX55oB/zx+59VFbggWC+UQvLfVA2nw7w+Di7nRd6fmJQi0j6hdptamEDA68pyA5RMxTsoI
9T9uWFqkUbtAMIUpQmoV4Tx+Rgu0SipxdFzOh0j7fq5n1MfO85O+xuDxUlUdzdHF/WMDgBU95z1W
p/1wlJg2qEB/M7H+sA9FkBVdB0J0ggOifB/Qji6rHq4xlBB/ezKEczLmppR7pqN46k8vDKIDfdIJ
LuUXA0NOazkTQGBMg/sBfN5xmuaLnz6LeqSJwOmgvg/Ghjtufk/njD+pyDwV09sPAT1n8ulMLg+u
XN9RocrCxXtfOlqfsKXmkUrK61/J1MMXiKt1qd/GkTFHoCiNAS4B5y+ZrYgN3ZwIQ5jP/pg75g6W
PfZUwjgIuC0HV5B5BFo1A1C9V1Layx686UWd6RKEVYzLc1670GeH+/fkSTg5M96EG9BoUH+atK5J
83uzbZBKGyV/NVXxDi3K7N3VRF5CU2iUZ6E1zYgvfyXiRFJnABc1ge/r7gw0wPKccaDh7C27K5nb
rphfl823VVfpHk7B2q+Pv4YdsK67//AEh0EHaCznKHvdrPhojRy5klt5rjAg1QM4nl1NmGbvQHbK
VdDUmblJKhaYZADbgHdRyoolQICW3FADYFM8D4FwD3Xgzwx4C1LcQ0giW433RXyVB5aUgY+PPTE1
t3r4Rts7pw9WNaqWUFwSF8yKyFGLuA9dB189Bl9gvXwTrCYB7BwRnFZ6rnMXP2/2EUmHthfHx17b
RasAyrKzdGfPSvfY4AeTLbM05eUHUKDsrcFGeAWaC2ukN7O81pormg5C+10svWIL8YyeBa8wBERr
bwyBuhOqxYuXulbKafiXbpAw5zVcCXZMmOi48oTyHGiaNDp9AuuZpnW/i/OXc9VdNNerbdFPPBeG
mpQD20GhaU8qGSAbrgkXrjmb33/ML/eu0HWoJy/7rNMDRC0YltY3MauzE8Faa0OqgnyjeV6RzNQ/
EGPWguhsTM25Zl8PW0d+5Ri5yM+jIXcQAI3b3UwLoknPP9ULH1LwyAH249VNTG4GNSM6RRJdflJi
HEVsDXqo/wZoH+W7Wn/nbUyNeFnYXcivBuF23UBL0KPDpwekUE1oYm1jeYgHHbvOSzperIxelgdY
FF32xgymZRPeU4k5G9fe8ChkyagVcipk547Q7jTiqymyrohxT9E08oNW7qsYx020hj0/AjWc/tGr
RFffGMtWMPVSd5JRX58lIV303oXELFOEwITTCfKoKNgEREEJQ2JCuT+FsgBTC+p349kQsTZUmxD8
2xb2cQ7UfGVltOgRTMo7nS4TaBWqSQGrzkSdFO05NtM5x+EKdkmjyUwo1kGEdeR4MWpbjlI54Dqz
6TvAwWv6wdhjQeqtqcvQhbNca2Dg1b2asiVFiXOQjQ2OmfNBcyW6/681wkLgXupCtpU8TYq26Tun
WDRgGWlw1PvnYWEaA/ySZNc+JvNHjs4KnkHo8Xvv/e2O/P45N+aNwQxiL2GhRw7iNG3rI1z3dMgO
LOvne88p9hxUBT78V9NlTQr9bMiHkuyzRHkYB2Qtbv0JcCZuuQeFafvruYFnfKw4PUOBdM0JBFR0
+9DSZE37EOneCGMxXMIt/yVm6DaXMQPYrffS0Eq3wEc35bYBkzFeuqZlMFJT65z8enkFONoeA8RA
Jtx3bpq+uDY3sqwhVazg/baxAVrHW4EeKhQNYy9f39K+WGxwGDnvJ1tBqt7zuhOhfHUep0Dy0ax9
KwBF8ZJRyWNxNvqj+znH6e40QA8ZloXeFfrwrnKkp1sIo+3HO/kE90As+Op3sx5VxqARnCZWRzap
diNf/yHq+K0J3NQi4EcHxf/kaNRMramlFYZGySp8Q/sIpJehsj+twktKAYB9wT0K+FuNQStBfWUd
e9uh1m0I/t3Q6cGxwwFOUBgy7cLL3/ix4of5pviUbsrvRp4c7CysPOi/KpFT4bJquVKefN10GPP0
BRjxnakNYNp6y3VnvbKpEZxz29AI6VKsUIFMX+ZGPxUtWm9oljBsYTiSsPYyc8XVKavW5b49C9yF
eDg+x+8nuE6Xsnkgft6yWCs45dXhU41uo/fZCI3IfzkTy261Go39VzmkUH7xEt2NHFx+MrwSuVmd
8f13NmeVPHPSEuv75kIt7xxb6FlzZxbhQl5utFQDNa4a8eDRihIEeGaZ/ZFba1x32IQSp9ABtkSg
OTNT+JguYfVNzuU3OIyQxizOPnHwNvBWiKifHt3o00W+mCQNoxOz9Cjr3U2WLoQzz0ngucwRAgIG
ZUGmkom6XpBSEaCyD1tGb57WtPYBYcXpKH9w6QLJ1JUNFo2snhBjuX56KhKt1zwsGcuD2FOGXgcp
lGsq76ZnwnV+NbUTJtSmuaXJfqDodBnjjuJ03vmBFMWPBG5lLghoDcJTCnsudsY4JpLm9WXgMqQz
tQs31qEQQdjzMoow+CJDM2kS+F9oTThr8eIHxOtoLVNsuw+taaVf/AHslqBwlwVEAMYl3JNBo4YY
QGALl20Kt4lsVmPuQTEDfJutRhVlSUAq6VSgNYC7/zHsGsFg93y5yhKe6Yz8kBEuwipmJglWW3t8
lozbwMhHmC4DHQA6TpeDN++gFE2V2QbPAYBUXP5QXpVgnGGVgrk6omMY9W0XEwHHTrXdBn6SegR7
rHCQfyxJYO9pYSZcKKadVAVYGHEHMFQimAiW43b1oTv7QOXZ6PznCroiC3cZOM5492GqDO+uSrG+
egLDj+UOIm7bNPwARL7z5YcpiLp6KQaPVIQ/1Eo022vccK6WTAF+X01peiSv6ntDsFqDARKmTW2+
y0ATWHtZfuEK35JSJ7hShf8+yhcq3ekjFQ9hZiYtkHNti1EV7VhIurLd8YJ1PKeTQ6WkP3UzZQ9R
6HxFLbVLk3uAWGmEwWCG0mmDgykwlJCHoPVNMmiX+r/qLNEPuhUpRsTuzApNadC1/afzgiuBaryg
eR8M3lStc6xXfhlRWNqTd3vTNQm05JFui/gw11J4FhG+j8DE483J3k1keM4TD/k3MDh9pPhEKof2
Mkf16bQQbl3O9RiBx04XE929CyHjV9Kee9ctT8BdCO2plTILhqVG3YBPndfi/pqF2c1EnQvOXvGG
hftJRtzkEB57HdGzQ6BHBiPaNovhYsfXKbQM01+1zb+8dTWFEdt8/enoEnxzFjHXFjMqQ4RIAapA
O4yWQG9Qs6LwtkEmzHbR+gbXihf/rYUyVNzh5vXMKKWsrzy2YJeOrPpN6HJpbmTuDTDnBJ2DZAH5
UVp701a3Qqk3bA3xt3LZuFjywNJZXDaB406JX7mCsOu3Hq/S4l4Jses0tz7/B/nVTjh51r23EF3i
rReCDW2DmAHHpzZ5fQQlQmr0VO1xYmXsioJOSZa6KJyPMuppMbv7coKo9c3FrYGV8Fo9CU94QJ+F
mFYFhA7r4FSuW5IVxeWjOd/slHWu2MBvVt7mYN3GWTBgLbCWL3CA8V0Q6rpTNL8Ww/aL2x4eq1Zb
fFGLStoz7zR6MP2qXCqhkTwv300azRaFHEtxTSYAqvHSVcAV4TQ/hVgbZImoMZO/puFXgTsic0TD
d9tRAARe91wriL+4e3BNkuEPuRc5c7O5V1Wx2lezPrCIMgIy89Zbz1zsSGN67cJxaDnPF3urBXm4
mdYPereuC+e/XyEOslEUReX9FsUVo1PA+B5R60DtELLHy0+vv8fQOAMQawqdLRNkeoty61LGVTm1
lTWlYHmqkCIlgB76tx/G2P9I0PC6UtatgsVopV9QjVxCtdISLaGEhIYKcz/Wj7nw8UAjuAGnmWRe
WL6Dus3MyK65WH4CS/kKR88ZzM9Pf6W9u0o1gAzO0OLt5xkAER4tRN/egXW0ZBfl5DdlbkSInZM4
Yjz294lQLqAoNQm35FQk1DnMqyLwN+xU9dOfNwmG5pXsBDViNsxVx7QjdIvIjU64YNyGt+/XSQHW
ynCRJWFPSLOYxrZDA1N9+kVtBFQyRM6jEah8CVHjkczTRAIklKpxhIDOVM/qvOIazSZMloXVjpbB
+wivqa9y1q6dhfPrp3yDgoe5yCH08YucRhpPG6lgvOBmok0E2i5Guq38+c36lo84OwWKIhZbL1WF
0ynU8vcfjhjKkyZCLZ2kAqucqeSpNTlKDGyC83oLPYypYHxPh0jTvkeZQeLKnMHmU0aS+S3cuxqA
clMhD17T7taEw9Y53Q7rFPfHZDynn6LSF+M7Nm9w16QPZhMr3tww3TCxeNVCDy1kv9C9pnykCWbP
fNr+pMUnr04tocaPjcpRlQVHRBE6O30ARLBTzsizPFvQP3LFWQXZ62mhTlT92qLFScCgmHT0VJfr
IYotMzFMFg5TTQovM6LJIE9DdjCG/R49sUOoye6gARAaL8PL1ypid1m4fp3c7HnQ53Gt7dtevP4z
NO24/rMNpdArlG8jPqHS3chv5npApoxkinTtDqQaUtEGuDQ2FQvPzbasM1i5GNlzKTWsJCbZBOzD
Zw4x2zTDdSteF2/IyWWPsbJ8iXHmFSDZxK+YQMAzxVA1UR7znUsfZp5e2K72kbs6bz8ryS1+1w3P
wqrpV5NnTaDzUTcqPzo4KXGrdJprEmGwo4cLgD2W2P06+rEgG9Jw4lZQX6j78xcN8uNh5z0pMKRE
pA+QLHzGZbjQlp0BGi84X/+bfeEK4QTL5px9wR2+fsg19oSWLxVVzdPM7xqvmVANG+ZfP9nJu5pK
wogJRoqm7JGlqppWQs88rq+kOeaIPUY/D677XfufplP4/G+GbZgc1MiAXVY8zoHLdz2kkT6DyjXA
WIl77rq1d5GRQq44TlJ2UmUsRdqoYNysFFU4Br9w5nMwdLEfsPpd6My7ktPzkSfcAQgWBx645Wwh
Lo38HprnJyBtDPCBjtTERKhDqUqMDk3mEzYQnukWaeiSSqfWjcxclxKd5e/veE8is+Ol+Vs6ZZAl
6jc/hlsl6D54/Wb3EWEjqm27TErz5aCoPWbHWhnXMCpWVpRaR1cnJln62agWhAiOr4oG0779ej5F
UP9aXhp7mr/v8gLNREdm2ftJTTgBmzSxdI6Ok+Y476t4TQokt0ACcBTeMCuyQMW4XJhGiroxtdR/
FYT13ma23BXkEdz4LQYc5PPQ6Rqj9tHjIXUmhIcMWrWsAt1hoQ7mGHMdz03Yr7tFtuY+1oQmAdvi
VspNIayA5k9SL2OH1nIT6v6tiN9vzjXTbo8iiqg5RYyiV7RkCB+QKTGcBxLixYjCoXDtRIx7trc5
+DkMhmxlIOdjbN+ApOZEEaffNNqRwoXfM5M2xLY+Rb8cGeV2wEw4w+ZsilBUpidZX1qzOwa824+c
EKtE5CCLYLYllSw/QcV1xF/T+aGnj5geTJI7uaVJF/jcpjlebwr+NG8toy5fe4ncWpWgqWPhvYZ5
tvFt2lF8J5+8KG6g7lwReZB0Hq0AM99p8SoCElwJluWbxSzmlyBrum1pa9QeoJXpVQSnfbDDt6wp
iabWiz3lckh/2fpWFgdk9PjzzmPb+uygmeBmy6yXxg3qujv4BjFesJ4W2QhLZ6NuPVeBwPXqvVHe
gwpoXz+mzbhuTYzXbXf3i4EV+jACI6gaTAcNRjvrTpl42f+W86MWFVEtIIVe+ikvlboFIztcVfWl
jNHuwsks76XCdAG+nSI/kdSr5/Fn/2532ApB4jCCYBoM0IZO7Jmiyo+zdO1RYoeUgk9rzbyHJUTN
+nfVpyK0vPysAxL1JiFReCD7Y9rmPykAUtIsrkDMfPARb+BRepXvxYj7DTxS2AfdgdU+Vx7BGO9e
6LdhCxhEtfyKnTaBzVkI4g+dbsqJsQ32bfEUgFU9xOMBLw/cHcy/7er2lwzOV6isaxchyA9NluQI
F5fb9quN5Zr+EWxFLu+fBUzw4R5jz0bR4j1ICF+CJZYcPQ0X83YekxLwa2jqd/rXCKrGmtdrPN6X
ouxkCKj3jcLLituydR7qHXok50bgg3d0BxQQfQd82w3jpDzcK+QMgPvN0qkS97Y7BSmovnXH1LDD
ZaXUrrpGlE9XcnDwIm5sSYq0CBD/i4iIp9icJ7t1YBLgdBDafon2296RbAZrUOA5bU36jKmkTIVs
UhA72ZZjsSK7Z4+hQPVdQ3G8swnMLiJ0gsXJvk81laKTGh1JhdMcXLdKD7508qOi5PpJMAY/bZ/H
9+73qzSBoTvt22HnTQkFDdsbOiSQWYmZ2OzNZYxY8pna3zARt5jECw07BJ0aZxlHaK+XwpdkKG8B
zNS6iGHrguyWUvSQi/D+vj5n9a8TspQpP+EtnGANY/GPAB5mxcfkrKn2tiBLg+rxfuVY30X4Gurr
eY5TDy2wVKCqTjcazOTrViHn5X9ltKp5debisNp/vubUYyu3UskwwTYhTRhs6MFU9bVRs9Xuojbd
WtzKlqFF82Izk1biuMcMDi2nSNKsHyQ/fyI8n9VKLWYZrQGIWUU4Glt4MNrY2Q6/BPkpBIyaj1W0
r06tX03Yc+GchEWARR6q4NI5b726I56tlcm+jvs7otLzi9R3RYhI0GxqB39aGrmxbVyrypDO+9dX
yvawKwVgZercAICTYsrYpdsSjtpsHo9xLiId2dulFFJOpij4i/RVD1JQM/h5wWpUub/i1O7qQtYB
wCgDbBCOoDaeJlrvVbf/KEQkdQgy8hDlRaUuLiLLfow9vOZmMfqKw7YJCwieLewKGYIV12HUDkih
ioOMi0D1CK1hHjtd4Q0uybLYsC5DmemAeHSdBAH8CNSeX5aFnwmjYHlusmb45j9WhafwEnkpVzwN
uuTElz/A4xJSzGGNp96+2RBJpGsdCzOJG4Cqlen16bbMmlJOFqqQLKct49WK406oED8z4/yPU3PV
ETiTgnlerT4tyZttcJzxRpvtNgpsGvEb/j75u41T/uwVNwcDFaSO73vgcx0VyEDXlb+84sl/L6Z2
A3lNUpS+/nS1iL+Zpp0ZcQ1B62/0xbabMGvuy9QHfMunync66aeDPhrd0A974lUAl5hiUaG/T0I8
vqlOcOPHFjXqcPsvm4xwrmxStR0a9QEKNfxxmL9w+xxIXVzUgvfVMxl+R1Cnpu1ErTh/BNlLMbam
IOaaIPRxarQ9nWbW2ym+qHZVi/3qWpDKN7T8cvjRdcA057nUlHrjjRgPEVLILRiu8cIXL2PugyMy
z8B5iyOsqbkAlkIHDd58RFkAoyOWq6K1WTBxLHZtOE2ZFoVGGHnFFkv3EibIeu8nsnS7r/cP1cj/
IXfpZR/OzV1clhKDE0b9Mv0X99/jsb/pAz9v3gpQxkASl6non3zl+cmDAIX5dYz1X0hl3JuPl4Ie
6na4zO15dDHSnK7zwAvTtAYWuwa6IQvOD6Nr5CemB1y71aKPjxJyuj4a5GRPD+VMRwjJ9Bld51iI
fY4/2DBE/dTsNK+8MxQD0Jeq+Pye9/o/V5GEuSo+LVgnMxyzR4Ks7HyoKXQi0nKoRh2C5oGgG3dT
Fky5LwvPx0Sy/veTLFlwXGaGR+tRuPPH39p3NXwrMiuLe5kwmTUKjQlKEHOGN7ShpLdf4M0iUolM
R4OU76BC61wnOrJAIWZjnWwUnk36I5qgArFzBmPxVPHuu1KeIleIBnNhbTaZqKSoztwBozyO61Y3
uZuE521C6PGd3on1To8t/StD4dfC7aAxlgTopa5HshemOOeKkC6MAzHtqu4YLxTvoBDIjBSmr+kT
KllrY7SHVb4HSlghbV+IwR9iFJOVMkTMrtM4fXeZSfnccSDgdwwzk2wcsMwi9s/YabFx+5QqO7bY
ZSPucuXyq7tlvg6zQ/vLR1BgHlv77qZ+UcM0WVYpc5GILJ6PsJ/AbXDn1L5oseDKk9YAc3jNjysL
kz8ka5ZMRvpr+dhQS549PIeScBgGeRW2Jsd9FZlXQ+iFVJGYMKcref6auKv6FOpiXESbIYAl1N6Q
qNhTa4DOlQ3Z44wbvhocwHd0FQNM0n5Uu8ApvxJdmz7Y9rrlJNQJoE6ec+xbfEvzJJzZpvR6coV6
0obaKQ9IBvhCiIOm8FbxX7zdB5/KfaWEZnZ/U3+3uyWG1OeRDHbVOYbWAtJbqvlo2+oghrSfs2Tz
N/tM5/LRPjUkVnzTVtaC52gY0QN3fXdJD11wEqFlPI2dOGzjKO93AQlaKBdCgB5FvFVBNdrGny0h
xwnpov/Do6lTNQRPY7VZ124cG4q7uDmVFv+kS8rTPHzR1hr7GoBHJ0rr/P2rkjUNY0AHJfz3ZYLq
nOggub6LdBVZmjX2kHO7ZsP033YUub5HOBHWsLWkeErncGc9EVmQLDKH1Epy+6RJVEKRNkzL9OS3
q8j1FeMT8XXvdCrt5GIasTqeNSjTxquNv6cpRPqFfx/zOt/shANyq4X38efXIYVdsap6Q8dFDf8+
xVIN/V0MS2goGI9fx4KfO76ydwNg7LDoO3kbfo4hpuYobsIp6LAbaKCRyW8F5+ib1VFLibEE48t3
PIRMnoFIMQdGIzxK9cIPWA/od1RJxuWLAHeosKb2Tibd2FalnnMPiYXUXyv0+uXKqe7LMrGYBkKo
aP0iArnWG+9vw59GkyTjJG6EsVDjVgBu9sxHH0MGWxGMWCpDG6iX1ubclhQu5odgY8Sj/KJctTf0
ZRqI2o/A41WCnWSZ5eS/ljMknK8uvoV1llukLVmLj3sp08c05LPwTNNOr9pzmsdiIXVPpD9hJkqp
OYy6ybasCSXfzmEut+nnL5pzfRobuUER77pYWA9r3Q49RZb3tB1SuKFXXnZbuvyDQsX/miKiakgh
tOF0gf8AMokNH0tB3plcwoD0Kxphp3QW7MzMICODqw0M5UIlQOFYFXfC8Va/wOMQLWdV0fEWS/Ey
5BbuHz3DNF24YmiKUkI8whCEgUChR9INUB6EJ1N7uMMWNTEoaPLX3R9NxxLc5voR/RRMZpK9bEKW
oOEVIiEK6dymenCuvKP4WQSuKq2zvwOtU1F5Yu4G8E7BOQ6jMd69GOr1CCwoqW3bRiGwM2p2fEY/
YcJoc8dm4SXaNq5NOwq71/FKtGgxj4C4QdcUsqSf+CQYLz092yAIkdc3RjtVkCPXU46RCiQcCR7E
rlEHopWyyShxL6aSQ32bDqyXmNETTQzBiB4tWknIkBkN+wrTb/3zgEit6yf+St/SPtfW9iow84FV
T5s21VAz1VU14szub0/gGc2JSLL6OtdA/zNKqMmbSVVl3P7bYNCElnbFSu1vEhEQ4taHQyOQfQjG
3oSf3oRpCs8M0BRpbOVlClbCKgiLm+HVSjtsGFpwWKoTM+GIPxAkQBF7fCytXYzZHeHGWF2FWYCx
21YXy/PROsacw7w3woNZ+8VH0Ia8XFXlmmx0TpLsjOexlNMNAkRxilhXWniGWGa8XVchE6+xbBBD
M9jES6Ao9r4MmleYWFK8TiZ2ZoChw+3m33hnD7mDp5ACVfTAcR5gKC3nxgRKFIP8QbD9vTwpA+rX
7Lc8/q7x+0SfGKaQo+ay38tzJaDc4wcshdM9mL9IrUrZEyn0JYCmk1BELHkx2eojNzbban62ZRkS
QmPj7l/hyWbL92qmwg3D3Xi+ubHect5WL6gw5H9b1vBt6e38yyuVkFGtO74HIuMbaXqU57AYTtwE
FkHQ+LHuQ6ORLGqmWtvRrN1/NIbzhCQ5FjJ4vOjnHz1p0LOkUEcnwDWUaZhncFpenPmDVM5YYqmn
P28+vxqNlv+LULfuKZkAkSUScrwc3f20kxluuINKYJYkFckVIgKOmg9XmV7078dSjpACIenAH2vg
d4x9jkAfMTAcgeloiCxUPBGfdYlfit3EDxOkNPuVgAjTpmZbSTmxTORYhHaMjsHFsy3ERkFr0Fy2
JTDOgcVnsvvJRei9GY3gR4T1DfnYTH9TgpDaxdN1JC7lL313bnL6CTIXnJz13BWwB8x3iHxdvHRb
yjPhyh27KoaVDfgjmzqLWYxde/HtVLXgVI7kBAyTawf/37i7WRm0g9EWQwtmYQqPhIb+JfXOMfye
tPzGLq5Djq4TFm5j6lhLJxt539wShpQBd+HQTFPBlG2VFefAuYBtu9HYDJ3L4D6YeY2vy92z7AoY
pB86JwXiy9YmpeEY/stDQEjsFsWK6fqakGMs26G7XhV94ghFSRsMgJuSie9qSRFMltmN7Ab5Xj5n
xVN7kkjRtici290fS89CAiLvg8OwQtgrkVLFhk/nSXm1tyE5GdMtKL1uU1oBI6nrNbVIvBROal4o
eyqCFTGqh1defXuNKkg1Ja3hsKyZ+RmZ9unQHcm43FwLge0Tf2rFj4IDKR4nz1swJnmc+9YzuXS1
zRDb5B7jtUBd2vqEhpnaTzSwydw3Qqo7h6t54Aim5xXb9akPgXJwuszVGKgq30Pf/HLteIWJPy9p
if2ZvRVTeldsOT6I1HVS1OCykqNw9oHPeZAlslARSvw5OG/hXQ9EjXp8cYapJNOH7eGfaFvpo+80
VoJhBU6JK18Y1W/f8wGU42a3UekOZkzVkSBBkaALZfvGQo7r8ztcD3d6olqVLiKIOr/pyeZALPzm
S3fD8mdU5SV5xGLTVi5HBFIeM1ZH++h9N8N8PQb11T9gurwDnS4CoB5NMDv/qKK7uj2TXoVCcg1V
bBpNEU0HtN42DWoTJ0Yg2DprpxoZHi4uuSQ+kIwWQY63pxmQ4qbAbaIBtWusDNs5JKwP9qyi2Tei
kwgtY18ivqY+5eDTUNC5Rk9BrlZ6EDZEPtuvkqhh37DVg1P/lmFfJW/3uusyMl6CONYM2057UOJ+
2+4eWyzqhwzSZe2816hFJrTAIPp/91P+cI02o6jJkNaCKXh+cE6m5KYhj2TN8lBVf2lm458WmUvC
tdWzi6h2EPQdutHe1S1jnAmOOP4l4FcTQOrxz1VIT7bPFF5UmibxPSuYLmiwhyMJNJnuIWfhdUEq
hJ2mzO3MuKTIN9pFnvIHii7FTzDOOHoYBsmODvkuSLifOYoU8wI6a9nb4ZZOEkQ9QJMOScxrjvnq
JqOIm9F49CGmJxcVBpEBPJwEVKjO7LmKq0VGi1+Q7Nofsjq+2/OX8qzyxwY+eOkNt8DwnoY3g0AX
cFRvdoYEvpKm51cGrrbU9aPhoAc88fy4hVotzCI57hct3chFvHOIfQt0fd5NHbom2g1C/mgUDSH6
eoPA3Fd3Wi6YyPe6uaR8wm4r7aCzGMnMf8oSEmMC7NKzLoW+ePiKhDEn5G5CdnG681INzWGtZ1ym
L6E4DwJodgq+FPdbDXwIM55CWVJq7JPThmt31tIS1G0WyVYVUIlkHzv7retN2g5BFaKa3fcrJdUN
Eqeq3MKwlSQBRTEU5rUhYDZgtifLKD2HicuEUR2YP/8VDi8J6YGa4oWURf6ft66ugsR5Xh+B2wJP
SdrMeP187MpgnrX2/qv562hrrNesK/8bmuaEbVT42Wnir8Kr+95W6Fq2ngnA6yEcHz9cRTGIWaEH
7eD3bu8+2sALqSUwW/KD8ctaZU76gbSteMn/woXKHZqJylq0Z7r6vPA0zDCADKNzZOl7TGvB0Gbv
ituOfY25ZZKILN6WMARQUbKtS2pa9fw1onq5ogfLPmtaxf4XCdCzeIVWaP53gPB4LWjMeEDA5hCT
G20vhZErESYfNP4sNn0kzbW8DPZOpW4NfDl9wtNBgjGIEcLdN2iPpTCIITcAGejypffBao2YIleD
Vo1sJoeAIj1iJpSvGFP78MHfBHTJL3X+ErYHkhDZ9/IqnGJExha5eGmUYKp9HA2EYyCWmNo8/vt2
WHlVzeIOJ2h8+fRNbgbBEIS/egq7qVmbyto/WPks4VbB9HGGdiyxPpPxU2njKdpUxLRHoef70hOR
/IHbN5t6Tkvd280qq61thk77LgBNWhwsdgJ94ha+Tnxl/Tar1abPspnZj/YMLrLX2Bv/DMEIBE/l
HTwUPQR7URjYMinva6R1wHMmZwGHYtP4Xk3ioQqqRZW2w2dA0CtTm7i7qiBss8YSzTDmuJKkqiYn
m9+j97hcmWio6v55n1shQswJJImgGbBJQL+RRBldYy058aEB4IeWDtedXQH0d6rIeGgmrVvcMUUw
LgaitR+E2WEfPW9zym2zgJLOT8eh5rHsBKYIe74LPPdrkQoWYJyg23Q1DyD7SaWayZNwH/+xaRmG
A4G4h6Jzc81ZRl0H8Sj16c0NMBz99+DJyLBppwO0pOOdSLnmddva27lgWYT4ZkPGzWOWBO4gU1Sw
tDOhVcH7O9+g+l/QhNvg7sap8YArTl2NLhmin0z74fptwONftiRydzdWMuTbuIP/f9rN4614tLE7
mWxcgvuJWgFiVOMrQwt2wv6qBdACo88vMw0JkzYgNj8gZsUCmuO7buSeiWASJLEKhtli/NSZldfm
3mKbtgPYGRTUC+sxO/uMQVorT4VX0+kpBfBzoQ7C+mFXF9AlQca+5mfKCaIVRGPUL3Da3ij1Ngl2
K0jER8aF7vqY+MvjGQTwGDOo7aAC+WQmuC3kncvfYfG2sCA/FflILqbqizsF98EgbvypUo90aY5A
BJRYqVlW1iWmcvgb5Hj7qp+tnlJmzpfBfyRWqBLahF9wz0nSSX4N2uGGsrZCi48rjrOw5ZGlOgqK
UvgYxKJinF8U3BccP323RdIer6kLZXVmQkSEdGclaqLadOFYicFhMx3j7DjT/SW3q8QYtXiWgdm3
ypxBkX+4YC7WJRpu2It+4xwLD1HvSVWHzQL6rZ3NI3kURrqyzTxSdkLIRPRKK0AfW6/f36GV9abK
rxMXLceYsFgHc9VQBSD+Tb4rPBe1DX9p0VB4cnYzC7ewzCYwRu+Cc00e4nLncUfNUHv7nCHAdybl
FwfA+mCuFO3C/XhnlA145VIBz9EUVYMMz7Ke7wKtwH6ZQ0ZkwNhXTUj347v0U0q5NNOG4Lb6Dy2Y
foIZrNz0fuejs1TVHQ2utuJGXZ6GF9IL/9yCc+pMXqG4geQpW4lI1C0ClsYCIvSI+m7BgHtRqetj
WfnnzaS5kSJwxSFtu3AIO7Tn2hEdKoXZjBRkUY+GgYOP8JpUx+wAYHKOvTz+3X5Dqf3mwsGqqE4q
VKl3L+S+tIzaMlvZFKOFMWhU0WtzsyGJmFlYXcBMdn9dFC0V/DwIsajPg41R4hnEPAxuxsoeEr+j
1iyXkb3PmECFzYSdgMPEAfcEZuvuWb5QcpCp2bWE3Y5PIeF1onRYCkn5tpjyyPD6YGaf2js3Iw68
BZj3fKCudYrTxvlnjK3pCT439m97rIC4JaxumTTcDmrLO7HSDxhDMdUlbntMmRazHQ44ppdrdLo9
iOAbJ/8EdEX/tNoS4y/CmcRNQM/+poOSDF8plUv/IVUR99cWemPgsu3Uo5G4N7Drq7KclgrofmDG
H10YD+rnK3dOPyehKtTWR3DgTWkN2pVTLxNtzLPNz6xmuaAs6km5MrVRxCrzNYqZ9f3mrGya71KM
LmnRNjQia00HKwSfd4JiOr7I8ekXgoDF/ZsL+Fp7IbKivMJ3PyeOYXhVIxQzcdVS1KsHlcLQoeN7
3qRvT/UvgWbhoks1oAfqimXtVxkxJDKHrt+nWeB6sTwLRh6wLIRBno+8i+iNkUg2Eo3sZ/l6T+6q
WhLw0o5JzGqO3H6NB7DufmSqJP5zeU1Tosus7g8Qgq2WLHQfz7sBEbx620BclFkI9JwZ0KYfn22j
WMA7PgeqjsrRdpj7MmJ0Ix1Xu9VKm0K5CXNju+Pmp63z9RpN9hId6JGcvaX44Av9Cq99e1oHhEK+
aW/Mn8Zb4ybN+6i6MpYhSgooFIrea2rcHwPAvdgWj+dBjHnlGaP+IQYEBML780E5/ce9Es51mpMA
6K3OnyT+rNlZ8XQUCMAP57y0YzhS9sT+OR6nt/GQ/ZsiNCr47W7FfWlgjoxUgL4oSqzlaBM585Hm
2Q+8zr0MINyFGyFzpLvYSBThl5R91F/AztibS52U6JKpoNeaO9KDYD5l3ugHqtxYQLqph6tfw9hR
owQud+V6dwb6E13UAUeuCneAw4p66/bn5QKQz4XjGAyjWqABqLUC8YoESsUbsRvHkiLbiR0B42Py
w+whCjI7pekb21fxxUXEQlV53VtbokAnQDh9NnafLOp3GGDkrdnZKsFePZKZQGnx/YGraXqmN/v4
lGEimC+ELQJgp24EBZZUdiGYQPcgeIlO6GR6eAY0tZdppAEmcuzQpGlT+9NJJcd7X0bztei+8AsX
DtHwvNnv1RrSrVOiqSDBw7hF8Fx1VnoaCV+J9tD4pQbDJOILFSn56yAsji9RMogLDdR+JeMbmfXR
hLzP/jvH7aYUtAhiNbZ1X4mbH34PJ/+huwUAWnrsFXvb+OhMkHVP0zW68EEGXc4mRZn5AtzYwn5d
dcacncmsaGIROQZOQleRu8hD1LekaQo4K54Qvzk9ApghLhEXCFrQ6rAPC37sA1saudnC658yq//l
dct+uyOK1KLk8/uWr3PHE7/6pGiRsQiaHjmI97/U3R7pN7gaRlXQhmxwKx9dqBkL4PiznIEDlmgA
Gc33cgGoQEyopcHki3eSHInrGLutQHRFhU4STOEUZMCZnmHqqYnO/PamsjkeRkDYbdvaAMja9SSt
u6HYealx9V0JrUFVaQ7OwcB+HH4Mxi11HOuP1D+l9+oryFgkVArgWiq2aSStDG+pQCmGHGzIrYq5
w5A8jGUWYHsG30PTuIDp9dyvXAAgv2vvBhMrEmE8R3DvxpxS19uJEd1Prcz7k24tyTflBGbbt+rZ
Ij5/smtHblXnvn9dt6KC1/1bbtRD9FtuPaNm307ezB120fUvWptkrSdTICwrw9r8tOf72YXavKV3
hYpapzLOXBa9rezJsy+SDHa+3rmrj2l+scOzivmq9TfFOr3xJCqg5o62xzvDnadeeNVu+DAVIUY6
KbKCUopbjvJXAAsG6Hz7rH8Es02njdBZVr0Ey13l6XofQ0n/eDWoXp3MVgKL7uhG48efui2gBIFD
K3vHJkpuVvUjBDBGrgDgbdExabVRFms8s5bSXf6EiKrTaLZuwtPHmwfKT2zaRhdhnEtA9UVVaWuH
3mMJL73S0joLuUKaLWgKo+7bjKYV0nlECLTPrLDlu4e4hh94N/x221ldSMXNXG2kRaZsL+RucTNk
dRzGm/rUAdS2IwLHFXg/4w9b7tT+Bw5mywZ/Cnnl6TIVcQkSiBy+oxa2BPlx5/DfkdVROm8dUl9v
2hUCsHNIKImhQ57e+Jvxzl7texRKIYjQbVHXuDKt0iUiP+1tH45uVYDv/8dbKZOiZtMRSJ1UYxrJ
T/2Ks9OZD9K3xeSeaSkxil56nZRYSolmtfu6+96ocYeB9ZyWEzaP5TNQD95LHPQCQTOEFIwpOozP
1ZT+AnUXD0EtITPdJd8r9TOiB5LC2ciy1DsraV9uJw7af8xWzuW7oZ9+wzEEyUxlBUJzR14baxGJ
C5lhy3BC4OmqyWsTApvI7ljRMaWJdCFQy8++oztG9Ve1WMkW2vi0ulVX1bIyqKjE4hRy2gB14M0A
vj4wrdgnqeBe4TXTv06YkivBMvny7mc+GHobFIWnqwaT+Ff74Oi9NuOOXrz35tCDH3CHJ2tAqNiO
r0Pla2GuuiLlnQbJwO0nM2iL6eYamTe1y/bMOShs9dCjzfcZHLc4lTtQd9nBtKI6xXwPdwgBJNwQ
GiX4c0/YXbKrUk283BglZ/D3ymNIfTXKS0jgLlcDpOZEDP8NhpiCEiPBIspSBDvuK2OJ3iaEkZFM
q19vACZnksftOzJB27KkL+ny5yg1insrT5C9ZOLtTdY97ecg6gO7dPBHLlJMijUyAz6A+m5NYePv
4Ior/MffGEHn7P1l362v+vFHIMr/ijEj0Q+lxPgj/xyYBv1AxsEuqhGqMm+WeQgwdQYvMx46gdDT
AY1alcxn+XgjsrkXXZYoKFvI1GtyJCYlDpudeH9ESedOBir+kW40gO/hYsneDYfu14yXC8/RWq4i
7OcYv4VeZmoib5W+mTKDn/97MUCATzKP+cLKUTNu/uPl0wXzJMb2MhoLHBnha0IatlOc8BxOpEpj
17iO45Gz1Ia9bTaKkTNfKd+qnRnbmsHH+d3ot2qLYRAKByYgzyML8bMmJI2R2XXRclxGbRy6OmH9
7/+pXZe8RofdQKumfGU5Da9M+vMxP0NjcwM3AUnIFG6pieMDlAh26WYbc7SdWpdaYera/RqkxZji
ADuMIRzRq0cR+SI5ghjpT9TM83iLFw69286stHK1ZS209Zs/sGz8ZmtM9XDzHZoG4xLYmf8ojSbZ
IqGEjkic+C7ABhyVyh1cv2AsZxTat2pXjSwTyd8Gw7sg1iajSZugcgklHsOj+m6y+whrOjVOu5jo
g2lKQ0GFKgxCl+aAP8C8tBz6NzM0HGhZ+tCtaATZTPj5Vt9rLz71zgGcLknEtfQ2nlntTbBZxluM
p43B0eXPH3jKB264vqRfsV3/scefrmO8q86EMJJ8vYp/2ED+TCsOQmcHvrKDYglrbLctBhN97HXa
fu8bnNcSoJNNKRwC6ND8LBT1W1GRg3JEqaPoBlTLwFkueCUzb0oHkZiGj4nl6BscKvU2ExdZxQ7a
9DcK/Jz1XODcntFTzFgVaPFARsDSgGM8Xt4Ux7rVfbQfaD6lNK9yMgwrpJuDtjZEfUB/l5l32a9j
IdyYNiCMeRI9IyMDFUneSZ3NAZphd3emL1HP10u4nRH3t+VOR+yHGpb7VcrZ3XrsnuqdsOtRlLrN
bpv1lYgW3Qj7zq0PANIbqKh7P0uHsR4PJxJ9bioJ/ekYyuqHT+EWPQVsZ8jYdO1gVLvHopyPwQsj
p69XdeIaAgKfqcdqk33ASyf8bdxXNcHXPZkXAZSfSn1wLAMVxn4obhmodX7wkJifT4rBLYNWH/8h
roc2jc7QAt259Yi9oKIvu64Xp2PdGSBnHLKJ8/D/kr5WoH9y5H8ow+rhwXk+Mo/RjxUbXs/8qum8
E0mYhgxS9XCRrhWwrl1slzyz1ror7Hj9bLGswDi7D29SOdNViAcGUof1XpkPG4syFrJpT47/u59U
ONmMlS1WPEJKeUVeY8KaZZOk/71r8CDzZWi7EB4EnYX7bQeGvSYLwHiGQnRLJiRJNaMz6hzJsxqJ
pdlGxshMo14QL8UH2SmY2wjkqH83dZXsdJGryFJJTk5kl4FvH6o7rCIT0kEN0jAUVsTLjBt4wxXF
q9Ol0J1KFgEG5ho2ze5W1bmuko850go9Bt6j2ZURXLzNAae3YxQ8eR7Jc4mXCYo6PsntMW1Etmwf
RW63N20OB8yDwla7LZ6yRS3b7tdNgxTJhmYWKvXf3fDO+cJPDEcjOBq4LFt2KbHZGjJ8R3EYqiat
1VxLgPj++SeEvRagZrd52a/qiOc4KtiuqlfhQJHn25cRNhecj3yIwa5H9nEXKWi0K8t1W07vyJiP
gO/g60hL9ZF6y0ar6oOby/b6z3cONCibdTg947x5Tj0zMXuKf653U+TV//k/TuKuNkeWq64zJ4O1
pCTDonHH9O4OibX6fTYU2O76SVJ6mZ4MItAjqM4DlN1wrDAoNoKxz9gekZ/hD1eUrsqms9852TQ6
rK6FiAyznqfNc7z+sXrFUREMktWJ3/zwnSzxfOq5JIEvNogSGW4zXSsxGdd8E60tRJBalXmGyy9T
e7LP/LSm+L1XDWaCKIasIKJPmRh+jA7pG7bmZVaOR/MpwO6OUSiOQiaqiUtsOe3/dJhhOaQv8VoJ
Hyz2No7Cxnichxz1Mrfdd3EoCrAuLNyoFjXKnklGOaJWXlA5GzyaeoJpZX9T9LbGV3GGnQMQGo1C
lhbb6wMqFfo8RzMy2jDRsW4NyvWpLPRhkHaSIx8Vs+GrhpjGqR6jYsEB0nSgfGAOE92+IGlNfzUC
wmaRHoSX2MTVFGG59nC4sc7RpVdVDcTVc4KP9pM6GwbH6fMN++K/Eqi+/F4brRrDEuPTzwAKW1AJ
LIuy3ywpao2FnC2mZ5BDvknEES5ot3+lmnvShSbSaR2j6CqHQ2OzZCuAZqO+/2Q/Nq2d5VY1UgTZ
E2Obffx8Zp6gtEnHnQodvnQHHVq4pO1vjA5AbzNQjuqOvCvx+j+6zDz1yuH72N82F2WRsT9yWRzg
GOEM484S6IVkD0F6ZPohhZeaQgAI5eDulZrcyttOXOyqESXqoHYZpaOeh8Fg7plEq6jE6uKppN7M
vxpGcgkljl205AVKMZOJxSyyQgxN1nrYFjxXgwVxYn9dVEEfT5wS+PIM+5E038lwOqOLto4cZyZ3
+oIDcOVfvYTivjoc1OTrBxn2HQxqiool2CeItFiKlAJ3qkMfgwC5RRFwl/2yjYM8ArMAfFewBpC7
h+g584nZ9rR9UwODrOi4iQERZr+JIsCdwerlR4aeoi2o8utnsLHKdyrWfykp3JKVZPQX79IKArdz
A68f6vbcPpIS/8niTpzbVkZdwmbo9u8RBHTvd/icHIBW6t50Yg2DkkqG1ELrFVmbNPcls6EXjK9k
dA0CNA+/MXHIJxxndWAGSHKFhg8j9eDFTpcRrc+FaOO5s9/IOuU0bG3OIXupqo84neGHmcb42B5S
KjGFt77FN3/R7I2HcHYF5LZH3XY2bBCHHiu2afjQolrdUtWXuMfSyKC96QNUDhhQgBgvoPw0yYPf
+zYFpW23NbLtYFJzFlVI33mckdkT6dGzIC/dXHaIepuXPdORV+3fFcZwwllCUWSe/9HY76ouXiYm
/VSZXPZdSTeGU/asUMvDa4lfd6VWMR0VVKT2udpTLv5N15UMcr4Zo/1IFWzyTYZ0urxPXAEt5ZON
h3mjnN5NZbpMwQtZaFcxZ+RY2hZVoQY51wWQnmFtNp2ff8jIaUMkjZnsrPVHrBcCZh7p/cw5yAiX
uyqEjhKIEQwjN+S+KklvKtLFaYvVl+IaFICVCWWAYnfI8G+IVchJcexABHLjBHUGxxuoDlfKjQNK
WhBbUY/RV32OkYFRux0JTGVCTLOmzRpu/4RkmJ2JOv0+P3q47RBf7Jg2DE4+RlJpfxf4DoGAznHY
BoZnOddT3jXyAQBi6zKLJi9VebGeaXX6ZBG8H9YI9y4PJrmNR74rwi8duF485O8U61pi8pELXUj1
YnTQvKekNyfrNIyYp8FjgrOwfKKpBPOJ5E5l2PZtOp8mi0pc4VqIiFT9xRNATedztW8obX9/yJVR
62WHTGaRFnSgtf8FFTl4EmulpKgWk+kxDMFyO6ph4vB0DNbyhlWQjNRf7qJOoO9ygvYUFB5ateCu
5wRaGP+iO7qrGiw2Nkh77F9xkYQY1yHd+qTqajitlKaCNz3suMF6MxBA7KUlm+srpY4MlStMPE8f
FHrKHXdKioKmMqNlmizmmlMnUMM4l46wGCWGOWSxhgdYpprNNZjqLKpV/lo8Ky1z2i4ZXWAK0qez
XjzQtOZ0324wU1ggQP4/vLB5inZ/2LdEuW3LhW0JqH7Ivxi55Jx+6bFJGd1Z0qQegBxarNlphUe+
fv865Wri/ju9pGBs5P5J7P7T6OufkibpBvFJv3cqcW5jWJVGLyky5+YqOXdgEWWO6JudeJ6aOMDA
u3TJaM4efZzThTOxcDKMvrpL8ANyeDB7p9gjCqK/74AHi8GFIVa5XWovjSxD6N67zs+16CGbvo0a
xs2yQRxzGqAke3yUoacNhJSb1yBe+hVpl2QWCum4mAh3P5dHKNueOcqqEx4dmcMbbmLk8F0lLtMj
GmaFG+WzfHJXt3Nb5J3HsXYp6a7GYs21cH24bWoRdDMg7aHuMpav7jPoK8jSe2xerEWRJKYijga4
Aa2Rhfu0zkhe/ccAEWTa9TrelZgR5akITEFozSymSf7YEvlru15ZSSVzSrDeMUfRSxSLyOMACGCB
VOihdOmVHYFsTnzXgb8/E8a/6L92Q4y+6u5jq7WBNaEecQVkBvGDQv5R6M9CHc2Jt3fm4E0n5eC+
WSCSmRHnj89h3RbvTQN3mfvvORY1G1GVbRC6/JdBe4RDwNU0oZF4ho10O6eWg7wUy2QxYpjH6zQP
Ao4yiEZuD7Ik4KVCLgx02ew8uSkosAkFre5UlZL/wEWhiRIML2tk83EMr1JXGK6DmydDK9dQBI/a
mgnqJvDujhVIwbPi2xvxFcuIsrDvFKojiMt4+992DdaERv+i7KxDlrQ9flLmmGq6TmNJaV4494+6
LSrkXmfDc6z4OHsPcb2+7+GPCQLJO0+Fs4BXKdqm8qGxPYKDXPUxVIMbxCoDBXUoUItKTrkaqQ4y
pvnft9NV2Gr+n3Cen628bcWHbeaG7bAbFxUyeHK+0q0E9r7z4VQywyCeqQfltc9MIsmWdt81YhcW
5OoC8WTUpPXfk8XTqEhUPkBDPLbPQFETiZV4FEKwD2lD+NQGR9bnPLgCuJfeliBAxWKZy1+1Eh/y
cbOMG3OUn7DX8HTR+1TtUbEfKvToAeNe8nzSXKmJgsjp+WtXKUhJfiVxikLQrK+mO8Bmbno60cYK
TM2CgKGqJBnZO0xzdWiks2ruJOXGLGlFKRVdtTByu9i1WiT/kNH+G5Cqw9srb1eCtH/wjWec6+8n
LWhFMyi6bDDjmTY3MUEYakjCny3UZHE46+/lylHl/X+vZLPZM1UNoIijeseY06FbipXng3Fn/5Sz
w8E17pDs/EEBo8fNrN/uebo2gKdBSIFSufTc4xmGHpmErwQrufR5Rn8uZAUn9oeO0NYscYOX26FO
uR7eqda948xlpRymPxtMtimC1B5SK+wb4vHICR1S5v1/p9iekJaefKIzQ+kpq2/yljIF/2FTrWDn
S7Lk8L0e7momq0Oh4+1On+HwzbdEfDXP1NwhA3gSId+/xOzeEKdY43LfJv2PLfxHhjCziMNHk1xo
/C5TSOkLRF9kJIfNmFEu9IYFbqUUKQFpbrk99dQgb9H2SfQkJ0pJC2Cddq7oOaUxre9OlOJqN5gw
gTtLCerXfuJTHjh/4nqIEKXMUcJaDARd3dESSRDausPVmPydhE3u2pRcYWFlNxR7gimZSjbHDesb
A7G73/VS1gDUZY0Es2u7r7fc5reGTbPdvrgMkpQVtb28NxQm+79EHx3NMg7sjLbaev2aSBwlpnT9
b0MuMLqh2KtIksRmClJ1MfzsSdDY4SIS+SbrFtYAJw2mFm1bPoo5CwM9lg/3pLilGo1XdcUTo5y9
m3fT5wRzdAoYuB6fvdvuGs4ePp2+oQuD+LM/5iLD/Lu5Tmg1v3Pr78avjqeeGTLN3Y3MVK5jhVzq
NImwJRPKeh0Z9medCkVrCTA+mjI4BzuIwrMkCCjdbZNAB4UxtnykOIa9kwWOPg8Uoo8X29021UbW
QwjWh9yRlvQ+dXMuFLY7CicJYWmITdZQVxnPNzIARDGhpR0xM4Mwhg4Slh+lfdccFWCDqBcg1P3M
WF9THKDG3nxbRYXdWOrCJezzi+1gGPL7zb4XZA7KSt/iZcoivptjoi/7101ol20Ttb2MBj1sLCmu
rY6RTHX7PdZQlshh+lSMgiTEmRDcYIjGMZlyfmznZDABrlrglrk8rJ03oZwNM/hHi2XY+/ZhbYrx
nm5vX0t+skM1nnlXDWp7c3Eh38LDQKhvh99ntJ7C7OY2YMnNjOkgZCAxyu/Di/ziHklGb1mgUBbw
mbWHvzoWwAWpW/C5cft+n3A/5CmqbP7dlDAIqbH3sQ4mUSu4yhLIhb4kxmX70MHf+EBBvakKPPpQ
gqcoJHt3cKyfGkgqqbAVXmQxpE9KJVxy823I8SinZu63y6mzURHpBeQ3vVzFx9W+fF4K+Uv52DnF
h+ooes7hhtuhZVwbLjyMFNd2nRoeYAzmgRK/lW/0rwVXbT1+sLCqWbGT3F337OUDfsHsqywuYas9
YRaIB0hCPKCbAlPCtQVjISHtyjACvC8TRwQgAQdzvWyPp52pUKffC6TxJHCTXGDkXBzcrCiaJAKy
Dw9Gh9rwjrnfzOq4ZLOX6RO40Nmbp0kqf37+1W9xC0c2Yfz2sJjjZ3+phwebM0FAifQRRcX+we65
TJZj5MMajm0xSYQVb/y05tcaRLDYZ19Ix9E/BsF43ILqSZT4VLUH0Vu/xPhJXvj5Bq7SmJ7l1278
RmGP1XxNsoK5WfrvzUxQv6QSzDWHmHXevOQguosWvxAjn6JBPD/fJ+OwKVECWD0gWMjFB6W/Lejy
7HohlJNilpwL0w6bjujtWeAQ8lXqeTyteZEQtYLgpJQi7lBNWpHpfjivAa1EjJFhxqlaqUprQdHL
t6NXxvg/yEnlK5OVP04FoulSIT0rdAEG6H16cczIzBy7WwXit8P+fLyl63Jigh4/4L5S2HhMYhwg
Kwp10jWZ2GcBNzijoc+o8yitM+Yu0Jf49c+fkd1ksIjcuaGTIbrhyBL0kmufqcQ95lvGo+Yd8SdP
Kod+NB2swsFaBUPBWCv9FG2JHd/UWBC0MyegjmOQKtfn4Pby9lXUdF4WdzhGwnvnvKlIj28MsA5s
3ev2ywGwl6pvN7NEuGANYG1AhOphbZu8ed0pGhB0wKmdmBAYNXihnMlYFskjtAEQoYUkL87Me46h
PTu0PxVrC+gVLCs6shGG/ambrcqXLqFjQFzLQWuCCDlG5mpNEzg4g+/9iLcoYkal/JTLu8Y2UUfP
p7o7tTV8anWs/JU+cZrCNnB+SzAbuf9XIk80vBd5oMAfMecs6/stLMvQBj6qGRgwUyRQk+qIgZ0i
GugPCXiVMAAD/bS+aoqV+oUOY8FL1Wu6MqdKnc5yK6bvGP8Evz6j9S4Y0kqClN7Iuvlhv+tCzPEr
iXB5sHlxsmZ5CXi1iUAp0cvK/att08o+jiOX2JJaSGcYte1ivBxgz9U3fwbaYMBsaxSEmXBlDAMG
/o0YD0ro8rTPKGtqQif8GUVagZQeZKdsBhhVyjQ0IE2Tef/OqNntbdy3olQL2bdFgjZ3YziHxGOE
E5FeHGOuV2ituhAelRH0eWbdjwxtTb6pfV57kPUzqBGFReujdCIQyyOUaZQfK1/pygP0uCIfJDJk
HrcsKk39btE9h8CI2Y5j6K6PqVGV041lb0rT3iD3wiLEtRMsEBM9pyACkTFnDTOvMepp1xvz5joP
dq3VnywRDobLvhGEex5wwDesUTCrfh2AZbAKzK450Zvs7LZ4grHD48dFk6P4cGqtAqaexTzjLz0C
EkweABjTgEXm4b8yP+mP0DdHHWsm0G1Qfa+GHPESsHXNeuAW0GE1/2IXX0AXfgwCcRIo/ron5OJ8
jcTa1QigRazgYiEKIuMRn2uUobYoR9Y1Lp60HJfJwBtm7fyi6WQdMaJY8OJ+5N+N+G/VsZtZYteB
Kq4BvOFDDYRtMluXEgtocF375UTKKFvlrOQ2gyD7y5/bjiLeiX7w7utaFF2BJZfkjBiTvzCkgZ4f
vBGtgAV3jbfM2hcL80fH4qeOmms0Q12UR3h4Ic1ZGneIudlwNmqbsNNuGN7Ayl3bhOwMdyUgqqYJ
Z/6ODZXoDC9ROOlU7sWR6Hq9Ivt4Y0b1cHmjJt3WAWOA/wdjvlk65J1g4nd3MJD7dbnWaH0ntRQ3
HMM3Ve5K+sCHnUNa60efEJb0ZGVE5Ve5VDolIcpJQuGXdQ1tveL39cplNfx3koncnNab0U/MiIsd
Oqeyi4EeFw1+z+fJM9TxR1hDPwN08+ePoHl4KowuDIGXynqC8MP9LhM4se2EJHClaqoOdbstZfmJ
9JEenY47+MfVmQGrQvjFmGoFYWcli9RjPzodrQGeC8PT9JQFiloeJwYZAGC/AWuwyIxXGNZH1pyg
yEzqXMPOohCN08zjKajS1XK6vhbUibJ8PTulBaYw0t1onNjVAscb0SZYAJuNCEVp/Uc5nPt/WxPg
WotH71Th0scCs45tG5XT+7w6vpcOqJUuVAGdAVMmP5WxsMpSHCJfuYngmtkYAZtarwrmj5GvR2sF
MskQQw+m/JIjRF4j5cm3103rsMfmapzyg0X0bygNzUnXNKhKKASozFHyZVbyajvrvEy2KhMoH/S2
cMz/we5EpJbZKQB3W8zZpYMH0Ev66AKsX7yd5g8WoO6j/qHQA22lKZulC4gDT4snE3HnTc4Y/U9t
py9yOyg8GoCZXhINhAXnJ0XYPnXi9V+QUQzHzHtcqBrGJM3WLQUnR2A5nQ3qzw25Udim44PBmZ7O
bdYlPj/fCuFbE/RBKMxuX/WqaBCmDel84pbE25tQ96GChxy+djtfVj8t/SjKB10l22Y34vg7m/3L
zohSHmj9a2Bbw6TXQWKu+AJ2IsXTefDWB2gF7ThBYrZwZiU4uhVBmYvny2C81O7T8gruQ1V13N+K
iEpOfv38W/hC8RsVV0Z3rGE+dEYCjDLq8v+yEoxoMkQS8WRZ0uX730a+vnOKUYMOdKaB9uTkbrjS
aiXtMMaYguA03da+rvZcLlq718IzeHtiHbY0liSTBPaygC6rICCpPyA5CB0AbUuYAiQGwoYbh7MB
yXDXbm2ZmXwXRLBmZjWCHDxfYoEuHsip2HSbMfGfignutT37i2c7HxRygLKlbHjcLPIsWNgOyi5c
pGflBmV+vdEYhQyXsjS1yeNO/8xnWCl8bnUt2aa2s72Tf+b7DwtZYanGtZazvD4Ff8DTi4DECqpz
PH0i0OWJ2NvafZ2Dk3/p9wduy5MMopXnxa0imYWLpcLm3Vv9eDfGi8meaidrcUjC/+hywBIwPYsi
LJzkIWmWQmh5SMLP6Af/YO3az94F1lDUDSOt38djhiy741+WGLyH1TVSYsUwWMCxbG6houZXl32d
bVaQVAnK/m4q9pVY0sC/Ym1qT7uZ8546MRlwYI166VV2BqcrbGzOkT4WF/fm9Rp7v2uBqSIdk5TR
1YcxIaQIGEAA7Q5wuYX0K7xergMnUoFBF7BVdNA1thDfn5Q9FqZqjFgasiUYEZmopA/ncVDl3vRf
RPQC4gqcJ/syU3hJS1FMVlfGue4oQK+febTC1bE2oT4ZaDyb8/JX1Yhrf/o6V3Pf7U3s8vAtP+sx
1/DMNwqGmFyoSK5iBicaz0cVG7HjnS/D9VWtse5d49Yp9SkOXosTsjyd+6kBdM4RXwDI4BqRHvrD
aJ83g/GNmDCBs4rkOL22uMEhfnYEQyXoGqFAMJq9/qapLEIe/h1iW4SjGGOxksAqCLie5zuQy4gl
UkEuNsSaKBuVauGrmbkfe7XK0+8rByp7QBzE934chHHbETHWNmTxGmwIUXoRwOM4uY7NvZnFmw3J
mcJc/IdJzxu06myW+PKZWEQJrYU4XKEX37Ogao0GQskE7IVEBZTiRdZkObHGakJsxj7p+Xj8aYXy
dMSg/5lXFtCXyXfXT3PH7HrhprqE0YhvqwWhJ7ArTgjVmDibD6TedyprtjMPwz2eV8GmSJXlKQTU
rqFNtdFryS+AKl93VleZsrMjdRvmdWgB4XWxjvWppjae+ie3tNBh6WzsMf6kPgJA0xzcgGTl0XeJ
05lgdDVx3QcAcvrj6397P0QRwS7SM3cuFqemZ/sfDF1tkGr6cIONyQFfTp78X7jWUYqwwryO5oDj
0BD7/6pOR0bN631ATe4ovc/+Yi2/l3evpywkDGNvHl/1BQz3C9vkwcflsOI9QQW3aGZSB9fQeY+g
r2YEEI+M9gSDc/cfHHZ+hYxcwT5MbiLRQkP5V/CHbVxDOAOy296KnhFVg61xPiK3l0JTOl0aoRtu
z7qdBC6wh7X/pIlUYZJhvYY9Tkub5kZFcHllxMntiifF4WGs3kkpPzALSDSOJmxUGBeH5vhLCLw+
MN1toAzSFvF7S235qOzkRe24+VufmRBFpGlcYNLh3ssiZya8GgxlSBeb+T41W8M09kdnv0csMizo
ZqfKzjJ5a/jfLe6emBaACw6TevOLu5ALr99JgkCRU6UtZakc8OwLh93O+Z6JE03AAyU2/eSB65PA
b5tB1lWdsEBAWNmHoGu2GJ550UhvLDAii3jriZZEal7bOzrcP4Pp0Lh3TSRzjw/Td6K2WqVinkN2
sqwZaLaz9noKhIRn5p6a7i6HWqIpwW9R5cm1RRHEws7FBYqSNsnSNE8JCaCQdqfaDe79vQXVLknU
uNuCtgu7EWnlU9emlJJZMEjaq1tTbf90pVseEpW5cbCGh4QMwAHMpcpomFRvT8OppAL/3RgwfvJ1
rrKrZ/mMFKdaClfS9opA53R8xVwJmodi7nYUloH6drnWLcLwqtqtHLj2pirLB+011qyqUHhiKCsO
bS3nFaT4dr1m4pGbT4i497LULLTHnK7vfOqDUskCdvS3XgL7f0hgJG7dSCY4AjSe5Goi80MSQ0gh
FE0zLvXAvh+q0bZzHzNkVs6N5piiP1UFW+AyJDkQLptrTQtK7fL8ERWQe9AxHlMh5OPfphaGk7Go
MTPQnaRCFtaA5wEfr+W192diSFMAmfdMXy7BbzSgyFjqWkoNU2nz4NwE4QRM1outq30kjYxukM+o
ZntzYQ9LpFDcrVQcIqOYRuknc3kEuZan9qB4dKGXwhO9nkTTjTO/l3zT13KooM9X+iDWMxhDpDN1
CyBM5/iBRKV2sotom7FVVZejdUb0KPSu3wBj0jaO6Cjo0M29ukGXO8+AS1QZ4rlq4JN4KqQ6VCpE
/aQzsVgCCYF+UqU10mnktLf80eMwIhUNp5U7tXU7ED+WJrBGJ37Ob/C4g9imkgv9dp63+TPJUOdX
MIaX196E7AJrejTKVIpmD6mI/09qatdD+QQTOxrmJqeTpPEVrPa4nrfR68eo1569JV+4JolKREmD
fPbUI0fQ/Z9aJKdiqsDfqlNKvsQGKPHzYoBxZNW24BfHn3ES81avrecGgU0DcbDkP3EclgDKlpiA
w2OdvErlzKAC9sujloDbPkjNAKF+S8cIB/gfRCduX9mny+crg3xxAkZ/5yAWV0+i/EsOVveZDBuZ
kte08rmnUD6RnZydwv4v0rQURBMDOyPcYvYUqzP2KUOf7DKlVJafZ4QCbXcVFyCv2eHXbPnWESST
4mVcsZmvhGF9K6J0+CQfGkcMz3U8IIQdHpbxlAS6spK7yphHt98uwCJWjfWt2WoDY40KPBaHNB7E
O6OvHK/K+/8URTZiV5bxsp3u+HPWx/8VAFCzI4Hv1HiagPWgMz4Nn8Mn/woRl6ST1W72SCo27tNR
QRvjuB5Ll/J3x3IZgTDR5g3kFEc2xGXTGylGoYX+PErVYEe1U0ngN8go3AOMLrAGdayqL/snEPOy
5APPH2sXWMyKRhGS9mDe3xm956bpaXi6upm+NZpHHRIyVy4duwmdn6Spm9VFHqa5QWIPIN9qwiWT
BlEoJTVbgE0ZxlEN/Lu4WARtvpMMaRNNGCyTc4aI5lwBlpWTvcNknhJpo7Fwf1GXQ2Y/Ipc+GMCS
K9FEBRWaAFYeFQtdGtlNwgBRSGifsqwXlsGWkzhVSRS/YaNnO09k38e7hmWIy5k96Ko4A2lJo7rG
kjVoA67qZ3kg2z6DW19rii+vPbaWD6bZJ34+WbJ+uwq9c+9Nso2s6oJgsZvdT3emq7XDQw8xXcRq
nrw4OT8awxEkc5RuCsrFYhcw1Wfum3+FuzJXJXUsZQmjG+rn0k2s61lyiA60SUfWsBnxs3hXYHxO
/zGinxNeIRKp86ldyRp4KrID+2KxBzhecsDfxzosihUzsEFKAgeoqCBZb85Hug7Bwec6D8TSopzE
/zY2Eyns9WMSU0UsRKg7Q91u79DSLqNfvDeNchihlRuqlPX261B1c1r2gY+7N0cGlIWzJuaSRF6Z
9Jf1P0HCxsr5CeOf0DD4bSv9AsdjcxmLx/4cZSt5FnwiTJnKdl+ZmKfVNONkIeEfkVf1EcGqmzOe
AEQT73SKuQqfsQVQNQk1PqhUQlfXUTiSxQkvJ+fef+UzdSQtGsHmb9wOdhiI2yxci2tOKi+Lu33F
M3SOUmYGhbJi53df1a83Y/dUKUzCVZQpGsr30jTbV/IJyWQV+RMijj+KGBAdMHtYsYfHJVz1XGY5
qTjm9b+NDqWSXevjZXjM+WkaQ4mUaGUJilaclz5N9Oa2zUMapo43DQS2XKTqfbLYsmJgdh4zPIGl
eS8EDQ3wpwVU2eo/VloYC1BeNfOel2ai/jsxoU8Sc1g9dgcJ+oXnGN5QypKnbP1VAdSh78Wvqly/
FnIXCeOWGHKBTJmO/u5QU7RgLf5+SbLWbGmspwbcJZ7E1ZF7te14a9omffDelFpiVxZ6Khkbczic
co7y+aK2zw/0jHuWkWKRo3UMlIxWTRSeBuL0Zp2IGGxf5/k/hdOH5RJwdNDKgk4BN8wUh6+Cc4YE
9+1camEbOIzdlyDsJihsURDUCF8bfLEFZJdCCpmRnBIeT4lohIjOSRmY6tYDI+mL02k/Sfy033tp
iUPVHfcrtDfEbkZxLXS0tOtGR6kSqyiXGgYEIBi/B2xnnWmtJ19h2XV65BRvJDJ9kdIv5HB4vEao
ks2IET4lYUNMpfF5IgQFSz1DBRBopi+49j8faxNKW9Np2YVhAAcJKJtYfHLmiYvEqEaA1glZ2t1H
cf+cTiJvX21ynRef401/HaBtGLBcVGiSw/nnQJ/HsAUCgKlYICzLx4MeresXAwdTXVAHGrP2QC/K
lrlOO1fobDrbjWkp8qSYw7tyY1e1D9TelAQ6fc2Zlhc/hzaNbTFpFAu51mwCeYvyD2mr+fujvk7O
doINindYf9yu2jmlT04jgDJrzVPJolZz6IMJ+ad2IBHx5/f21JwF5rBmS2rShdONAEO0P2+2nOqw
AeU7tgN6rjTOuzsifnx96FDFeS+792TzcKFwedgQJzgkoJzoLlYKLyGV3+9tHY2w86QxFsILOdE9
zuuv8S30cOMXvw9oCGLJNu4q7pu8jCEnHOA5cpQOzn14XI3HKB+Sm1bL6iDNwBV2q/CQAeQZBzcb
srbftMM3vtgk+R5/+6NvSnd32Q8lFsQECdr6yzjNH7B65XBtBsb0GM+/cM9d8i5+YMWcxtpYwjub
U2Xc5FUTLtswiroHHluRqgZL8+m6etsdAqC6OPzpZKqSeRXsHEFdXkm61/SuDeFHvQyE5RO/HCF1
ubys17kDv+YXueIuCK2mCmUM9q2RGLXc1ynk6JP1mfyt4rzDsaYx9NA3wCUalmqYBpYw7XMgs9B8
sAoOQUefUbZkzNEbAjlSSoBiIDJQB34VTigCURELeXD1RyLQLmGe3aqSf9N2SPU2ajNxA6NCK+NF
IFC/edRvLbfssq7teH3QyaTGDHna9ZIJm9X877TpS8kjSo4/ClGyviPQDmF4B6x3I1B+TKTagExo
QKOXHa8497cK2Ex8aSwVduJxQCJ0HkVETTOFR2x+Wcw7joF/m5a0LatJQK5kzYYWYttQO8aODiHD
0kgQxfPavdJXDU+mE/xYLx+vurfNYVFO3vC7rRUTQQ3yBvPB83+VweJP5ihwKRSb/4TSA4qlN9m9
idg8CcN2rlkhNrlYpeZnxMG4WrzBLtQFHZukRabaGC6QC7MVeNTom2nrbY3B7+0YeRBp/qlhqWm8
H6TqeETiSXyTtGjyOZND7j90yOzelbGWXaDq4A1cK2/B9d+saNOw3EKzfMLuilQWAQMoXDLQryyG
WgCF0s2jOzJihv9S+3VgpwLpkg7ahxgHI64FTtR5vihzNqpvmZbf8JgxmczYObEUdNnFI9yghxfB
gE/U6JEOADhPP1Ed3oUdkuR4sSBGNVbPpNwkz49jPlrQbNpNFewpx3NmIP146XpM5iSIEKdiL1oZ
A3KXAVMn6kDvioQe55lUeG/xnc2TJaad8ihyxJrq/n8UA+u+eln/Kai2xNvDIqugnDQqaU2tPI9f
i1NqApk19K1crxq8UQlpmQHsjF89C0IypmmmlVY888XgwL3ACOg/V5hghJMw48NcEA2/6sCy+N0t
smiNtuX4cEjTEC088reNR7cOjThElN7AL4ENa9+KiWe8Zpg8MudJFQfGGsRpz2dW9Zi48GDII55L
PceY023ZCmnkF2wS4lcFfKCoNNIZz8vGVgdhYQyJnL+lxeXl9+q0GRQRbZUdA1u8HjT2tIwkY/Jw
cdqE29SB1KEV+PdpUbHzfz/MDg4+74dMd7kxjyGxZL55ZfwNobW86abvuVvM/gjt9OrH5GrAzWT4
lfsWXtn+MSomLNzQQMa54pzZjJuncqF4Bw5maEPzhNToWQ+z2ELQYDNxx/BuSneoLK218mKpYclW
fT4OgE2z4bKLND57Pqb73to8JV9ZHQPskBruKlppNU8JMJIPYG0NGdHG+uHonhphP9hkA56LYCo7
KuFTzFx+CT25u8XK+18TMuvwTh/I5Awcg/Isfk2T4ryHl+ltRkl8V+plChtKvF1YHIgbiIO0YJKl
1kWn2M8OMWBTi4fTSNprR/CV8rDgaffL1Mb6i12VU4iRcS9Fmd7axC+kk+II6ghqHSoqCd0bftgc
iY3E2PkbTCqB2XaYOGxEQKODFJu5fDAIflZnrz7ylCK1wbCjnzfZ15B7ib+FxKVOWKIfH70WWh53
EUAgABe2nxMl0kzpKkOatGMPpCFh35O0Dqh2+qLw4+crDtAMyfqlnt1iFSLeXuETDaHFzJtI2bWZ
UpwOIUBwj9Wm9Laoa2rdgtSh6oJxp1WQX4U4I6qoVUzu6fjHw1G2ADd4Mn8Snqa5+GF0FSxjtB7L
YuPihqEF4ltdzRL0hVtZrHgQ0HMsUpxCKYIp/DuRtYaaHOBZiyIU1KST4nBpH60NmaAQJn99zbVv
ePitAjHOQk7bPFS7X5HkJEcbKgGgq+OdNxhIdY9a4IwSJT3PJsZ7dCvhmunr8cUzQL/4nlLQ8bZZ
ITsfMFRFqw0Nd9agrBkN5Z+oEiTpwgCA0wwP0NkqRR+XVzDUN0dS7wfX7hi5sx4S7wJGOopS1V+o
aAcapC2llTDst09ijS6k9ceQrjDpanTXWYYja42OJPQVMegjHRx+6p7hNsIchIxDU88fHtJz+esS
a+TJ89X8YFQQG6GvS6WhwpkIjJDbsoBM26ui69xtpwDSVnxhb/ovoq4Trtn38ozzc8Yt2SllRgA4
r40Qxu109yx8moaWc7MtmKfn0CowE+RnjnFjlQKMBU1wlKtaQaabo8cWYetqHETw4ygeJPqVBMGO
wEBCHyR7bvrGvH0VbQJBm6BeTQw2NWfiDwcDKODKZUmXTPB6su9bD47Mji+/0qtO0JBq/kZJxfeP
DzeVVb18QqwqB9CSEtN/UvOMjzj5UTQqTN7cRkSbOt1905Jt0fFIhbd7emDVooVpah7MlQXK/RZS
fZwV4AQI5TDRfBo+jURSFWHJaLm2ilvDFXFCxrexVzf/Is8mjnoDSBF+vO8uApYkJsqd+z8KJjnV
mXM64sdY4N2JknI8yHjdhTY+UikwIdz35KCZEGlyjZQhTcgDo+gmvNgecXkAUx4nQuixEwpxaouM
7EAEO5ebJij4lMD9C9ZlpHVXph8Sho4JArmkFGo9oEO5RCaSz3RrHW16WhCNe77Q03d7fEUMySJ2
8EU17PB/z84hwKGKt69Q/dKJG1XIXUEEm2AauExQr+oLZq1lUfk0sLbP4+m41lK1OBk8Er0Ef+dG
NMChaUKiLvfIoGwBcJNMxhHAmqYrF00hhaqx1M3JXJrWvkZTPAaJLeTxWYT2wpyPT3LONFW4V6Du
7sf/frjLtwxsFI35BYLsqlFb1qeMkHJ6SaUjtq1mZZ84sx+/OoQjsKT3ybC/XyA1Ekr7YsPxAP13
E7uGwTb7WAHDe2GYIUVA/twmOlLO96/l09h9uR78wDO2S0KmGxpsZnXNBuFM6P82wcNrU5vRUyiO
9lNNoB5wd8+NLtK7qNd/cZOw6hIk+R2DmcUKqjCmDtS6Iz5LMZznMG0nh/4+AgzOBSjylqWCifYm
7CfwO2KcNyfauSIDRROxjstbD8RS+w2OdQtTk3CDVEjBowk22o5QFPcItMBacg9g05Crl3KMcMVf
Hfhqh39BCpyYCSJi12w4BD9CVI15RNocvuepNKtrT5lHl1cB0GgG65C7NAzzCqtJctHLjxj7ngL/
Fd7W7VSeCBGOyt6G8PqxlSNnaXQ9Hee+XhTa9gn8NEYc2gErGnNbEe+Gq4DVbjhexGmJn85YHTFW
UYd5UnQr/5FwqblBZ7ZrLyxS03cvJLnh29Wt7cvF09dRZ05RLcIBsYXNtS4LRIwiSrP6m2sqwsdF
Jjx0JxbBY0N/2+Rk109wrNg8M8GPSq01fRnPaGQa654vxeM5jGcXK+MOfif/tSy/ACPSjEa4J506
MW7q4fh30TsbDt7XRKlE1tHvx7HMw3SW/0SAZ5DZl01vb+ZcWVpy7hG10gNYOgY+h7WGmkD37KjZ
+tm0YgUPXRVOLQIhxNRoUToADCLIg3MCp0SIsPEVZwEUnL1zTvKgKZOEQ5Ta9GQzABFke3wIGGbq
1P+mdeD+2oGY09/DA2XJNq5SbFoP5QDk2NoJGApIZavPogeDXg3WEvek9xu2bZc05wWpI2nLNUdw
S8EFdF0qFdsr21phzmrwn3GNPrsKniE6REfXis9CiMTlG3kswrpv7FQZ88qXXM/owgC3aDotdR3G
gQGqIGCeThgpgcuSRaQgwp/cZ0/oJ3SNt4o4VVvCIUq3RiwZ+1IxGlvu/abnX5KbTmY6m6RCmHjd
ewj6DuDorNbmlAMWhj/ycnp+IjQa8CDelazgAAeihqWuODusSMR1IFJqr3FxJpCGkWlxjsUAWsRd
BjrRrdD3stTa5DWRzo9mOl+YxeqXKZxxeOMTSKDI10ciUUPJlFK13tFMlVS2apjtStpomsD3n+Wl
EPtBgpPg43G/MW7U/8EVnhL+C1thxep9Jel2VlZpnk8V6rrRVM0Pd5U1epEy00hKZIFcxzZXDyOO
s0aGcKtqUOxlSRpy/vSIbiUTyF809WCTfUvtb/E9BL1+U+huAWhtIrud09JHoxCR+VaUIPWrn3r5
AMIewUZKmNAf629rJW8lcQ/vXR6vSMqkV6peWC3Lv7V8WYhoRZOWTacmG4RuCwGrKmVGEiizhb5x
RbMVToULnUlJuDm+0Bum+HGWdEYJO5cQEzxr8HrZ0OyfELqrCOkCVr98sWVvHDNAGg28FTKGaZTz
U4tqTKDRgomVnY38hEiicEBhL85JvMOkUbPE0X8KFbLu5tkhTYukiN3XFnc13pNwHdwx7lhRKfS0
rLD3+QSX3dl+Sx1PfV9XD6ik5CZ97EDhWylF+2tWj1rrIOgK5/ia0YufCUmf6DSUlmvWQwStdFT7
dblEP6Ouug6Z83pSIT4n6eJ590zNfooAU+EyOPAKHfS2cAQWTueNu45quenocm17zM+4b9PqhqxZ
Tj3wZICkrY14sY1BpBdyvSfSM4DdgypNyoZo9oI/S9N7X4Cju3NSy20rl04G4bV70CPXhmptfR5T
hHL66L4bKhUHWSVZ+cDpUFOTQT7qseAP4c7dodY0kaCu0NLwoq/FuHTlzC77FY+nX7miFHgJ2iE4
2Eb3VoqekBBAV2tKllOmt8FHjCD3NW7t8/H8bdKMS+gsmAROq46aQxzDv94oUeb0DZUfHoa7wOCO
N3ESaMkkCDLd/btF4uhHQFiLinwEHvSG7ZFV/eBnIr6HWzSt9Ltz3wUdNz295RDb4oRd8RG3qQy8
PgWS8OvP8k9zBvwIP8dnWZwq1Ewtog8yGvcTgmIl1vO9Qr/0/H4rcyRuNLxrHb/u7Yu7kd6skKOQ
4Qnw9s5DQSjqcyVn1agOdxfrDeyfAQc1bQtvbcexpEP4cA6gnH0FGW6CTToiflm6Z/Pa8wZ/Etqt
u6YUC0OW3xmOLDetoOceh74zgcvNvoXMiIHp68ErsUm+NQqiSA38+BTw+Kmcs1EZoX6o81sd0w0a
+axqPuRtMAls768VTYqAzzlbHH1dsGTVWEQ5+UnWbBKC7/QZ9NaJZqP8JRBsjc/Jxvl5D8oMRsCi
DHOEGw/bNlBED3aPhc1ED819fgk4TmNIltn7amdx5IeAr75yQJDCSvcimyVFCvx2XV1k6mHkcTxX
SS/+bv8ZmjW9V9hGyO42ZfeMljiVAvuoHaNV8veNqy2mXbRBW/vHnn5ccpntFW7Dv7in7gFB1ReL
on8iwYzKOeq5MtaIwfEwC2qibH0QZEGLyOLCfpombRJxgDJUcpShqmNdIuN6ES8qnpCRfos0esHj
BJXEN6G3qP6dIUzDFpmM751kiooz1wsjA6PSHQnIfN+ZuGdLaCOwMdikTTlO3FM0Y2wLtrxyd4jm
da8QU4rV1udCo2J5P0FQ5zYbgJsxU7cDgJLkx0vowYDMIfrtKqDGGSf3UPE2noDi65lk2MO13TBZ
6LTj84MCMedPiPLhN07vNsauMPVoMivCflEy9N7lLenUBoBrD+qeTGXKjVJlvLahpwtmMseCg+qe
XojYqeYtKHoIUCOgiJTVcSslbqgYjn7/ztlHyFW1DEAj16AwJ8Opu/H4lc6/L083JENU2DESAc3G
1gSuZsq/ks8V/W3SOkE9povoMX3XoUHODMrEbbEBznxdnBQoXmqTBwBgmAW2e0oyWF9TgqdivwaL
+0g9zvCUhleFUFacy6oizH8hcrNicdePFvqdYJRxr0+mfTLwBaSYIePTpXlmolaJOpSyGPyZUdjb
uB3drSEpZQR9bnZdggEyyjh92W7TQTjdV4HlDXeTZXuWIyW/jtXt+2Zp5LkByKihOmh6dJlW6GLg
uTTp1b22n9ujHCucAHFWeYE/IVn1yfEiTmKqSQj0Zn7EUDdhLRAD7hHw/8rIJtFHXVwM+75C/0nq
IhwrZBYh0otOJY3PCVIZcLg5oFYtEpMpUzuHbQ7boU8soBfEDCpLj+JoVE2tlVgHjIz1n+nEQKl5
TcX0TgGm93c81L3RfmeMGm6//CMTwCT0sTXQHmxZMlKLLP5aKlN0ycOXiNFPDojhozDJNV2u5SlC
0KVm/uBQn8tRzrBfGCr8RyhovEPKRbXz0Q6nkMQxTFdnXnemf8xAp5cnH54c41ECgkxHoa7Cp+Xt
EUWrs8gtGbK5PobxRE2uIe8GvNAlBDwYgjFara/Cgji7gP7MmFjmfvOZ0HKV5Gx4u2ng/NOPZeSH
NMU5h6WGu5sDF7G3Q2bjIAqcjCNFauCuRlS4Mkaly/yv7TkypeZf6RDgDx+Y6tm7MvLqYQzJmI9R
/2zg5ol+3pSIsxsEHbqZwXUPImAmCgC/BW5qRyiS1tkBZp9KHqGX6gM2t3EFmTFJc9uc88u5TAVf
OftggLPScw5UZnDBm7ItX+l0dw3R0s70hAe5brf8Q9+xAUhlhjUU5q+/+a5Oyn9MHZpFCGBafb2k
10UAhoIFp6nKDYIgwEQ1eTcDSs5neZFOQJBjNWwrV0sxUV6Ecmj1B/bHIRDZazB6EG4i11h15Cfp
jRx0+UCsnCUvdEQdmVIy+5fxI+CgVM3ruN9US7mm4+6lxbibLo4AzWuIdRfnw2dDCfsvrfZB3/22
CdthXJQPfI25uNWGZ0tfvG/P6vXxjXOtGpZgTWIgY1VTgjz1D2jQqqeNdlvR5z1+BCg7mByfJcpp
ODQFY0jGk8fzomiT1EuH9LvPi+J0eCZ6Ap1HqjIh/p/WdoORRPlqfB+p6XZhq5nCziE/t/Z1XaxI
/1pFbjnL25jq2mR7w8LJ6oTkbeoSxZ+uLrNGxwefH5Q3C9Zz5UY95N2ffMkZK8/FnZflYzrw2byW
Mt5vFNEiU9uKif0hoELyV1Si8YgFsh9Yuy/i6Gfl/xa2TXQ+fXeebSnQA8GEWjtL+2zfJ8AIWb9I
Nt0eLEH0cgzz4kAPDzJXOwuJwz3l57U1KlbXk8KUWirVCxDFLm9/mI0XovXEQNo93oGo6vAmcu76
rIOSTDbceSt0BmIhM0YaxpBp6MqeQOJrJkEvPK2NAzoa6n6EtAZsabcFgx920OJ+3KQxL+opIljS
vs84nsWpTdD2Oh3LT9eNH0r90LSjPyakbsrMbXZPMS2RprjL0qiv7jWP9ndPi5Wkrt0CBW/VdhHB
bkH/lRcUD3TetQeg1YKqKTuJjeOujgyM3CU4ZNBsac4li50uESo9vwPOkVFDoJJLs5XqIGZDBr22
whfwqnGKaEOlUvSHcuvmQX3idKZPADnJb8fnNyZaTRkUvsfFgez4oxozW2fcR1Nb+be5868JGgmw
FOPGd8fo6McjAZZOFfNIIMxPwm4Dc2l6KjvQhY8NRWNZxh76kf1Y6VOqA9hP5CSIoQ/Z6GAHe/Ex
Vwo7Tb2Dk3nv8rQrYjzKN5Ev6IIq711uo8qeGI/LFDqI/6syi0WcPiC1j6i2BfCKvtHVWkTtxyqW
MtKMt8AaMyKQxpnAiLkx1WU34GMAtc7KAO7MV2facXn+QujaMGxYRmoS9OEuHzdvwVw51npJubdi
YzHi/HijeqsLq8P39J6885LtcPWoidDZr/XBrozOC/RQMdoX3xJm1S6VTXcqLhjEpPzw9tBlJR2w
XmvFOpeQQ/Sg1RyvGXKL7d/9syVj/BQKOosfHgILMcTn27YQTFYoV364tLSJTaJWAfyerUPTK7rm
w0tqtdWi0Voa8M9FKLk8PKasc4dzX/OfHFNrPg69ex2Ee7EzCe6lxCn9MHc4GHDc1hPGaiClR9B6
635smWdPGNft3B6ufsMY2xOX9UtKw6ijoCvnTriycA4Jb0cASP/qT3S+tg6oVxcDuRvS1XO6XVz/
AIA9zaCGwf/EspErLdy0EBscquLbwzGMom7nEYFJfRI4H+E4VPHMm/6N4P7Ae84RTWR4wQvnM3YH
7HSC6t9PaXzWAUkkb6qeEdvqCIAUaj81jK62M2a1VbYEgcVJQnfuafxg7xeHGepfJA+O4MSyhUER
uh+Vc3OPNoL0D2uWRXJS15DAW5nvotZswujBcPE6ShyaQwvpfd49EkhN2hsFxlCGP2RGcUUzAXge
qzGv+WnCBihGhe3ZmWC2v4eb95kVRAHqb8oyG+6MPdI5lDOI8ynezQFJCOpm49IUA5jn2r2pl3Oe
mTIAnS6azCxiBl3sWiz0sYfdvY/oojs/uQwp9NmCDQqL3Uiy3LEjcgTJe/PXviqhdH6TVhJvUJXw
X5MQ/1E9rCcbpQi/2ibDOU0j1qlMCrBf9wjUEezhF5arp8E307pYwfweiLwHt97SvAj4mM1p0vVf
x9zNDarwONS0QUYd81ymQmQM9SPnl5YaE30dMWZELdE8juXU6b2EH11AC+84L4tHrU/Y/TIL34UD
owCriRrNDApMz3VNrk2vqKTAho0dXDWcEwCmG1lkfvYuVwqh+u3I9cVM82umBcDGtTPO8JhW/agG
FcwD1jYRbNIjS5SBl1ftLxEBhWezCT0haGaAdweZenruxOgVqN1ttdq8U5DNEuYQaiIkdfQ1quZA
yI2PmP3OeyROs3JdjyUlb2rBbGC/K7YKFZ0xx+B/NfAowVhDwC3MuuDniKdbgqRnjb/ExTGc3F5r
quPxICHIW+5pdxxHJLc7wy7NEnke9m71WYk8Y2pSbJzfzFyVP2GWsMgt7gycoZ06pkc0HsaL33er
nRRziHrKWOzDUN+14U2+CDRa9gUIbiGwAfOHZ2kmXf5WcuCH9RjyPDm0LjBcCjBWonuF2aJlrmbW
boDPOGfm2gI38YzjD8Eq/QeRME/VjwloGOKh/PHs70EfKF99NWtvTEKA06T50hAvaOl7qyoQXDoX
yLuXA2hxXywpV7OroSilYXbOqKXkNIUKZHszEt5R5HMOe7vsVSpJR/F+r0hmNWqhM6afzzr60AhX
OFP0Trx5cPh93J7BucND5oagV7Jx6eko1D2V7k5thOGfRUmYSm/m45l+wz6OJjGyTr4+OGCiWaIw
QEfRIjVKiWmQZwMG8pP6A2Hx6521HaaHtrRURyNaOg/tNgglVrPOUuEF9+I5PorCzplQfkb3oka4
JZHu1qgzkRJRjdhXfhjEjICK9C9ZgE1RVXrBzucG1sl8oilwXFBajERpwHupdoaMNIOPI1fS1lki
O56eAP2QxaPMwg7bk0anpFbCPUPaUTdDfNA02QsElOc7xqs5+0/w+Ue+r6KSCx/poV65uDKg8328
l/pYpT+F2qHTqJzXFhDOr/OrhIxUecKwtH1syECx2NbzACvW8rvn32MN4MCDUBTVRpKv6EnC6s67
2emzFju6BE91SG/HchOeErYB2L1yqAvW3J+oi+wOi3PkiCaoMfidQBYZ+6EgkWL9w0Fq1+oKAV9h
axSXAs0IFKBVBEcaXbNSnEI5j6wcXVZkfhlm/wa/NK/eZQTKp2zA6Tii3eCpqa9bUyUrqly6dang
iXL2eGm0D8rLuItOqLWWuKq1tqA60dn6kbia21rLQWQ9I9X8Wh9B23gvh4GJ5w5Vwb0A48sJLHpw
OUB5XPm6af8zjPxXcGbnmo5vkXfhp1/FdkgJQl0Orp+OkySynaBknZy9gkYjeLZBMFK/2y7H84y2
AOuYA47GOWWMfEsnFTPk3kEpyr7IORg2pnRYf57oWNqSP0MjL1pU5HLWdlYBelyz0biQvvp1rkUZ
KU1776Rg+eFfqz0ppGex89gasrBHeUb9t2AM+sxicgEyF+jCVgnlHxM5InAwx1bLVJJ9faKlI+Fd
0If+pzYWtlOA/b1UEUvsYx7fGdA7OZTNRiFguhLKvkcwVPCte6O/DGIqoi0gOVGBhDmZPdlIwFGY
Pn3ZORUFnGqXlVhuMGKUuwoxgIfe53scnLRoTbls6Z9kQ6HzjR7Hw4QOW4VR6ZnzMJAlevju+Duq
9zPCVj04dc4D70CD6/MlRHY2pVROqiQ1UyquMquxb/P0kuWTH08m62ZbYz/S0p/hxHS0OKasZSKI
v6EFgPJmpg3GEPaVKyTCQle0/L3IFDIpUFJOP2pR2RT8W0tr3XuV2/c1AubQX2J+JNQLfGMX6moD
1Qk8JEH4UIijrRq5rVU9izZihHZjNe++BTlmnpgB959QDZCoyTfIMvmHWZcaLcmBf01p2ddxk9UR
XdohIs7Aj+oFrGbUeT5rLq8NLKyaApccVWpMvZyacRxto/+hwHxVBA4IShV8L0d3/ZDbSHVpNwoV
UoS+SUgFv77Ddc3oIATBgTVApXPiXCPqoj4rBAmsUsKThsy7+f362SK+ZgOcIOjrnrmK5m9T3VFw
X3aWwQKHfpNj2XHNrV35vPaEycljPDWNtwafQj1I8WgcTyFY4DC4uQeI35Bn7AJg/8urlyfTT65h
cgerc80QFS7GZv1nHeMudKsyx/X+3ke1nM4TRrKrxAo7ZBdqv++eCc/pNrwtFpVbQKm1tlIAW84B
Ke2WVaGjBUvnh4t8wPEHcK/sqPNGBFA4S7wq4ucZZLWeqg0x5VuFE1GGCs+rDXwF7XEjT+B/JbA1
mQuBaxQ82tv3T2WNbWGRoW+j+tB6t8oVeC7DFAAP5rj/vzcf3ldyIlA1AKsKe+ztfmHkm1nh3H/Q
Ac/jKdS8JdIHrVqxWrQo+PtIVwM8uui4b1VX2QTZ+xjSOHvhK9pgS+B0KlaAxM00kojVD5k5JRo2
SKcDDc3/r38PafWXK9WIHPEK1BI/P5CmMgtj5LtUnTDMo8mrK09RY3W8o2rahCtt0ZPIeOkbRJu/
IqYsNEl5a7ySNpVuX47XXaDvD6E/9zsHuh0Z+whpnkUeQiQgfrIT9W6WfBAWmeReYoe1c6CXduKs
m/HFJqq4ZMRVc1oZIwqbBYze8neZrgUQHBEOuCtVCOUJJmOXUrZqOhkeD3xZbJDIa9/0ECrVnq9F
0KI8z7Tne861NKCup8MpV/XBOk5qc8rppLlyOLxGq3QwHvTtGCCMhyk50is8J+r/1+O2RpGYV5pX
h0z5MLvOBd6C0f5veKjy89r4DbMZvM3bUy2vqCAGr56gUi9Crg4lG9Vk74b8AZZ6bw8vHv7VLdxB
0B3b0drzTqdieM2v/s14Glgr7LfOL1gJM6SqmjQo8Pvi/ybpQKuLcydGZg01hr9lIzApQ6dYMLbm
WjZ80MIMKDvZa6iytviGX1GUuYuLbe2RL295YQfibxDPbrzmYo9/bRAtmzEXBLyIVzN7OoIQHX3k
CTyv2wXlSph1Y3BFvPcVGaZ3VM+LdW7DoD58cPmZ+cJrUsVbO1EKncfFj+hvj0OeXw3kDhQUMBlH
oxuOg4v1iIvXeWpRuzuO/2OZ8fu1GmBO+uwVgCmO3HkQtejNgDYmdki1/4FvSr6nU+jsLnM+3msW
OiWDIrV7jfLhENd0zOF5MQ6hkh3j6kH56IYBRccAZ2sVGAfZioRy8aFPjTwJD3QRDUTqjQzx73fv
PAi4H0ugpn9oJS55QSSSo868Tpmrssu9q1up1H4xaKuvdzsU+VIqGuldYsQ3nw1I+GWw28Oxy/e+
5Rvq9CLr2TGXPzw2VxB2ZRYFdgnVyS7SE9I/I5yZQlhOP7s2XZRMdn4R2OcZ0nH6mcsiiWM6w04o
k9nSyrUkgyiVLhKzGgJjz/KKQRsiTetIlS0jNHQPbhCwzf4tm9+Z07dg4UJotDuc8KidO1ii06zS
4XEVhNSycurCTqVvpoBOfK+lGbxJ1bSuYzxMDjEG8Fxl10OeWPqUAASC03A0Kr22QqEgOhFHqWJ+
pObrfrjSFog9jtmwqpjTqRKamzkrQhHvGDHqmu1VYfCSz7s/eKjNJFvPZF3s8IJJjGDQgTsHBoLp
LGVpI2EAKsRfMrQ2v2WE2JCdXE7iPWw50J+JBN3JeKDe/rqv4CVrUal4gaTsyYrDDAJGkkkKRvHG
AcHCqKg9c1uOiifZe71XeW5ybfGaXas3bmxAng8f6+Floipa9VaX+sbrShGMdZw+4Mg0P1lyKPwp
0ZYh2/tv8pTMk3jPif+Yno8IKS0LoIM2w17O/2pCgqVWjeVvBXG8qBpUMy/2QHDlgH3W1gNLQBD7
XsfnYYbX9Rdo1eHYmxVTAS4bSx2zwEA/QKeAAeMvoRUnplEa9YUup/I548uVGPfSiX4MGEhJ8i9p
UN6fOiftxDtJ4u3zBIT5TVLGSwKueb9HvbNnt0oB3xIXXkEutV4AtTsHaacs3j1jblsvxoZLRIXA
BHOtxz0Fcr7A3MUgdZFx0soW86z9QwVeaRXZufDHRi/ibDRaZBBGGLsblkwHOdmtWq/r6eQNfZy+
pisxQ5V0XgwNw1riQSHu8DmpC5UJqy9WB9xsF7YaI7RSPidzbOvuAnc8/z2Uw1L2ovTOM3AuAFRC
wD7Vsp5WuaFibaHoCiqF5x86duvmMPgzvjaIBzl/ecG6DDVGT+uQxhTqvpe4ufdve/iBEutGSWcZ
CVCDycQc5SRs0D3xFmmfU0nZirk8nms/dR8SIByXrAVDlSmCz72g/moRjRVKLEi5uhcQG27yD4sF
8S1EjH0NcI86psl9cTVjGwlOfSHIVjhfhlq5VIjzB8Ty3cfDczNmhE6rJ//8eT8AGHz805SnyTdr
N9K3/XhgfUj6seGn6dye11jpTNSNwO16zIheFgb6JnPoPqFCwQP5Frzpg58REuEED3R1uE97xXzJ
OQIFc1tRowDqqdJgnHbDO9/ikptDSIl1Wd6Pa2WMqgFiOdSNAG3IkU3I0IL0mJFZ4zxKGdjtrFGg
IGz9opdiuvgxHpEyVPGhhXjcEgpCpZX5kJRl3tdg2dXktX9fbupwuxphzgjBB0B99gFZCqMyrvuY
wnLqRnXs1KVdGVi9BfH6CjhpyE+8zn68sv3S65Q1eJx/lKYupink/Y6IOheSAseQ4YPk7lokdDkV
kLl860k1G6wOf9e48DLV9krzxl+3CvXe6MvXu0evdFJQd0QBR91wUPzEts7PK/jwh2/gJl5S5/n4
M0mBw0cFHnOuOeoAqt8Tlgh78j1sJ6cAOoNNoGvY2zFkIa/I3MM20BP6ADQ3Jt6F7ITs1e7spj+1
IagaOB/0LBCztBLGVA8gdIzohDjc9U6nMSPFhZqP764XVFDjWO5nMqYqafufcpDOcYs4NfkW3sWZ
DFjJevFjo9tJvSARVsbg8bzt2S3yqQAvLziC15d7R0ekhQO8CaELpuqVwGjrcpe6XZYhgtBi18Lk
WRUGFsGCvAbIlFbPgWCioibny2ah4xy3wq4+/ApLR66SmIYwphegaQxR2gZ0YzxOAu6qKflMcJ69
2wPvbFtCGnWiRazxuvJ6Vuuz01AIOsHfaUBpsegcDFa7Ssjl6P3qc6zBzlJt0jH5tF7lY5VlZNlH
zhOigMW33/R9V2duG76qf2mcbUp1eNoxTBEiOuaiVna13kFWrkkjYMCbzZ2imJpjQliQ9TPM4qiw
gao9NSHySZPYMn7NtrY4b4CSgnET+m8pHVnyvizy11+pEnQUs86O4hoOacc/vnH09bjsTktIxBsb
uY2mrBTlFJvgJ9CsuWm+Sck42BBunZN5cta2OlUSIGi1n9BzXU2mBIvxkUX76DIEad4kC7sdEE9P
BV+nysRctW7RShrKM1qtTLdXzsIp/Pz6P8xXGb8qRuuNs/p/eaR9dShOWpeC435GzdoWJcVAQKkW
9PRAA89rOJD/JVo5pUDYpgJvmVse4tcuJZY3oG6sIPqYC+hPqbO9ZjEmtmzVhXtgW9JSAC4g54am
KbSgdfC8xIIh0LXSKCNAY5YoBnAMCg5ncbGUD9V23Of2bt9TR1xICpG/bibWyusIUjsEyrTHd7IB
wUKBW/8dCPIJeQYd1Ii9osbwm6atSgfUFup2SVTAejpWqkhtXE7th/9zU9lhS4Eu+7G6pX//juB9
FMWv+QBbXiZNAnFpXNpHm5OfUx8OqQcZ1rqWelkXzOcLJVa3Z+DZiggAHYuTQFQF95UkecbjL+Tm
eZmyhmqGacdjEZNbK1CqTrSWOdaA2Pz7JJW62Dsko0y/i634LIOty7wv0zt7d2w5P8YdT/6SGw8y
DPLwam7fp3eUxCNly27p3j0H5YXpLayrCsNFcyTChbRo3ipTjAdFk9SlkrBeeVboOvImqRzsbkAk
q2KpyPvLRyF39iiRw1t3hHaF3p7k79Q2pH9eu31GAntUQYYka90gvVriMvsBCOowDZYSCC9uw1wr
QL//h6LB+0KY1aAAKOjNgiM//ApaEfhNhf3v+ye+FHLR2+7Cq2XFbUFaZfNrvADJKeF8a9lVRP+V
Ve9jEng8dMSpF1PXrOC0IHryOHprWkkr3xKOk4VtR6gm3+Sb1GqKh4EiHvhhI2aAUscyjRfQYfpg
i0aYYmpOU9EjSZT8vAg6QKDLEtwQniuzmADr1H/nXyiIaMTqkZq7pEQ9bdoa1tIUbKpaad3II/W8
WV6D5VDAnEFdyqT9Dcc50eTEh31Uaj+zlrz1N8pAXkDySHW01gjHnAMhYGad6oxvdij+pkZBcYxy
GLv23yLF2UVIs8gFHaVMd6KiKRrXE0CL6cH2HLeZFSOh8h+10xAouB2EcwzRQu3uBejB2MoljFmB
lA5HF7tbVJikS53PSnCWPFjX0D1vocHAzg29K9QuUoSkaj2oJC9kQHhIp9QC0oOu1miuePPvkHzy
Hyi8HQrRHJGVDAuTSjAKLqjx6V5peEpTlrjMWAhnKlnVFLbD2M77FEiWmvFAcAT5Lfwa/1DEhvNi
Txjpg+ls/BiuNw97IPC3z3vBXPxDYAYC6sX+daKUij03+BOzEAy6ufm6XNyAgPyDx8C6wOVeG3ue
INq/pKMnd3MgY7BKyxLfD8d3Gu4p0ZgIYc4zvpAVERZZlb7iMPYl6j5L+g0m/M6n5eH9Wjn9+ugw
hbtPCoo7QXqZ2Ks6G3HUMTU5ERo8aBxuYiX9K65Qyzdy9Ge93QNoe5bcRj9IDjxMlwXV0O+yYJOB
S1n3YHRL/MLMBwEcRaL98C2D3JZnXAKH3PzLLQ3S5sU9/x+2W5wFhdA9uNhK3juKuWq6Cv0pAwqZ
z0p8bhCjBTmHRXtByl39biaxIIaYrMNBbyTI1gqdymF811zTvtcnN/50TNw/g/smUumRytF7KWpd
nsOCkBZJYN6xJNS5RrjWAQ8ic2Yxuq2krzqlV7f9XIIA548qdLHNPH7BlQhgraW58P5YM7ZXSw8t
ZYwEWxuG0Q3/sSSabJ7GT98hiY9EpKXIkkVp3XjXpVWrEoMV49RBdSbSlSEV8lRhuOABw2glpFmD
KLbOPi2zNNwVwQt9adYwTosmtWHtdOl7F9xXg6nCISG5AP1G0eWb41pHooIR/Zzto+6X5CP5g9d5
ZOUHxgXUf+cHiIf887M8Fhs8ZtFKck+EkOm7flgoCYQ+meNNTqbnlw0Th5s+brCCyXS4AKeNxr3C
kPi/CRTVTA/AezCJ94dpk9400UzOgbO1MM0LruaJvRjwN5K+XdM0zFKE1gg7MahjZZj1lYxBB84r
HHWg2ki8ucsxhvKf2NFsfb7Lws1jqwIv2IJo4Y95PFVNk4uaWgoZn8VU2X8+YtzTXOzxrKc/fBcq
6k0ut/vgCD8GuR77IqQE9xQ+sVndmdEjwlm9yi78y68UVrvB1hFSD1vPVxS23cEljz5vovNccbi6
eoMFERAZ9WtLw31odqOe/Fez2uF2wyDVDVAMpTn/smQFjLw5zaPoehb3b6cs0Ez6OG3kdnvEoWSY
/PgQwyvmZRhasKnIGydICWkVGVndPdxXj+qJ+XQbA0pU+9R2WE1qWnHXC4QVvCODtw7wI9GW9npY
Y8ce0TGr+kVim6/CllyeiLavIoz/Ea4tdpv/7YNHgUJ8d8l4UbbD9NoSowJhhHs8pjmdy0JBwWar
K3cnP87vXzEqvkB517PTTzs2PzZnTPAcZ7tcGKiwZHq5ZvkZSg7vnNwE1bePCanl6I4GcEVxmhe0
IZAYfHJIumCuMq01gC4OR1N78RzxtwwFtmmjpL50QS03nBdziHQ8jnGO3pUWVQxGb5GBDwOTKbKX
YWW5NhL6TzDhjqT33yTMBMPqT6OyKqWonDBnW6hSVc1li6ou7ipmROvBYxWuhxZOBenLyNL0XBlc
KtBUCx/AUupXFVezvqHtJkHCMVlthvr8mph/tyRRYsxY2q/2PiatW1QpZceBRmAsztvR36XWVXvW
2lCDHhBZTxDzXpzAQn+gQAOz+kjw8LP3lfiMZ8m1o4lva1u6NMdL/qAuZvRjFldtHK/y40AzOAb5
AE9Ei4Gmag35r6+ZS19Cop49QKqwQHnUFVaL+8mmeo+yUmsBIhk71Z0kb2x3GIo3D7fJs3irPw2x
aS7w9npyU3BZ4aNwDI9tzNPStrZfkMlOeZFsvKhaSKCKqkII6+EwJcH7PIzR9HYvL36iRcAkK6fU
UM8/0lyygtHr2ymaXq3T5/G3dsJwMw26NnSqdBin2aC8WZRgYvNuQN4F97mXXvYYhzc+AyO4UJhN
8Z6ipkmpAr1Qx4u3pwIS7ZTIe+C2ViiqpiSor3xNb/9WeIAxcghLIj3DyN5h7rmSMlkzKNv90xWz
vMQjC0L4x1AIhzgUfh38c3OyhbPHolFSjZOtqq3FC48+eXdOjjLeD3nvWmVts6nLPc22o+YBoQhl
TLOfHdSDTGiSwxUnn7TCUJMrGWhAuVYQXFguYWCiR+YZQy7pJiz6rembo1ydUYKcqowa7kduvMXZ
kSxIislP/gNVBKMCi6VqYt2DPUIIpW/RVSdIRJkbCTLyrOnJMh612b9WzRChzjmXoXPox3gFFNeb
x66Nd9RYXwDqVJDj+ClW7pA19V+Hwf2tfu+EGAEua1lu2H5aUge/wH2AKyNqJNjYvAdqw7bEmO6n
ec2hexCdPTfwyZPgsi/T42+Oa/k5k47KFcZpy163BSemUBBFu2ePYyT+H8FML3xkYzPycHCw7yGr
e6VCWQl5oJ96iFu4LreZt6eKK3kH2lQzv/4Yqrkwxpykv+15qZaknf56TVIcK8CCFp2tgacA+vtq
hJnrnF/jxaSDqDIKbytC+Q3DmJ3Jk9/93gCip4QHvoLqf++TRe3PlvvveckHu8pgNWY1I3hvw8by
6V4nTQGzLLNp5wbkPyERpMbzMIhg92M4/0bgIu/efGkhkVKcBD+s5RX/qPArm5ehHuLlzLUEV9y+
RzZerOSc/8uUSWCdQzG56YVyu+0KUwoIqAtlzWfPWIFk+QsKZfQjOAW8LraVB3uzM92ZJd6HrBRR
2zGwnDyU8SfulJKTycUsPSgQw4xHmO6j4CNZxkmPfVB2RsPERgPgLimDUAPRGZA/5VefJfFET/mM
j+6XyaI8/aMGIHCcN8DjGFSKF02RJ2j7VIW/EBPC2fV/KlTBsEbSF3tUR1YzdHv8snpLO762+8tQ
SfiZdKD6X8sqJwSVtNAo9oEAt5EKuI2NSYl2M8LWO7JA2TlWjCeAPSiaIOrDyoPxlSrCbdNlqmrr
29viheeL5ab4DUXdq7n8BiSDgMoX7Wz+3LlMrmz1drdoO5Vl6aWDQNE0u0Hp4EbMHpRwf4lNcC0X
nuqXglfBtGeoNilPcMterq8JqKmV1nkzyaMPKyf4IsXF+t3KkV37QNJAmq7nBHM4r0cEtXG2EcVL
CrEQevSp5ljeiYBuVWSLaNxx6aZDYFrY94eirW+mtB/7yZ/FmsCUrvGwYnj+INWxS5WYZOIPSg3z
y2DSjkRmLwRIBbGhXkzYFDB27uthFin3p8CiR8TtW8B+nBwXcqRDYG2SpQ6Md4K5diqeKTbzouTA
VwVENYixi0YZZyYgD/mgBHx81RM098Tk8y3g/0WEq0X8/ZSmoVo9q0leT0qZAfeq8Xdei0Rf64rg
VQMTWODI5zsQencbo4bEY8GXEzS/C9vDGuRsGJG4u9LL5+qr3G0Mhu/viaja0J7lC2myrUm+jbYt
nYueGCHc0czWTNW3IJ0MNQx3VIvCjCddz+Lb+XoAioptZHydyOb6PQyPgVPOuha2PENcajHklhdx
kOCrf1KivSSNqDV8F7SyJpmNlK6hdbq47XmbOwDw4JedpiyCKVYVs3MJw4/Vc1uRctuEoVDWZ0Yl
ba705oDCroXYFh48jA97Nx2oi9B1khMLci9bUsln4y9cvHCULFlxahSJa/Pd3dqy71EtZGc7jqCR
Y31upSim0Y2Az+nFBDKufLrlYmRTYdmEIdnilbaVAdUtvrW9/wynSU7eD+SdUErXS+7EP3xWYWAf
IgV/udO3YkHUFDLzL9ydmSuBFo4FqsB0G972XcZBdCdjBuQzrO/0m2Q3s6lJ44ZMkv/UMXmuraTm
Frm9+vk22xZBE7xPMuG+jK6B1OS9OUHqWeBwSA+ssajIuuWCll0ELIc8mZuXyWorkaoejOrCUsfU
DqcOYTexSYDvCLKvBzSQ+YpaIqEteXdWimL4j/dSHqOQJOJbxFKBAZW8xw6BjOIlkfE3dGw7WbVf
bf2TSp9eN8ms9hMSS6Cgk3zSRaYSqahTGy7rRSfSI+iw3kq4+2BY6VBsiwwBad5p79QqnS1yxbex
oSxrM9+acEWJ7IRTplA1Re1/n1ULw8qKv35PsIhx/yB6nNDnvHls+FnAV/As0Fx91pNo4Ysun31X
JFRt9p+zhnamfPjRu9IxI/nrmVKVLRfimGJNjexrAyhK/Z6dSWQQG4jKO/wYNVuGd3x8oOhNGbzY
nPt8urudYnoBRf0celay60c/lj0LRumXw4v08tsfUTok+klbD159jN9/kLvsHVPkcONErAYoUavU
HTj+iNQxylugj+bofi7k0zFchYAZWLN4k0Lq23QiThDLlb3XLwUlHkoAbQx7sCXPmIQUDDimtpg8
tP8xsVdQe8r2yw+Tl8Ix6szZXOvA9fp9tOG/ZOgDag+TxGbIK+AwsHvB9kj1C75PC20MW6x97/3S
u5ozv5p0uO6SlAjfDJwosuZghlRhwwtqPIMh20OqW3Ppet6Q9HFzQ5q4MA5XJkwvgBacamzk0+3t
fRcR73/XGmKyZmIbnZGH+z3p7tgnq4f9mtkwSdDT5Ur27kvb5NJ9ocgJNrQT8meVLQul7RCUZDMU
Zjr2o2NS/ExtGblrxUp2pKIc8siHejEdfAHilYQCGDjhFRee/EB1RjEJ4dvKUcJ0TRioNnQ1sgg/
BtpyZ5AHQH1RYOPZACFRx8u1ljGRzaLuAr9z7WqJoTFNsz/NPg6uUEY3zpwEoGuwJXYtG9Ez9R0h
fMMSFhcQ7RX2FmCn88yk2wtm7hc9MI7Y6PrWEhy/5JcbihZBx84O453MFM7n/FfIUhJajeBgN4dW
fErQsIKrMQtCatqrgcG0vhCIk4Ejy6BQPm2DpSVHuS8GUwmFZsiz3C1xbdmQvzJ0UTq5nBqOJnXF
SlWHEZhH5Bwb7cXP6GYbEeebs+pLK0cJsx4Dx6tla5LaWE/u4VPV7f0sDO1/OAQfEqvCGKLEJ5nv
EXC3QGPsWaLVyN6l1Bz4mKLVgncvqx/u6fdNNLH6KB2kf0cePiMYTTvHMfL3tHk4eoIO0ZNJ91U1
Ke2EsLUJR0veo7o6BrxtR/j41yOE9DFay5smEfbwx3kjjYJbLk821dYf0yFXaSIF+fneskD0AZ6t
4VY1F0JBmv5NbIu+46yyvH9O2He1IkCFKjaAEdiP3bvSpXiz+cMrWI0UOMrdvXMGaaqcj809w327
/57LolzhAnCaOzt53i1XuqbR+nFLq7ZDdKRtS2EZ79Yg+solZu66hjL1r+h30eC/g+VFteD3sCls
1sl1epDpNWLyFPlc550WKvcU8rihR2bbHTcpIdp7udY3ORPTjIP05u00DFQGb2+mqoxEnPSCEN8S
9SZnLks6bMQbQkp7ohuvrdnu7/J70I5/v04j0E6QKkZ4iKgzBOaOud6WMNxeK8DZJvM3aYM87xwi
KWACexJAGzey6VtteShXfwozX7WK6xlEm9lqAsUxoyHfSnCw2+tbeFm6FdwCUmabTNCtebqHVema
nqJbc1AjfND+vQEQ6AOwflNBvziLUBeCm3AknRENTkqfzhB/NaplgP/USd9AsRQzHYTIUajjERQ3
u83CrvVyN8ianAeGk2b78TVzqsIyI8RD5T1+Qiz42L/rI3UaVvn95vJNiWkRMduEpVZa+EAxvMff
uGZk3VOQz4R1FOTtRhVUoII7f+8tR6xKUUBPk732S4P8AbP1HWWNM3G+ABupGQHqrrcr6bHC9aWx
dLEFbkvmUG3vWe29Q8AXTpEJxgUhCda/NDMbG/pvffTMxrXbQbcyo9E8upww05GYMsgT7wSSS73S
6riIDPsM6u8S64uSQmlsQVG9lC+Vds9TJvVmIJ44PT2yUBlEpnwuec7zy6DjYqkxs358b6EtX1Hm
kUj04dEIFxUNHMZM4v4nCnZUlvrd7L4qPJsytDaTSRZOdijDz+nBdTkTAYGikIErlq+Z69Br9oIW
4KJ/6zXK5G+T5c7CyIpsuHUsjK9cFel/AGCA9YYILEcdlx8mxgAiw2+2YAGjjZJ+nkMuSJRlhJNU
ckzKYcB8VThxshM2KujrSCgWRC3ZERMedtZEsF6w80DIKfY/pEKibIVYW128LgCoxROIU1Xuqhef
YZRoHj3Iuu7igtYtZ2RmWDPW74agryAZj31hm2kLZpxTOe37z1t1lbkRdaeoTuMqYpWHuwslzqtv
W/fMrtNyab5fEk2a2WjZe8a0nf1JkbiMjF3T4z3Aj3kmbR4xA10xqvZxnH5ha2qW0MctaHVsN6eP
ngyzvhQgClRvhOEVjNyJd9Oc5UI7RU5NsuYC3e/fOk2itIs5Jvf3haJ6n/yq/uAV/nvWqZzN1ZaI
6nnB9kt1j+5OoOLF4RLnCpIBa3Cc6YYePiz2uj5LR+nXVOxcH4x86y0TlFgrFZFE2NKLi2IaJx1w
T2kvjBFb7uuRnipbla3lRqiNcq8Qmy5lK0ZBy5XhHEXocJ3VLlWMiHmDCfnUurgDCAbTzmgGQWxf
EZDupwzw9RJ0fSrOUs+qsd+5jWAjs6XdW0EAUvPMPMWvpU+njNAJW11I2txVNdDG+FCzX4dCkhh6
vGxqMVR5rxVz/YJWTKHR+gBGN/QXHIjr1FsvluQGACOHEQtPIDnNUDEYY6Y98vuJqA36iHA32ukr
9lCEO99owsrSz7X+IoTiM2K49D7m4oqFXmXrgTWH/seoNvKq6jEAfJxAbSDcllz/3Ix8XLLNJ+Wh
SVG0XTUuQFQFl9wJTSLHjOfgwKD0x3M3oQBQ2izzgBqMgxFG3dQCVcSXSoYU4ifAyA0t6JTXvogI
dpV0nPBVb7pgAL0UA0z8TLn28wdSV/pen2BPCQKzVka7FiwwiEVza0KPxeESzzRlcjCoZYKVHjLj
+jk+G2wnYG2JkG69iWt4eLiVrMbF5SsK+XcHujC2PT+mJ1Uk7LF64utxHysbAJSY3gzZNmhOP8P4
WEabVu6FdB8COqkrUkfoBK5KQcbziKQGcw5ofE30QI/AuU7nOs9YQ5oD2CQ4q+S2wvHOWv+NPvVq
+LAtWNewPMXE2mE2Aa4nS3tDKlYbsFM+iWaQ/e9fSZb4w+wGgwk7UbSyX1H3EJFoFNO2g50WrtNf
fSuJMD7qElUq7n3uHZDgYqI3zCNToT6GfBqyumfVor9/JI74NOYVLvqEAF1vHGBmmK13cN8DhdG/
lc7jzctdMDAPLJtJpFEgqpmX1Tiz5CCTDIgLia9Eb7qBxhUHMOg63QSDrWfT7MOgzrxSzTd9/KhH
Td7EtexXxEWEY7b4Vq+V5LhRlwEqCdOLFg4O7vCX5Xrb7ilCgiZADlMmIe2ZgZ4tqddGjWZsEh9c
KGXG5Oiz97CsW61jceu6yX6MN7/wOJtA0mkFC/NhQdM+/eIAUrDBi0lLltZ8c7y15lnJ2yrrrPpE
9lNQkFTmATTTW9RNB9jW+fO5H1MZqrt8TDqXTVjoi/Vv2jKGQRXNCbeTi/EmgvDfwHl8xc1NoX3Q
FyS2u5Q1hffswh6T1g+bROuA+p2I4GFEesZ5qp0qHfEgDtoToRKiPOU1qQbosteqVaj0JvwfU8hb
71xGYazw3OZbuz1EwnUjo95ht8b3tT2A2xhhyvQvpef/GlVUR90/ZoAdTyJM9oG0CXcmAcra41Kt
HX25W/FMtSyJoEyUSyTTib4AnAvQsmZz3W2AyFzFewkQeJLcRZGUGytihu3qPPxzzyrNkloEE1Jr
6jkIcv/VW1qc+ierG46qR8HLjtkOYbm+1hpb1bcIsDUhoHUrxk77XtPF6d0nmlp+EySAFhqGJQfe
Q6wFO73i8VcWN5mXZ44iQuVrZZSJPaZaw+2UT0qWCg8Nm2ZfkGChyaDEDwFP6Scg8uxZysh3s8US
fZ9dJ565Mh25KdUPdnMcwurvtok07Q4gYU89g9YPwzeMlYX7fiSacfGByLOFj0wx2bAkYvYKHRt9
jXktEwCgp/o1hKCJTfEHPsE2H+nCpqLghyVDTyV5E4RNrafvjYBpAO0U3JLy4uqP5kalTfoNh89X
zuSgrNSlzwgzGNPbfRfOmLSR2N6II+5KinRs41w11ro2puDXFdwbYT3LMV4xrSY4MOBxkUYIqFwq
5/ZAVBpgWON33q7MjMdXM+2Vj4Wxqa+t4srwezq5EhI6s0L1kYeCxz8bHDf3UW0MPwt8AbTmSF+/
d0L+p3ChJI5xsp7a4oKmnSA1ttc+OnKBO5W+1ImzOLpgO0BEkzzpjW7J0JEpiA6aS9ProeKnTdWa
vSQBPxXDfnhpTgHnnH6T/N3PZcT/pFbUQ6qfuM/UR9mK38NDG73FOolF055ChpKeQ07PkCxGHmHL
J2wIABnkvDUtW7gtDK7MtPSfW+CPYhoP0LpRbUMk47LZRUx6NEuA8AONHwJyiaHDgXeXwIUp/0ds
rsYB6gjb8/K8lNy1gihPGmr/nB/+t0HFV+K2hmfeJizxysFa+g47cD4PMF6c8OLHUDeWwiDAGoNn
NESDwnVW2T8Rkx903QXmUZ3rd9UkEWz1Y23cwQ0z9IFgqzjsJFjalPuo77hvnEXNWMNS9IWGQhGL
ryL3EUsJwOHsAmuldsTWGsNXYeag7JMtTrURIE6V5GtCYjsKY2i52eDii7bCPXQ1ZN4/7c/CG8kc
gWPnQAhboTaMpqyOq8bqXHZj8tAteMlYXG5+AF1sHqz+yXY0c+CXn3aSDqI42va0tBIoBMVn1hsM
2qmeCVBw4ZTM3VxkqseclgamwHLWy9V1QAE4VntCdFoa4PE+o6QNJby1My4W2J655e6auuVWmKzJ
qPVsBNPo/vJudXQ16aDkcTyEUuiEr6FHN1MSpiT3EC0D0JqIBahFyAGAe+LdjjaOziJ7HOvstVc9
mCYOiFNU5bydNp/zJrgCQVT6kML7YPY9MguMoKO31PojZUno0v+GfB8J1zbyWYA/RI2gB86U0RYZ
qodE4AW57v/P4VFCN3svsBHLQuY2VbLPM6gA59zL135SdTVK6mmZTt3w6J6kQM+XdYVeIgvIw4vS
KMPE1r613wy9t6tV2PTSSh8sYpjTkK+1+rEvRv5ZJ/90A5piqY9L9HyFoQZl8Fecm2Yl4bB08zkC
iOZUSO6va17zqedwaMLcCcNwvODELPEMAuOOOUOxTyA2KN0mCsBjpRdoXOVmx/HlP9FNdwoKf0uC
PnhT1inWAZNVqLPmRv+mzmnS1iKrHHMZePtZ4FYYRVeLosHRVr0BDXXdOSEf90UtvWWuq6+c/nUA
qwzr2kOdF66Cpa/S4+ZOhSLMcAOF+1X7ztfmVhhFCxEzIKeB9ZxA2SUsLT5cgNLwqbXVUMEl5xFw
gdJ+Qni00+x8z8Ld7YSGwq0IeAVJPpDzel9Ec2z9j38NH/0+lqnuLD/86hDNZXtZQ2tE/5CXpgJj
rlebgap50draPt0vr3y5AxuWCZLpLJXX+Wd2A1IwbOgHrJwO91IiDtC6bp7KN2WBpP3qN5AOlTDH
B0vCPYDjkpBwkE5V7PweDEPQEH2MaUId0oZ6Q828I95NX8cBSP3BlkRDaW/iJUvI9mgQCttBDhOm
7AUBqP3JOqOQyqe1ewNupMa+MJdYUne7N2jR4z2Gle6kszhYdQB0kdZlFMGvzZwzlGkfb25rNDxN
cjecFdze+ncmdRjtcBaQhtwwPzNyuPl46hkhEHNuEBOitOgOSeGVp5vw1nA1nX0SbTUqSdi6qtMb
H5FPqm0n9hOQqOBm6vH/CP58+zPXMgDFAQhmXd67y17l+R09kF4OnSxn1xdVIF2NzngNVnkGNXST
C3kwQzFLH208NeZzXCErdJKVlruXTDa6IZq+6MN53LPMKThvIwmTIYYoVkxG0bCtJLV8KydAtCgu
a/OesyildyUMQiwUvtIbb/OGHp9+j6FCZtTVpTq0QmWv+9lTxZNGLcC9ZJo4wsyN87aeLNjf5/Sk
7nKYHZh/tLcZJZImxZvdUqRjowGjCRAf0P2bVpMGbn/7Q7gNqgl7JJbt26ClMrxa2GpZbXNDEILk
CBdBx91W84I2O0UE/Z1750ye6DJKGNuX0yjqNq+HxNmPQgAnoTKeMcuzKwJ+4p4UVwaTHpBOpVun
EQyZrvlvA18vJ7xXyevm6GNVMTQUSg3ifrdD5ehKCiYPE0Bs8dHCNBdMrQcF4N/exuze5jMqT540
N7w0S8goyCONK36dQe89F8JsNGAJOWHr0q5f8gUMHJxkdcHEaCGbr31K3FI8usCXDstOywq2POsE
idcBg63nMd6wHpV2PSU3NfmvVRzC/vlc0EcDi7L/5fLk/JCTbYly25Mtqd6oLdne1pIcN9zSdDsU
z79u8tpsGx+cWQxoaxNfs39YWQAXfn6nGhZ2Hj6qdY19dUdPRWyJSNBnaO5uz9wBkpwUIymb5j9Z
mUEKk4bTALoega8Q0JbQm4EG0U2p5fV4avK+h2UKKO8Ew/ejKiuAR7uIOndAgbWT+mqzoTQsZJIF
PnHfjV4yKOB+cKOGvwGvjIVIkYibSVKW1WDvaCqUJq37tCi05VAiBbwhtOeMjmDtSj8XBw+leZzk
hJOUS9T65tSlao7typFhqzB5wyUZW4PJXwllcZ7BFBav+17/SUWdplmfj2l5GG7gGXihuLX3RpuZ
S5npJ9c8NnP25aNwAZUSowuLnv5BccDNB7lKk2FUcVGMCJhAvbtQrPgwq9ycuw1Z4SXHRRXdRKGG
atpvjv3jC9Ubyx38bNix0ise2xsolZmRL/UFbHX24VmXuyRVuxBWfI3R1Sbr2gSVVChsTFUatuqk
o/jlILxKaPuIHeUHcrty9VZWFw5jqc30oMD1rheQ+4Y0GV42gggYtjSvCNpbVfk9Vzk51bEMdD50
kitr//BA7JDa5SFHBHHm9R36a0id1equXdGGLaupn75ZzH2qAMVy0ll0zGSkFO2KkCUlT3xbUveh
CIQ8xkbqopKF+yLGZmolLT1V6e/0csiry0XjhBnvzzdw0AkNtw6NwYtmMPbJcj6yNSQDbrOnySse
VwVvwHqcMwMtVK5+N+znsXCVg+hE6IQzRNEU70WXf9HepjMaaA9XJ28Zs/68LXHjsQ7SY6d8A6+y
Jm/QqQl9Sh1bBiNnMkn7ud16iXwOVWW+XVFVjw76QRpBNoQrDucNlXOQEl3NFQKiyw+3osEx+Dnx
ad7JxHeKYGKY3KnSWOu4QaMMAC5xlvePxOhf/TaX1noSDVRWba4aeemJ2rEK0iK+zp4wKIXya6rE
PuYvOvw73Ea9zPrFehVNrx9x4asy84iujAJgWC3v9X0p0VsK28hQurJPUVlmocVFp8/zP2KwgolI
+jto3PYA+FuJU/GZlGuqHv0spBRVJ02v/N59UxsZpJLyb2+xEaVi9L5SZBoBK67gcFpdEzt4D23n
JA7x+M9CR0gpVu5TNVFvxMOQ0RsLpbZu6ki0RZfSNJ3jAgE5lVet2jFADdMtaSNBSFXhjAxq3JDT
5D3wH6N1i6sMSwyqFpvi18IQgYLKzO1BsyEEkFevwm1h7aVwN5LVirHAmvJLvoKCNniL+RspYQhW
mWFiMSaP9HTFci/pmJRsiwGzYO4yzFLMNc67ITmn5Bs273+n3O9/sYLyl6oZpjxyEuJLn0VjftG3
iqBShkJWPyPGwZnJI47+nw9azFvM3m5aitomblkp1oLrbRAhJHMjLuNTyBvL7Bmjj8159izw47q5
8DTDXLoYqdQBBy6tmxxasbhQEGNb0+tq+7/u9po/4CATPUYI6QzdJJHOCL4cTPZXj8LpcoDlytcC
GFVdKnJBSLrCip5hYJ85OzLG1V10ZilqJLRhp+u8H+EkS56Ox669tBkLWFEQhtbp+qfXUfHIFbkh
SpEEBxbvdeozZmyODkASj72dUix7Hnfym00xjI0cwcfr21PmWFpcDpgh0U2AK3Ns0xD2Cu/pGgxm
LqogznR8gYxIB0Lb3u5ciLlGEkrpA9+ri1X3A741Z2o+Q4lWVf7FptxoB0Yt+zauuHF41E9x6j21
fnILM9r7zHbtq/6BTLptPKYR+mtLB7feiYn6blviOwXtBzHHzGWIHJc19DmfLe5JnkVJbTYG84k6
RNN95n5JBy+SVR9z6oP9fiApMb+c7vi74S2DiJzfia0GgaxGnGAVvBN++e0nmKOqa6KDlVZNl/Ro
RE/2jRdiz6SJF0AP7uFT4vGBvzUykfkGUo/ag1MuH0YDdvWyNLVQst0uY65VUwyh5bjxUmDh+wrI
93r1PvS/lsJBwzN6u/G4Bcxm8bBmp4qybDs1cYpVvt8z2h7rXRVrIGdwCJKmBnrL7ptbZW/X+vNO
mMI4dQrfTktzkCdu+lzo9pw6ntBdI8Y1SNtFoDNEsw480NMJYyUoD9q55H4J8g3H9HQixHdhxww5
RPd2FKpxJIKVafCghOM2lPI/3FElwkpT5n0r8zf6wP/+FjZcpYuW71nFqXHTAdLABNPIe71NyJi3
/5mDhg25bZvkTQJpc7fU6g+nkBWN13JeoufTStX136rA4NqwRVu84J0hY1BCBu+i3C/6tt/u7pKZ
Vx3MR6DtGUwDNpvOdDO1FC3d04Cwts086CUUMEhIrb1AE79TXndTy+cbMyA1vv0m25CAjFaBdme7
CS19x/srfVi4M7emwc7AVQNIP/ZJPw9TtF4quowjm6Ie6grAoAw3YUeN6rrrHh0oh6PPA3H5uZOr
UTSrJmxQklhrMduTvGsCtMQWhLMmhOwb4oTb2gvObYlKcOGcjhuWYD4UrPAphnTiZyXHXZgJTXM9
JjLA60NmbR1xliek8lWkkIH/YrslQU0U0uekCwoCq2gNmqWN0LlkWnu6C/QuM4x1OtsSot7yW61B
26ZUdf2khKvdWX2h+tkmj3rNFxWk8JZhdUOLGxmnotHq85VAneSeN8PIPJ5OoKq1WsJyNURMU5ab
uHysh2NgcMQlFvda94O5zHghg6Rav7D4LOaE/qDtFQdr5yO0nm9vwuwSHBrmA/p3XcQ/D1jsmDmx
Mg7MfFy/xm81jEZm4l4RtiePg4E4Q95+0VwTY4Ge0Z0efspgRcyBk6257LpM/yFw9zdKZ4SCpCrz
kIUX0eOHFUPno5FBYmiNKrBcpK5HFUnYfSDrsExkxkHfN5zueZG8AljqgfxI6wxTVcIxgFcZFx6i
ukxtaURKn5YURghAEV7aCSojGms2CWBVMw1UEPu9gkyuwwxTSpWKDwdpAtcOwBKmPf9Qz7NoLHgR
/VM2bBoLRZtupeqnMlU4995hFZ9gtN2qlHwjwTUppmFotzur/vFTYiLbcwqZ2aDMxCRmpxNcpv/h
Jozz/nskl5vOPDQ7gsWt+fO7MTYUCvbIIPSMzf7DSyXRCMyEPV4qTjfw1SCv3PdDMtlpIEnaCwZi
bM2ozjgeYQ5HaMjXnKC43X2CJOQWFkgqo0YfNxAHC9m+OMqTQnRFOKD3wOjXVfNQA8DkFhwHrlRX
VVfq16iMv74zYEe7HSkewelKQDB3S6vFuFv95WGHCvUgzqCS7oeKCkGpud201trzy1hAF69Y1Y3H
ou/FjIWTXZEv4A0hA6vrL612Mjq4z6hlbKDA57YCWEL91EIlTsTSgd5Tn54YexhAsAPvE/4XrAQh
jH+pekA80qUhb9sRkHC+cv54s8DqgG0TzeVtX9LGSVONACL3NZoC/4InsxRvTE4acTLnsaFcsvJs
MqtF4wj1aO+PwwieN5E/zY6+EVvaT0J4kMfcWdksijctKZTrFAsFklRiKNZF6MsRvhxhgnL8XkVz
3ZmwytdLa2swPxQWI3WM67QwkoXZjsIT2fRoOuRNeZ5mS/DMfB+5P5oOIuSNq5qCWCUvYB+qUgtR
02dnux7tt0qm7q1ssTkS7XXI0pwOuqVgoYFIKHmrSalZodvPspwH+jC8UFSzqbApcdOzK099YHL6
gUaHiVopJoTJt9noTRr2aeMzGHTcuDDJVhyCvvtcKp5lVSPPkG4UX6xWTXO1Eke8u8R6J+KLdzBW
9apG4uaafbCEwnPDiWIwoSHYLJYJjWB23ppy1aNPvgcq9KZjvej5YPHWUxjae/Uuu0K0bvXim7bZ
AiLlPTfWRgp4KA5yKlvq+1BKUzlLbPKJPqFRnxmvvibAqSJ3Q3mC4WlIKIni4vabqzuoEdggTK2K
GAU6ngzeuD7m9f4jMxWJUdNeYq6LaS51XKMlApQ83pOsopdFKAP65f41fM4Gu4977Iy9Rir9deFp
MuMU1LN10L4LFcuxekrXePKYIUVRNzTkMkpmI5BJ5tgV9NgAjGozHGai0IYWCXIvVXhvwwZXGWM5
GeTKmzx3EUndsOM+v5trBq7HgaBP5aSV5CX/BdCnUs8UCh/G7GTehQbNSl7qRGLM+vSRmkq/m6KU
6rdo0ATtEZ7eVCvaNKUk7bllj8dtgAgC9CCvlYc2ym5RttEi1JYDo4eV1cqVgYI/f69ePH0w9Xm3
9Hz48oG01A2y6RD2paovURX8rT3Zf8B+P0nZ08DbSDOS1ud1x07ZRKWdapwWOflgNgJFrQZEGHIv
hbCe1nEjxNUNkdn3PTYX1ZOX+Rz2RjqYPXn3ZUANDLUqSoXjvthnAcv/ZsHUnzirtY/3Fthuffpn
1+bGATrtUmqtCMG3fYOC43UFx1+oXHqdtepQXw1Auv9c7JmCJdKevOZRgAEpsOuiOgDtgP7z4QhI
6OvV0fRHKQ076FfV/Q5cNGc8Z23fSo2+EfvLqcoNKJxJdZCx8ybccR2YKFVu1AY72zVZl4bNPDu+
o9tJktJuVmZsEAWFkhkP+59G399ltDEwbCyziNibkiWYNIa084yEcI9pem6yxxP5EFLy/aySeYrz
huZopmiVAVRuLXdYr7Z8gzPGk/ZyLoZokj40odm/8tkHF5Nx+kVb6OZ6YDgSLK/BzLBHHHZ1GdFd
atB5rFGSxQrzeQSKNKgT7FHqzjIoRTMMuthXh39OZLzjpGkTSC13obyeOXSIgCuzP7TYov+4gMqI
aQxUmKZzZjgvU+RfCKDu50Nyw1nbiDDQKzQCxmKvNyouFSM+42euv4fW/HEcAHsjCsZXVTdjm1FJ
O9sM9wpqTMqBOcuaK8ppER45Xs23dPI4ZxUdXeaK5dszbFVUfdX0j7vRwQmGH+YQSkdAYLCA6rIe
IF/Qvzs4mUPpWEpT1dBtqsWGcZ+UPhxp3T/7wjvxMagiJC819EMfuJ46wfMwgAOy1vvj7fEzSvK5
0zLa6okAonG4syHbEc8+M4SZ42pku4diGFSN7w2XuQ0cpim2VoSp7lf0bNXSVdhcnrY0ghdkV4FS
Mr2iNbYZ0G/ESs6EVohDpm7VezRqrGKOrnXLS3qn+Bt0Ul84z6AquoiJHaittIqn/VST+RsY271a
120LFJwZRwH3rsp6QkYbfq2EWzqOJdfCML2NVhJ9rs8Ogs2Y6FYZbpJmqP8gpXBj0GFw0fYpikOR
DJCBDUcwrfPtsVKr72lslT4xNq1eAHWbD5/zk/F6ihI8NJpjUA5GqZDFXt79i4htLgejLS+XxFwc
A1JBoKx4sUzjK0cZ/RJDVazFEKJ62cAsz7K1ebIFuOB+4lXxvSZ3mYhw+2y+bPJT1HIgnmMspjnf
d8TiQxek2X9uyGd6c8CGETLh1A+ob0khNdESNu3u14t+5cMyYKYLLDuPw4S6cPjbNUtXzsWNgVMP
9ThEcKP1zAK/wlQLhgWYCiFNgWs0/ZZa1r3Om2veoKc0ml2pptkVUdHOcfWY2qAEBNR3M8kEgovG
ZWJuJ1oB2u2z6V89M0SPKU4rBZh5MDIzf7yprbvG9HHERK2h3S4wBeaTYfB6yAW8xgJFddB92YOq
qU2+kMzVrqPKnd1PIxomUp5X6MikSnWvOJyqUUNxLP7t/06l+CQHtFCJtcJ4iCmK8fF4UBiN9gHM
TXoO/8/qOHANfqTBtVzRWi3b+DhXVqYrpf/P7h14howXw/o4cIMHJDab8XMA+WjejpO46aAOdDxT
8FCUAUFlxFkcs6yBNOumOv4dnEBxvjZDcOFflfg9Dpenf80YuoyMoC61cpHgN2IcEooSx2vWN8lU
Tcr4ZlzBRj4ziJruGJSeVefkdyXuj6iVxWqhjrwendcH+v9bW65YXsej0PwXgqPSmcshwPZYC4QH
L7BafPWUk3gdPfh51YqPSSGsyqKobjOPtOwpFd1wklJq5lUYFk+0m2kzg8Qxx+g0yvtz3p8kmqNn
nd7g9FOstM6cnvc08957a3uryh5bNVsSPHETVp9ihwthJ+1cyxR4f8l+tTvJkBiH5kMXT2IOfX15
Gywt2YuyBnVKJjt0UlzosnCanaWP1haIqfOW+IFhlfsO+tiMg2LzQ+vJ8PfPMd5bUwMEOgQ2WpwF
pqDuCnoRFrzgzCr5RE/X5U13DQTJ6HGcuhW/J9rITipI8XQ9zyJ1wEkbPq6daiB01WXeQNx+H0Rz
ELSSSvxkenQZ1vRauigMoxuPrgkkqXm5YKwEJuaCapx1OTCW4mcZmKjZFh7Y6H8OOw8TebDv4Amf
riYN8dUj8ajQXaE3zZnuH+b6ZEfDONX0Tj2fljJv0rS9gM2p9DiihqLhZQETGnJufnQHXWMWTjKW
x6N2jr8nhWSWDqQE5YHcOGL9uF1D8gbWi32pEuv5kz7vgcrIGON2v0E945ytdw9A+WrmnZLCSqTo
W8ojZUhxkmRkgjZPZg8VSXu/qp/NO2hD/uQ9yKzJMOL1LOEAvexWrhQD3gRwWTBRsY0Qh6ExcS+7
5DBmB14Xkt2vGQG6mgHaT/N2obbkAKDpZXNs+R7V8BY+Mc4Od/+9O0Gq+WperanOOSqMQ4JToWZH
QV4YkwGHZBij0QP8JaEHiY51Ny3rrNw2BkhFJCHm+VOz/LzEjw40MGsD5ZPCvoecHeDOCieGRypV
EJNlqBYVR9dO0HMUjje5SKg6hM7BGmNO4TNuYppuQhz3WzPRCQtu4ylVa8Q45PHR+ujWmKD/QcRS
YodMdHzlEcJeprkjxms111ToawMzxikjcUkD3rRjmM3AZXvYTWyjY0YKL1Qy3mW7fzKFihy7J3G8
00AxbolmBMugPqE0X0re7zmzBdoKSPfaG+BPD6toChlK7ctrgY2oFw8ghFfe0RdbNUrkdx9HWR87
2fXtYw6aLj4GnWqDbZTb+a5WF9YTooLgpygaBsfkk5zsmWG5+waKTZaNBNFRj3LKX5Pa2FsiDmsw
vYw1zy/sinLBg6r+J5f6UL+zDpx2j//jbY+mdivr5oPQXzKovOP4Oscvj+KL5giIEV6PTy1Ws2HM
fPTb/oWSrbsPeJtKvc0E6bvTKdbRiaZF5E/iG3TSYIjhNGwxwtShY7x6Q1UeN59rmOWjXAVs1tf2
zPKbk/IuTtbditHv0zQyfZZiOhPz43yzjHp6OTLwUqXRBHPjc5XzjzQWYccnN5YmgOLkWps6MSlC
1hlKoaGBCcQTA36+HN0e3NFYHH7yQF/FebK/BBdTuX1UFnTgvbZLvLsg9WqSDfNMIkZgEOMKzUs5
2/sM4AG7+d1DK9n1tBPkGnSA5gs46jp64nGDcF+gkw0RSeu4GjLg2Q0V+xTuzMwgTGxJXmg8/+OV
UOm3udGpijfY6XqmrnxNiM/ztXFCtkAZOBzn0HQFywdkdlIrQ1Q/LuctiHj0UzSjBhDjsYedYdyO
IkP6nDo088BbwOOStwhou+SRBvgbkGznjlCM6r6bp/+ZZwDiz8zXypJ0ccvBaPgnjfyoMY7RUlnc
pIn9Y/9gwYGOCM/x0yoE18Y9qbjuDNKqYp/JRdjd1HQfOiIDcaARjowHlk1S62eUdfHOwhSJxcnf
L7so3BPm+3ZDZNsis5bNgyHfl668LOSdZMk62Z7/U6/sXGnrCApOkY4dSM0m3sxM/MzQ0HQsLSs3
4zyZOOkEFB9OvLmOGWN1+4KPAC/0tq4jDY0mBR5AFR01O+ISfsjucSTtJjZH0iUH7f3X43lACYVj
ZPWeewDET2dx1rKgxvSTnRh10znuwdJt7Jgrfw+TbbLO1+kVcscN/cynWRvLfxRNMPM560wTrwXM
0hP3IygiujAcsK83KFmi7VvjxPBCz5MMgAbEF2mqG3yUJxHdpCqztCVkf0w2gujheD0nvmNaXXQB
AV4xj0aB35fVRMFl0db5Bvz+i1+gVmIu963GdrjzfmkYQG4PCesn2K2pw0YER7VhmVYik9xf/1Lo
u1Tylip28IbNtz6RD4lidn1i/W5nBXPmC6qQCx+imS0M8am5iFXyNPQjvZUtPtNRxn1cKd7SGmYn
voeg+ajzgmfe9bNEDqQJJwjfwJcuEAnlfBAwPAyee9+t9bKbXUNZQ6GcuFunM/BPIfjEgub8N0ww
GJKRpZTvblyM45Ai0RAzpHLimmi5q41yOCFUkH3sI9X8C9Mobd2u7nW6uniwnF48LwP7wHadL4dw
gT1ZPe81tAuGV0mPpvoJ/wsyCHc8wrYRr7vS058bB5XI3pqFvPB/ejIZlOrw2Z2W7H4ZGQnKRLEr
dcQas43i4Kh0Ua6WHJId2bZsG3gqqk+ohVal9RQeSVyZChNkl0GCGOIYqto/4PdcCeHzwj4gIfw6
GDjbQZc056GVLzXqvyVMvjL/ovXfxt+a4/ywqnblQSHakNEDC+Du7hrlpw92sPQFiQaceEvWuAxW
Dfej3vYOOr6MC9O0tCSn46JxlRVOuFb2wHmtTGy9KOC/o7dn9P33XuPe+LDk4Fp7vUfnd7hsWaXe
PMXXcRX65F+NONakCNsI7Gf2J5LABmjzrOKUz6GYFZ8RGyLMDvdAAOWHWG8Nk6BgVWX1l0Fy5kpe
Sh3kInn2e50GSrDOSL5L18HzhOMqMjJ2nJNM3jMq0uJt00cFYrPskPQyUmxLOXm3tV8tYwzI79Vb
i1O6fxdGB0Wr/EJ8mqEesRUO+iljvYyOdwXfpngGwbHeAb1tIqPTqeP7VIewHW4gpgFn7eXm48kP
dEkHYkNROiCsEC7Pdjr7F5GSMEUgup81gJ/tgAHp5E8g/0pzkKmDbJGN2L3GMIoK7TgkkwGpoYez
XzfT+AcEiU0Cat2zk7zGhzx4IYQECLd64rSagSlMMz0b5Ij+jUcIe+j65MTlV+fcoQqjJTCVr/Zp
H1ZRNCmBzWDzCLTQ9JnwwBGJgXc5gwuUWH0fXlISyPzIozqqOYwq23yvas3nQBTduJ6cxJTc3k9J
jNB+MlUYMyjeb0H0wzYt7Z/ELHb90NAmIhrYNvsTO/PIG4zfukV1GtY+c5SnI2LY8qmO/nDYVjR3
Mz7BVcgwWIsS6ClJptlOnbfeGF1fhBWeQESipAb9qCUeNhu7P755CAzE0RaFMFUYsot2dXS1afXK
Dn2QUBgYLA5xi0eLlZZ/EMmVmkOjpQuDwWeat25w9/8/czqLmwxk5gNxri9hBNRU/M9QW2cZr+xt
Q8y9F/bEcTqv0AFmG16wDXSzkjShLcjgLoGTDqmhI1gIqFLZC2h3+ueeZzYLgyiVlYo6wGMELbmT
Dhsm5FBFA33l5fsZwmA6SYYXPpLmiya5cPMnGhJn7cZVEDFQ5FniN5W03rEnmeFLas/2TQ+EPFKH
MrU8flTG/cdyJyXgDGwmtvyrcP4zmDisG1NZnd8LAMKdUnFuvd7aPDSLVgZIO3j3sO5ebbpA8No6
uI4+XqqCGWrW7WATaM2sYkmM+HyyDJ3qoQT6ohDLf0t5fw8qXABub+YLURv8RdtnJracVEwOOhQ0
QZ4ykU1DxF6moXY8Aj8tX4Pup5Ftq/henbxIoG15xj8tVEfj1dWMBbZYbCkBsiqTLIxsOsRqJtZw
SKiKlSqWdazFZ+GEJCQcM0dxw+/Fi4hVC4ISMx4igWrY+50Z1bP8LCY5ewHNk++zYelaSrLaJWes
t4RA9tCqOqkbhCpfltsz5yBkqSHWxjfE6IGyuDgZuSvtUT8bPOz/KlkOjxFJD/FCBSqy54LzW6ha
5Kxm4n8TcqsJn3HGUrTlNwQDt48PcnxorXsgcYRL5c9pHKlXHPTU5lT5KPAd0z618iQKMNEZsYMB
D1bxKv10BbRl29Mm1bmMkLGRVPMLuQcOGbho9OozRcsUy/fokxhVxH+hjfAQTHICvFot0eYcvk0G
K8LpIQrRPg0Cg1iEe+jurh4kM++/Zmpwo/6oDGV9OltYZW4UqTs9eXu2c4hpC6X3MxQwZJK47Xh1
etjTMSRTF+kwh5tlYYHUXM3OWrbujlDb/0wo2E2jYk5JiJaEs3S0zXzJoxPfwEiEgpkJFVT7PbuD
Xz1H3AI+Fu5iOviWAW+jT86dplxgSwtiB5ub8Z8C4BnG5irXNkK16fr8uYM6zOoshT5TPxIPFp9l
YwnNTyFNsc8G/uysTKjxtn3N4ns2VFfqD2CiqVyRIdZVIU4vdJeRA464W1vHTFOBpPJ9gDt72OkV
ybuaz3iLF2xVYW/8Zq0PLHXp0Mb0jVBSpuORViZ6udA5VFj8jvlYGuQG8/rr08Z7YUbjhrL0FnpR
8f8Ynx0uZZNFJKX56aMf28FQN4brYjuBYMvT2dNkC43cDD/C0X6DwIDCrIRbbx/xS7vUNajAU3ms
yaqEeXRI9bJVTRVYo3Kdil7snXSGen7+KdL45PFpPX/DcCOq81qN1pNonkcd1HnlitOgnU6+GxZE
ia82sg5uE1jRi1wdEX8+EkmYEgc/JdBMofEVFzvEvBANPz/9fAVWHbOtDU86Z1z7phAw7H24PHvN
/BruALUyyQ7mBATH1nZPkdsA41dfhnBpSWBQaDwVR3Hj4guJNBmdsx9VwtI70qHtw1ZoxEhmmZ/L
DXcUi3nIM4dxGyztd0z+OP6EXwzxtpRIJ5AQp68SfhHldhCz5tSb9tLQxVicM6umeq6EOe9ABNSi
yRz7kZkv2rIR30VQBHPOgtLTY/L/CwXSSLaKZAa6VxoP66olkfc+ZjClC/fYj2ywMo6ORxrC8Xsu
wvt/IkRNvKUGqjZsHPf05aq/3wF6Zgby1of+xYNVZfsgbO0ejHHnUn55Oi+evsg35VFQO4ozVGO6
HN9Vhmz4t7bHRkIZFCE8EeYGQz1wlpnF4sXYEyT8woqrP90GsVVWU6sGzNal9/+1MjGwa0oYyLhC
gyUt4pJ8LAgtieys98SOnm52MjvphQYJgOoTjGo0sKO4eyl992F2ztOyofIktKcYDjoHGspYXxQT
6N5PV/i/5qGrV+MxRTwjEP6lzrkZOv9W3oNd8qyouQZDFTFY/NTu7S4TQeuNy4V0pjet16yYAbb1
+YWOmyWxez3Pll3w/7cci/tH/qGAHKQXUxcTf2zrQKEvg/hlhgzB4ikPBvR3U9CntHYRK8eYRLxi
u7wwr13aVxsFlTdoykrHZjMfwY4xF6ADFSamgSjdDqClpBqQ1x7spT/LPA9/audKBza2EL2gUuxX
5Q4ylL86YXc5w/ON4cXGktOZUPaaiVXJeD8zOeFpJrVaMehQCgPiPtMBJPb29qMbqMyS3LAkEXjU
e6bkJuCQeBSvFAyxO3xJto5Rqn1tkvZ7eA7SSIyFZPnLuseowDpteGacLPmQ6OcYObMpI00zQmbW
O22ysqAda7pmRfAs4w+sPK3jIL5AzttoWmjYaZLETtEsPQHx0LtArHe/ZxKc0C8Kt2mBf06jadZe
T+ofJtMXGAYXXSYCgogyRv7oIvhkpxVD8O8cJoRt6wpjRWgTFd4Q14FbZjDD0380CRRSKZ24S6fm
Yx17JVuq+vNc+vLwDGkKUNJaQunsZpGKtdOCTJseDxari02H0ij/zwxmh+2QNci0i1jOzbri+eXN
vEFiNU5hW8um2WP2lPWdD7SnYXaJOxOS1kOuW5QgTtxmxND9HZKuTNtqvKuOxTKiWKTjlJVGqgeg
RrME8Ns7drI0N0WWo7+0EbT5TOclaRePG9sPluvicgN1/+IUdYRQ0HAZwaQbLoemhP+afPcrlqLf
4YWz48cRlvtNVT+FYYjGuuJxxEhgNAZ+arA5jEdMYqv3GAGBJ1jHT/Hmid5kDIrIq3Brl+03mwZF
/Dt1uMKVDmPqIpEK2mmPgvqkLCDnCn7fvEVALQFR8vLS5NW+gaYJWk5dZNTKcjCKJbxbTTNS7tZy
2n//Dn7Uv1pRlqZ93gq1kNwiLnfZMCbEF6QFruPXuHzmYQhw7LY6Vyio8yN4xlkV912DnfAIDQYZ
PF0hjU0l2zfQ47NtEq9N3w4GZQbVSqjbMUkdol/xMefWa0EhPcGeBVeDH9cqbhIJp7NfEZ8z4fg4
mj8P0jxfq7smFrKS92ihHVJcf512em86TlydO9QMvbwy3N0sdSo/9xM/klbX6Vcqqmd9qThQfjPd
HSwZNoGzHUHzKyIjR/X3QmD8490N3V2VzW81skw97yCa6NkN3nnsGI3xv5EuZzVI/1gqd+b+KLb7
7kyuVQEB+V4jJKzW5MOGXLE6YoTKnFMWe/OT2YBmAw64UNwK8wxM6iE1S1CVy/klvli2KTHMQAHD
AQBsEFH+HV6VDLx0G3mvnDfaPIG0bm4L2XhyTD454TnA3XGHW/WOyJ0PaQsD/u7AYkjdDCwQe40o
ua+CF0zNKazIsn4eVI3P1WNeDgXb+5aHDOO/9aFwL7KMgBKSSo8Qx7fFvX9ufoSiSov4MyXy5Qrp
37gjHmurBi34U6+uGH8ACjfEIPqC8zs5fa+f7zSbS5ywwTNQQ5CiLLr47TScnpjWxn0uLCKFmSWM
8Gny64QqFSHCI17TKkixlbL1kDER/ivlFYIO6A4QDk5bwT9RbOAFpSDYwoRCvsW/1ME4tAEljR09
BqED7VwXHkQC1x64nSzVlmrIimWb2kgSiRxEeLM9ntrgxVVlpPU+/rJg/94yJCCmljClnTz1mvxT
t1DJ0+IavaCi56Mnrh6bovtWMIzfa1lN6iGpcIbFznEs/b8GhB56SxIXNXB1U1Vw7ReIwXYTRnV8
jOUnc0iYNYLtzrPR71c57blBgVSyY2bZGU+U33mOLFsqPS3Ae+hpwmoHY0kv6Ct8Q5M6PIfrGBWq
/zK0Hk7u6jovilmvSWSQuQEvpq/LBklaDO3TpS44qYwKzRxrT/whEqgd5HxaajY+QqWJhEY5jKp0
1yoqH2qg89Tlpz32Utzc8fFjMi0KYQh7PlDS/wFxsAyvY5xmCFOz39pVGpt9XEQnBB2+hEsWI2kG
iV+ID1Cb06PoU/ypukCjZ55pEPn5HSp+l2894E/3vCZebL3NnnTkXHhuMOk029JUQcYTAxyjW/Jc
zMf3zluLgp042POcotcHw2IMdeUk0pTN2Osw11jyaXKhVpX1sXG+hX4EaVKgotC7LYDALUUZpTzc
ssNE4RdfY46xhZjV9IAS7h+yAOfWaYnNUEUb96asuFeuqVLoGjHMTztHT0ih5G2sHqShL3nXx8Ad
dD+DAgLYyZID3OiDd8AaD9N67q+9+2jAJ/eR7D1OSHzvYyh+p5MmZbK+mfB35gvdEWwnymT+c2yi
FB36+IY/fdqza1QNJlTp3i2IJzz3/tGLqm1q7oJE4LbmN3AIl+JLIP/pca+lkJGOC80ZxevmxKUH
0ch+C/bdZTrV7QFP/yjGKu+uIzKs31MyRx15Kzn0WTnifLPXGSim3zyxeL08UZFFntI+zoW477uo
2Frt1S9raaWQpMDNS0KL3zdPv5wX1LdjajuoC38/8PR+uyGu1cnAO20bGCSQWUPSqN8XbjK0gD8c
PxtlgMyvcwGjzxZY/1NLv9J6xSDwCJSASXODhKHscDSEboWS60TM5a9RF8KRK9rszBqTj45imzku
mA4+seXR4x0ygTOkX06yEUhW3zz9gpdYeDtOOeZYavQMztdPP31FtV1RvD/4vuQbJ+KLxqXKIrSs
JjbvwtGNTmr9pdrYXl/sOioPjFDXnXoML66H8fyTdydRJpQkZ6gEZRJJwcGyqwEkUoXyQ8xZ1SCW
qPt0Bf+kZrV1uu2xHSiJE9NeUn6Aoe9FnP7pYu7K1rmdUHFhYsNtDgZ/W3fIQjLkjESN/Do6cYa+
iSl63hsU51k63uCEZ4dvZ59YYV2wt6DyqsgyBE54i/2+5qNLMJVxhcSzOWcb5QISRCCTk+f0CkRV
bxxUhH1HjZLC9LdwNEAdIwP0zTL1akXP3g9FJn53lB8eoTKp7Lnv0+BbleVu2EZd3URQNN2Fz6uY
xHePUwP4iqGxXSne+hAuT0eyJKMQnD8Yr9VKzAoUmGPNCEdv/XghMWcNiiIJpyLxeRotgggpEbA4
RI+T+T1ZXetN45ORMV9VOHFOUtH2/ZiKNmHPZGrq0EUOFtLItdAgyaE78e7FiuTsAqH4jKdrNItb
56T8VxmRzgVMpVDOLRWPMbluYFRRDMbvLl8bklBw9DBUMVGhkYUZNbHzNGMifj0++CSMhVBtCPje
1hbzkcyhW4QyEVSVp8J61aS4GmRvRl2+GU906XWqk+IfiVTIiX2mVHnkLUaz/41vwpxQAbIecp8z
w1zhfSmFYrCCn6eKjbhJfR7b10dlUlchSowaBMGcOTpc3ohBYpGNiKyrK/RMnRfq2elZHou08Bqm
+pJFZNyEZSeLXw6Vw4wi1RXa/ZDba2qisCrN+PgMGPMRavxMHyNC/5fNNlovgCSgbQ1V6WQFQgb6
vORkOTZuYmIxsbd8+Y/ikELhNzR9Mqg+X9joSE9sHADW0FaEddKCLeCtQ4dPFS15BzeR8h199h7d
Gu+Yz086MfHSDe/I9JW8/f6+zJ4ssGl43NioPo6ZJX9rpkPF25t0NqbMan/9hOmvvFBecyvv41W8
MPsSnAYX7hhv9OG1JZmkCmj3wNTJc2Eh681diyne/QHgeklWJHF/QiZSokEidy/b9mDdVPLG+0eK
+mMNfTfC4JYoMZNhFB0bg/KO4thtHXw9dFpe9BMxeu1gbdEziX0e+3r13kA8YOXcBPXTj368dtA+
JIhduOXNWR6CYRoXnLDbmyAhmp4PaeHUzgogOaIJtlvD/ynrpmHMaFsgsZivzWWtpFhCcw+SMLCu
7EuQftww2rHYtix4z+/9JHfj0DKJ9dz/7Ow684nCNFQFiXrBKtkXlsuBps8l+g8HAdOeo3GbPdvc
/1RnhI3GkDpnSHas0W4IMFk4jxjaZ72VkD4KAHylmn5AfzRq0HOMcJzqsg0QI7UMi8MSbD9TYOt4
ztQAhdrsGSRfsTS2Y7MOWzOo2winx1QoaamJCBmxb0gmkp5iFacyMvDDqgxKUD+z/fBThrHSDs/F
C/fLBzt6s74Kn9cxM0Vc+W7vHcNv//ZnqvMPvl2wFaXsuRcWtr5AlaRfxd2cQ6suD5Uz/ttpH+K8
v0lknh2xzv34WDAcfZEX3lQXOi6d6HZbG7jYaARqb6ZL0DgFONCy7m3hnIg4ZtjXs4f9qmGvKlGI
I3U21oHktlTdGPaxQpQFPyHWG6B14IRBlfyq32zDdnYNe3l1n7WjqTQjTaKz+b2GA4F8nOCEFVTc
fzqrOZ3arvm5wrSfy6+N5OrZkpb/I0mkhlHcGV/wwFBDyfosnL/xL8fr4gcEK3GI/n+1kOKM+IoA
OsxS1gtHVEDfCUHweHjBCx+qTTiiD1m/salFNutUBIbKO4Qpa3oYK3S5hLIenLo6A2j3Fg380AYW
FkZdZ8AlanlT1zrunm50TiVR4CIk+RTB97rYFoVDDR6HJVNtgsh76j9jUP1S5d7Zx9UdQiqJVG2+
JeFbgLTSfElVsb3S0NYFh360OBe6rUF06hK9YKqJ2+GOG1MnUMIfsD1lFwOz++IDk+v841ydn9/j
RFMSWCteZ/sJXRcOSFZM+m7PA87iMhC7XIxikzFvi7QNQGfX2nqrJIFszdR93fRBe8oqsVecPD+S
sU5KgX+HpXfZtslDsbCtxpWMPYjLwLSwup6jh9kFRyxpAIncwJLN/9kmnECJ0O93WtQ5xqZJ+fGd
hjl+3gjtLk8UZp9HCpNYJmvZVq2m9n+sKFoHQXKHvugURqpHlXU3oTdzc18KDYrIoNHryA0xNr5H
2mXpPzJK7Z/uWf4ZIgRfI6qNpxiVJgQUVduzaD/RnQjXzdQacKs9ukpjMaGUPbm2qFLCe9+zLp5o
4x8gbUq2CEAGQC3wgMUjRou+EQ4Icc0pAl38o8p5vY6OGc7APXT6HIHu1bJ8lfCOORqdqGZ8Zqbb
sVzEoPNYTIhYaDC3VDPdWu2RloCogOgnLomkrk4m6uAHz6fipq+nG0PXHVju5xOR6zjNhBIlRw0g
lPv3S9HTgTcZiRygDVqN9C58lbSGCb5WyNpmm4wNoV4U8D8/cC61axiVZijlkiUUHV8P+zz6UHEQ
Kv3mkM3xX7dAEFkvr3OGntb3rRRFiATcAycJlY7ydEW6e2Ab7x509SvoKoExcPbwNsxeLs/sm95T
eRbUidwPGMAQHQiHPN1ifTPgllSi/9rTIdd/mtxcFw7QBtpSPQ/WEYGwvx3QX1sk2JhYYr88qnvw
Li0IyHljdl3zDmbPZMT8QRcamwItkncJbvVweGttd9QApD/Oqb/1fTABsiRQQQREg/rkf6oeIbX+
ggm3wyf+s5JFtx3tN1nmtfUTsUE4dAN32wLjEsvZDlnDTAxGVp4a5jgbWftpO7wWfouwIAsnMab/
8bpdJsJnmtS5iaHg3EV70uvCiXRY13yd11t9ko7aPwf/jFZRufxiyhq3TkuxJp0aCToCPjsbpoaf
+oeydTnjiFP0fQW2yQGUeoFkwPd3itX56EhwcWA2m3YQaD22ZTAoBk3OrcN1TnEFdsAZO/W8qScc
DCIG61oalm2ZvX+rYh6uQ0ehBv7MjCVsjMklEngaSvVeDsd+qg+8accFY21B1CuMuL5dnGJgP/jC
ni+0OPXSzWegzDF/7S7XEBw/fT4/GIugaehcfJZ+e/ew8plydGg4UTUFzi4COgLoJkYHkbLoXERh
YBT9yNKXJp4YYWpQREgTE5OLHisb5tMS03htxAOrO3I5GmrnjWgMdsyPXszd4At6FoRw9ptBWg6e
SPZBfmVVhm5BcvxnS7wbGiFUDo2mt6eY58Oxgz5QebxUeZ/T4RNhfsukr4bDlaNVsLXZcxrf2BTX
vSCxBvTGR8b0ZNdzFkH9fvpuvWRNsptdS98ngPsRzvjiosnglt05zvagzbNN26901QknP9ov0sIb
6TGkPaThbjDcnz2cumkDAVebnn/wOIenJoIA1+AdPJwFmrspJf8VPq7ceQ1Zt9ambUCjTD9frK5o
uFLes6YoBOOj2Q1Q8eCSN0FMF28gDywWh/5+kiYGyPdjyzyLWpxewE5liRVtgVkgKiSw52vjmJKm
ltmsB6+iBScDTgsVQ+lBkSKFtV5qd2UAcNUqUoNd8f2QQ2FuKZwWONWLNbIbHwr1KVcxYftQ170t
uzGOCspXtONKXo9Iev5Q3bjw3ZSZc1vxsNt1Xfo2lyl9Hi166a22dXa9MYNhvu8MeSMM2lNyURFK
+YUHQY31LLuUVaqCQhkXMVy3/rgqnaPLZmDvnCO5Zqtdw2h+gc6iGNlC9K62xKuJyGKA0Z850nzh
bJpR+lZeyX++0exTE83upNolt0a0nCcNxSnMKsJj44KBaSqqMSyzG3hNJkNfTqoFs37BDGaBnZBV
OBmY0wPvK1wbvl/O8OTGtJr4xpv5U/Jf985Rin1Ct83/IkjAGVvK35u3C6BpcBfhybWQlyJPr95k
MfnTVCHVXFOcRnzqPRDHLuV6S1uvgOnqCAihAcbgD4P4T+miwWf/2Rgb0UntsvqsR/6vqNXpzuA2
LlbjuBOuyvqll4mPp5mF802VaRpaTYG7NfiLpilifQyd/PsL2qvbNNFmOtCq1VzPi5nZMmwbDwif
MEtX1pysl8YGKd+eEYTEfscQCD8SjR9rHWUBQaM0RLcFPL24Y35zeYTc9SeRgejb3xISc2q3zFhr
FWATbGIJLDnXV5QobRaPxkrRYAHQN4oHT1+ewu9BEt1YeOvt//OPJ796xuYmGldRycDj+eyRkMpa
PcK4SeX43Ucr6igCmOHCv2aUaZNv1/nL9BtyYJGvFW0vb5qeYVmbQPqPkrp9XIQ46lkrB5wO+gLy
wURoF2+AlrPoLe/4JHiuGalvzU6PJCXE5kEg6aWs+y2TXZQWe5N5tjF4aq4sUsrRu7u6zV9u9niu
2s1N14wkejAQgz2+FDohWczKAxOfo1ndTrR0qyb/6m8wYZ9AIP7vBp1nB7+AbPmHZs7dZ5SjyPRU
aLr8jvjlRwmMoxceph2ph2taOVZgwvXHf/JMXuKPsdglg7+Da1asEqz/SZiZ6XYux4NrhHDn/mEq
9YaTWhAul6SsUnWSDIig2pKoN0DuXCtngTdbrRleHDw/s0/tTXqphDGQGk8t0GzGGTmwnssKUXQJ
7+YMIN//NrdW2XxfyANcK7SGEs9CCqBEYzR4W8XhGIHxnMq1s3FVdQ0AVAGp3aIWQ9TKC9bF/OiP
sZHs93QjlxqpQVPutEeEnJ3Xbke+B1PgjOHgxx0FCKK1wAxndbka9cvny1BD9IXV+/cbTHoSOVBh
/I0aMZm1WAsmysnYbRxpi5/imMZ68+Pq073OoUJs9UlT3U69TQAnbJddiZCP7Rqx5+gNtB3C/o17
dyNIHNUXoJETmCLCE5ZPxesZeGVp/FCsAlDuKkyhsOteyOPxzcWeD436spPFpLRquNqy+MafdSL1
WGUUdYHjPkgYw3zud6NFMHBlpU2GNxO0QpxLzAVjmexoePXTC4YacYH1J6qSSZy0xvokBaCucsyj
liJ0APxhe+jTnbBVqGkWbhQDfDpl/UwovRUa8MtmXXv8JwbmMytdvmEQFvPepwwZMh1Reaiw/JUS
6pGrFAi6lJryFq+FCrXYt+Un4GNsbEdmINYwma37sMPIEdkLcakpezgkwDD0C9BtZBaOLxrr8Lj0
V6yW6aI4K4PsMr1lPpwm88BfDv5247q/ig9HHmhrsDsA80kKDdf1xTrfyb1b1w6b+Wzdeo/Hwxnp
/0+avPByWdl+p+wu//czAf7yLGz+pkRhoH0/SAlWDeqH8E5JITKooei+Dq2DxLre4XPemrbamAt+
QfW1fF+TtNWLFCwXszkqije5/KHbs9W+XFq5Qg2VEoDe7mgsFkeXFqll352KWW84PzvMXWU+BapT
VcYhhCi6PRmDU03fUI0qorpl7JUr2T3QHf8pybryZUl45Zl16hnpmsJfOE/BD4KJs4XyGCl65zBp
ufQyImuDl+RWJWNqNk1mLmE+Ek7bSRFP+098dEkX60reD/pw4fm2r0hZQU9UK2IG7f/bhY1EO1KB
d6onrZUxvRMQQVCf9mUkdY9KFFd5EpPr1Oi5ruPVWb0ZP8ZYCIqwAHtqIKx6jh9fc+NhNUOBm3TG
0TvOyfdD4I2SP9+ytxjIqO/1umftvhz8vg0yBZsVpVk9lG1vMpri4jVALBaq4a7YWELug5VoTVfz
QdBmzycRxxYNBXveBn1Cn97FQs6sR1me79IGNiL0wMbez/hRY7kHpGX8qbO2R27QciKMsqoFMKFM
yu++CqrjqJGbmkCH9L6a5krI0ylIV1j2rfBbwtpyy8r6bjiKF9Z/r6bN82fQy2uJ1zFIrgXmdV64
nUNbPCF8FMv4hpO1/LXKehUZZ4aHIZHjA27yjmdXPLtR5Qcl0r2ovEoX3NfeBrt5/nKwhYVAEPz+
gYYEW3sxtJhvTPGSxkaDKh/QTOOnCmylMeTxyu/9TiF/YBMkDB6WMz+iwSLagMGIQJwp5X5lt8cL
BAjWkiGmildrBFin0oDKJBP4+f9nshzyuDVEHymDpZKVuxVQzd9VeiBwKZgz8TVKdD0sRVdwHwMe
BqGAFMfIpQg9qWQXVAJd0LtN65mcGJ9eHEeHMe3vucKhCI8ZhOXubcIm0fXNrkOW+K4nEMYrNCBr
Tx6CGPOoyj6umaj/KapRvpUYUMbHoInXU/j3hcA0k69YhvRGEG0QPtOB+AQiFS/6Dnws70/DGIcM
WI7aksE0vcf+BDlsdSA1jE9olpJFS5a/mB2KSsH0WBPSMr+PFxkFr/lmARsW8Q5yFS9RYJjk5kPr
IClYG+gbIG853DZQXsgSU7308IhnIMuD/y+uxQA7ug6tWareEGBjrUVk4NF7eGG7gb9opjhm19rG
LpQqm5hQqliUSAfq9ClpBDTHcTW92dyHy+e/CIyo1tA+CV6Z5niN6IzDagrJvf0L3AjuIMnrubE9
3w3pFvuNclqHUGbaNTdytBcuZvsT45ae+2qcNQ6nfFyqMsAkfUGWfNzDRP6SjarmQNHAWBdT05IG
bhz/nJ6n+1PfBQYjsls5vhedWrGjxclcXcsN8Zvyp5gHeLZopBwps0H/O6lpcRSSV3Z0YD/WyUXm
EKk1tPmc4WfRXsQxHdKAGZDSX9E6T4Yz+n46s1MEnW5pVi0EMVjX0N2It8yG7wnC6Hyz7UVv7g4L
zgYo6f3n5zy1aSSVTMJpenIGa4/+RefMwAEZQeHAtr8I5wY7dNnbQM6D6F2HfTcjikDPmsrZqYHQ
KiJ5VZJHu04j8MHchLAQOORRbormGNhyB8ZuIZvHPkVaeq/M/2XcKLsu53+0RRcQ7ZlJpVbXxmy0
PVIKdIbHGLa73fmnclkWd+6rTKtA1FoNbI0D3yAI45Jk4LR5Wd3b+/1ZsYE5YkGP4ri7AdAMikH9
EYaEDOHvYOf0li7zdz+E+oeuzgcunOU1x/tPrwQHJKm3C61FntldS6wuWN41lFdoJMdF65gdkKB5
ZNruQ/rRWnFeNPFCTD/mpAo/fzjeL0neqzJH5SgQtHyT5Iu1hN2UKvs+az+8mnJDz+sP0ytR3v8O
CmwIKi8xvYLw+GFnN7pNc262NgLyUDIP6qqtFDBhM7bx+GCiq3APS4DcgS9YTGh76hn310Izu93I
Ttx5WwZzd8RPXUZLdP5nGASGqU0OLCQVH/7pQaq21pBHmRwi4Ml1Sr3VnC0DGSxJTELZoQ6cfvcq
Ewv2Pykb0DaJpS8/jAD2X2F4pfEF00FlZjW0wDFON0PZsU+mqYzkTbApWXuzGKvrj6nwLXzSbLTT
XfO2dPoMHxh+CMnGo4DF6u1rCSHGHQ30OyT0KqDM8Q2SwZU1tp0TPuoA/qezrzldYNt0tdzTYmvA
WUg9YaK+zjABaP4vHMaY7xbMGJVksrtvWbSm3DejfGvmzILQ7iM4vOj5Gdv952olQaUe4MM/lSvn
uEB5avVcNlXZnNwp10rqx+uYMJtThsjALvjwn9oawEEaMlQS839jsx+urMvgIQpO+o7UxSQUwZ/s
4Kg9pt4v94XxxndKNd7W9PAMcF94TrnJ8ZOkagzFD1lTMl7DZgFyjM1dycUfwhUVvhyxsSN7kmYU
9f9Z1bvkePc56y6dBWqb/5833hDjU8ORcFDFv5/wPUxDln0A3o7RD//26uRdOKBbfv6sweJHzNip
dWiLhyGIT/c1tjQ/cuKatipsUJ4zXRaOsk3eA17dBSSMDEMOkkaXmxTtT4TCLKx0eCj+ZMUo3Lrg
QfKbYCy54zQ3QYiM28Jiy6H740S5hncWzBGi6kZERS4F/rTNtNlFzHJSfb7bcaSjz3R2htLqKnUb
WxIAMHlX7ptKN9GOshTcjd+BZYzMMK91vUNOrfd5vdMwJ2vnCKZiI0XjgnF3/OPq/5z9bpyZGrAT
eLMIIJzoposBAgHGu89pZSmq3dMWAnHb/pKw2+azwCyUqfVs4mH81Lnyec7hWCFlCvbnFczWJGHq
QJS89Pst37JgnkEtpIr50vqZ9lZZJAxyN9ksgrXaXgFrZvL0XHePedEop03K8HgUsZzcoUOcOl8j
zVkh81YNcdU8NfxalAecqbwJLk9hqqxK24ndOyD/VtSpmWMlhrDn//IP21UmILlJD3D2ZY56d8UY
ROiz9SK5SJ65spLt4qxMh63xIzf6Hs8Mc8JXOidpEKzVeWKeIJeayWqiMNeulW1nbt0nyahqegcV
icshNQdQI9zopGkDkeaiwIagALZAV33I4+rf53g3gX1WL8puRMXZfieaPXq5ZLpHdcXjIqLcPcwx
POB2xCEzuUfbbw7EHu7UoIT+gDmcgN2jWPH9m2jU4BzdMHo1mWtfeQtggevbPu6R1I4siOYbgQ+m
ukYkQAaajc+z3cLixFWgV9f2+gosMgjSNeM+zicKjD/BKBqeSxbzr821GLWBL1r+aryPWMGqpNWU
0uYqImZf6MBSopbipdcHxxMbtBErApCT/EB5PEjrVI8aTwHD7FbdRxeSBWSlCFD54b9kDSO+8hSJ
F6OzfDVuEav+Hi8B/iVkR3f4QRAElBI7XR6koURB9CSJlWyDE54BI34ZhcrOmeIt062jqGD+mbB/
x63FxpdHJH2MUVIIAx004h4mSUr/kj/ARKc54F7fnp5mEQU5e3R8fyGN7FIWDeikyG/aeSu0FubF
mmoAHfUG1F93Xv8WIoozuNhAlowelQWkZfug60XeFPyQUkIQgQvSOIOeqQfZomXKzU6SajDinYgH
GssjI70QcRxkZ78CDpr/TKNw58TBN9yT958r5lguKTW2rlDfioYmDUJ5Gvb1uwRVG7NAolT7jiL3
z6VP5Ptu3aqp3qhqDOBO3N+HovKhdL5eY1kEDCrfrVOd9Z1bp3hLNs5MnUI2ZJg3+4fwXo9eHu6r
fbJ2/85XkZ+5Z7a03du9fJ3p8Odtd/RMvplEzjrLh6BD/KWwQwdFnRucV+C+PQSLVgdLswjwZQrB
fXPAsSYWySfYhVCgKpbGV9mvn469rPUjbPD5ZzOgB6b7rd+F0zbPcjo0PfSMxwInzB3gLTvKBBe0
SA2U8AO0kmOLKR0v2wW1BlgWCX3AcYl57SjEj2OETDhVSjjZgM2fOH78fzQBuESUu71NSdIT2O1V
E1vEtIjqAlkPOUV6DiWDRs8G+8Sw5zVG5aJXVqNVZxWdNkmyYdfOv/iho+SUTjrSG0lcXvtkz9hH
Pzvy18h7XaNf2fQZxJNZ98E41gmm5kZpLpyZA4+ZxvOptyz6lMLzBanSOufi1daDlnXdNljMeTnN
wMkKk4hhKA7PXYDmeld5qpGdpGfOcJpzGr8qjDQ/X8J0r8DnDrbnbw6l3YbWRyIBbpdxbLpasR4Z
pf89uASSAJy3yiAlbowlPgq/kA8pyHw2UyZgJGirV6Mm6VwvgsHxkuPNDMzn6dOv7SCERyr0dlgm
BoWOXRdmbfvQ3HQ4bWGWIAz/5uxtPtFzuNSVuD9zwHdb/+hPf9H5nDLQKydpyzsnV5U4k2E5pH5U
dYYQlSDeCs5RIHBFTE4If72e+tqRqGkRQ2RP+nG1y4BkJUNkRJbnb2f+yXUcP7SntFiemFBsSzH8
A5ARFiIYhFbikYX1NPlGgwnmTpvIbzS4fRIwjSPy0inbBe6wr2LJhE17/y9GivWrESe+5epu7bEj
XrMl/otkbB1YJ7heLtTyozDf9jqDQmj9jMc255zi6dX6B+G+wNQD/0T229zJDtgD80BFZLqScoZz
avfmhYo+fhBqqK+aoSGCst/71MboyvWr0tQw+FyuAANp9IWiqLXr5h3VBIwp/IVZ/Fg95hijeUKU
LDjO7Wpf7K+lcCW+oqKt3d0OchXKqMNNTIQV8U9p1+sMQbSH85/kLTBXge9pF4VOGDM2nnRYfEtU
exa64OnRdpgzZJKxGXU3u6UfPLq/kiLudaYiq9jzuUwWyw1e37NnkF6a+U3OlhuR+xCINjZGIWb2
oldoKxCHQrSvgz5XSGHuLpmoeLcheQY3Inw8cn9rnGc4HUqjs5hMGty91IYa6lAPK5PbDe/e7t2O
P0kA3oF0cjSUOBF7NOzgqjBIlKV4ZC/+zI/q3+6hR789AEP5LYAIcts8q4JhwCH4QDT8lQti4wHS
5vAFu4K5xzrlJYZsixWsmfFsRBzHzZLM7WMGLjEjCDX6pDTvPgy4PiHCENQODBBfbAWHE1iY+Bdu
MlldscOtL0f+UTF6EUAQDBFX1ywJXMjG5C7av2O5MDnUi68ULkut4YJm4sunSCEGWyL/BDISB2o+
EatTcd0auXoC0ZNNx0fjsAYD+bvJcgedeySfwkY/VWR6BFUlR50cXcof5j2DdU+4caCHTS7OwGGD
Op/MBa75F9rg59QI36FWCzO0ZX2Q7cpI0ctTQhQmrd9STOIcB7d0FYZq2d2xM8+dK6px5jpYCB9d
XFWFCuxyLrmvFMlKgM9ZI3zTYDiiVf3PJ8KOTXGa60NzEAixaHvul23kOVch6FzVOX+hWqvf//5A
O0+e4q7quJZ427n5YuDZKCokhOjb2VQ0Sp/1Myc9WnHXoLwjTThk4u6IsJuJAhEZtUEtBhFEAVfI
copLW0RZ2ybzME9+C3eX/aO7/gt8avrngyD/no+Eey4ZAMGO4t//GnhbJLgmrSy2gOKqQEy5OAZv
5IVYrbkHCpY5Q3areCE99T7XpL/IvNZQ2NobzvhOTSWHg9XxxqLRlm7Mk5ZkYSeIrnW1mQV+GLL2
drq7/SH3DhWrQqFHQa7OtrUkSf9cwU38RfuWHGGdZ6z5lxOdeYuzC5Vh9hS4HUWThoQFvnxVbY5n
PaKiN16OnlVJtDC/XFPZH+S2Ty8BHjMdasMkyWIDRQJxpIBMKaXb9wvZu190XuQRGeyQHVwN5H3P
nLA1WawCz5ffTEICRdNvhkGDk47/3a6kdsmKiWUo5gyUj50oBubxEH4ZKN0/hcoZFFL78e+D9Lq3
lFc5uTgkrRNglZyogtpAuA1xM5p7qWcmmM2G18HNdkJ+cNEuHdBVeMmDh5HI6jrtkJFcBtXBDc2p
JVdxbaDy/D7SFDZB/E6FnGlKMaewG3sa2WOUWoc7+Ws0muRhlxO0GlaKZ9lBS64NNO4AvlT4Yh7J
O7ounGy0oEsLj9qttYMI/jB19MH4Ce3mqd2+/tBU+igwIdaK3JDnkCj3eJRmMKH9lCCADnK55KuW
Aoo/YX5O2DQDafa1Ey0i/4Z0N6PqSO0w4sX+kNXrdJmrUi5j7zPl1QdSPA+bweQoMGytu2g0l257
O5MKWV6BPYX+b58IBmtBV/hESvSzqhea7ewXaiD/XBYsmW2aE/CcQsCOD067UI5FsgSXQzXygyBf
xwHpe7WIO79NiJ99lbI8dmhLM5OL7xf/Vc4+7pdqZwZxdkKK3CrvH1imef+O//VTKv/893eG1MvY
zYyiTWT7U5FifQrPkoq0AXyxOu60c6N5qzYdUkCmVZPSCJfXjx82TMthZk1ijXqFfw4fP9hIpck/
AChWn5XmmFBdFVTRC+QmZzFBk8dXL5dO5LOi8r5u5nqkwKLJsebm/MIyFyQ97e7pUlEzJoW7hhid
3QlWucgJZwpw0iPapu4GlyUi3NzHL3hCKcxtMJ/KkhmRRQbQMMO+jHR8+76b82GqejlAyXcRCdsZ
7mA7luR8H4yXQn8UVFS+/hU2NfMzXT50BFKqIAMWgOighYakB7CAK3ldhvLhR2crQ23/q7njDTon
7DgDtsVYWpFnQmrADbTbseEkfy3X08qxApy9WFtU2+9Ri1qJM6IJ2DPkwuzcq2trghfhoUb7goMC
ilgBzyPczgCw6GK9Fc9xvYjLD2Cx2NE5TWaDLh/mBw9pGKvWo3meTjBC6EUgag8TH+vHJ1sqv0hE
0yCz9z/GdNUymWfXHeHG50lWjRpxTY30lzZwtf53fvLTXS7zAqXBMjal72BNA1dIT2EWD0NDi52J
wEjXgYLkZY02Z159RlIVobXuo13t8D8vBURl6GQryIkNnTudy/+/E8BHFMF4Hmgzv+wgvD74+hxa
J5t1x+75uMZINoxA1/F/azlYWYplOVp5J2y5ZdTOd617Yc13D5X6JU/3oTNYXb5X0hyrcSl/JgLT
7GkExh2DpzzKVzO6OPg5fwtJ+k4QaoeStpfYPclwA83OPvHr7R4kxrzZZ8l+Fe352C65FBd92mXa
k9U0A6UYcLTLnSnhTFvCoaLL1MQE560IaHTsmPBGCMjHRYhG/awHp+0oxvBdIXhYBj7DdPFj7PCG
Gh1X1BKQtjpZvz/EqNacm0HIR8ypo2mksyt6xCVBuh/CWe8uVSF9/r0IHSSm3q9i4V2HSS/BiccF
J1LisVoargxVEQg1Zbuk7yNjuMjSUtKn8vRjmQHbrZKr0ZsWiE1zvJuIeJUXJoC9Id1va2SzjayF
QaSWsDCy/zsn8wWuX4fvVeOrHMdCcW0UzFUIjZw2D+sbQHus+wkdhSyI+5oqLGsaESIBT8owh6nL
QyC8DFmm9psBi8S+Lczw8md9hN3LS/oHiXfkkF/rfJMtipSNdCIpF8LaEy2N9eMtqaFNYplIESQy
HIsGqg1ShjSIGP7fqkPd3O50rd0bVwjyxbF8dUGkG2sn9zNa4NVfaZT+R4fQUOEyKywh+AA2bQbz
idwKtGYKtedZ2feAphUn4V7n8a4Ju7yuqEWbcxEQ84mVX8TF+FyQzSIxThesS3xRbv2/D72oRVld
H5qqSvkYjdrWQIICHhGtkGlXux6sa2TT3qVELgo0b/4uEKS8L/Zwi8H/vw5bY7YI1o/30cU8pNpx
PyFiArSv0dNxQXpZroW3XX/0bbrFLuUAZCej/0Q/Vlh6i+uBArhFHARlNwixfQ49EKWx3+EY54yy
Poia/OzsXizLt4RKyTqE3iHzc/pVNMrPtkvPI6fWR8CqGKFLm0knjgk0ajhnAZkaIzUtMC8qX3fV
T/gevx++RKxGWCNo5MgbX0SPp92qzd4p1MiV6NTrMTPsOsxfq2if0x9c2QlUVY6FH5Up2spELvak
97NbXAw8MIXtkzSuxTXwiRBWZhW19VVA+EzUNK2bx2aCnPjnqJL8+FfA0vvJ3AxE4Sb5JoMhhRhw
SI4V4oRpqdr3gJIvtONls4F5PpJZfXy5oVTl2N8W3UOELotCa3TpP3nPj7KRQDte7EIRpcVxkgrZ
y7ee8nNk4pOSwcA7ZP9AW+Vw4YR+LCpOUc/aLMqVjAxJO1Z+wS8/eJmZ8JY+M1uEW0foxqAJEaBK
0wTwPhEgKRFoDj9QaMTbkzF92NbuLCuRTMEtIzzleMJH11RgqSN2vHoG7dOapBwQYiXN7uFkaz1C
3H1KT8ar/kFdQW/D4L6koMGWA0zzkqlRjLod8B7VTl+yQfPjth2AAyqCV6is7HRbjiMVbZ3TguUO
CCrKMKlxZPPvAPxF+ziVTUSwIcEoI2zDzNtSRLK1HY1kVgkR4Wjvgcug0yiLY43QGRJEet40h2vH
aSRmZ1ksLgMrkKSgiobwf6/vyrib/r7H70NfhWhTLuSwnEV9eRRLmtPHvnR3GeqbUI9vZnaLo+Zl
IxLFJvhCDpJ0FJXFHIwVGo1WL/Y8sd5I5M5COSalqaLLZBhcsjM+Y/HF7KHDga44kJTgyL1KoNI9
cMw2NcxR4ROdTDdlk6dIp3XzTGMl9fJ4NUlzGttwNUMnk3wTs6rs7UZ4snqnF/1xrdtHHw/mR/K+
uhn3OqW+l+cURQfU6oYcizXrin6wrkrmq5VX3EGAJFzmoGxq5Ra/jKTyFdKLs3ny8MPlKIw7J25W
Uz8EmKjZk2wEi9sJsVXNlWvYrN0bjRoeDx84jWOOzBOSL5fB5mP1ZTMD08YWGNwdFerQaHc9JKfb
6Cmms4KQ72ePg2maiC/UR5F3XQwmRTyHL+QbEmpE8pk6TUHsxK2d11br34D0IEsv7jUiDbMaEXeN
K0Z4ipEZUkkoy6WBH92kthHaKrE92x/tgITNQaDh5u5ReUJmGU0sKPsZNx6cWiFN/XjGKU+VGbUj
sy7wfxK+9wqGoJsbL7IvENk6k3bmvLJCgBY0eX8FjBJt+lOBOtbZO50XMnwM789+hjDEoz0Dupfp
o8QILkGGkIMWFAFs8DAhaZV+26bNqSy9UkY0SJ5ZAshCQCOJ4/tbphCjwyBpMdr4pLPWXYJPp2ZO
fOzEwGMf9BnxtLVyIDgmkQ5nylQs/PBF5FxqVBxQ/NXJFjzHLGVy9G/Q1vdGj58EYQIjyDQk9neG
VQMpXEBZogxh9Vq8iC4WZAxR37YzTYR9QhInso9vfqx3GOxJC7dvtPbD3oErC/0hWUWk1aF9z4Af
Iz9ZV57uPf/vPxLhhxRB47NEOK9dh/O/rhrausQxflfVqzbud0hzRnaFNJiutU6ngs6nqkPekYte
gnM9rFl70FxFv16OGpoj5DtDmrKAI6p75qakaYB689S+tnlVUiAuelzNR7J1AfJF10A2uVELt8wo
jt8iOmKfKxmKPYIkHMoL6cj3joWL+Y7O9hvGUmY4XrLRhJ1wvhNtzUlaInJudTOmIXlqoxKzmmfb
ChUmiYnGRjhDuGz1dx7le9dTJslY+baaYWKQ7uCqOsZVTVmot/r2Myskw2XEsBxF8i4zyVR0qv7i
fMs4lOl/mwTLfGEoMKXdEbD1fsRb050wW/02IVkdGdMRnA6f4uTXmJwk68KmQUyyx6zDF0KW0w3d
Y/OBuVXaHCU0vvhBR9gRnE7pGYzigEo7Yo1FjKaVnhKTdHiHBVkUUvpRp+iQhoYBvsLRJVvSdxcF
AHVWKDbjdauNHfst4Wecg6uEgXEyiiAEJWILYnKpE8mc7hGfbD2/ZWxFJOFYBTjYXvvSSDUIR1+h
ClaXcfxOHcxhpmGsVOzKmJly43OMBclzmmmVc6gw/GLQKzGNK1yYKDcCNZaJNsTSTzoey3vbFrNS
wbN6sf2xXZm0c7GKCGYKLn+61cSnuX6Nl+GS8KveY7/qolOD7Ah9gPJkUV6xzBJJLwmPF9NK+QYs
KxysiIRX1NmrOC34cSG3c1b+0bmiXXB/JZWljkjS+OH0x/BJ/xC4QhXVYpdLZd0hRIAvfEg7TP8J
Rd/DwlzvVymqhdDP1cYmP9nPX8DRBIK4sUR72kjMZnhu7gI1GqFTTU7CznyKeHf44vhpMGE9xtIc
13O7R+heQV/zLro84FnOFih362VvKWQsGOWdchML4AC7NLgFvWiURO9/a0oCNIzAFxxk9J/9IhP1
UQVMDqvR/dEDsOVUw85Qs6giMGPKgEKqRgP0B4JmBB/8MZ0N8qf6rV0MZfHn8vyHACzFHY8GJHrT
oxCgLAZkmNNv2aXROFvYyYn1Fyc6KZ2UQJYJiEE7J8/NVpzG3wBYK6GJ6KxwYicehQQXaYTNBxwD
PB6U22c7bOqtF7phR/BQeuNP5zfzXHVcmWklx44g8aF6BhZ5XULnX+jbDHE7forlViOE2uQlQJra
+kt3S+m6SrrfugliERW6U9APzNuZ1qwpgaxMs74OmuLbG1ETid52dFRMciTRMF2xHBkV70PW44ZS
9BLr6pDtwgPzHCLK+3/TgmVcqljB2cg0qLEhZcZGDZg9bwUUQFrewc8QhQzJ7UZvNQv+nEbAt/1J
khurOAwnrtkxme5OF7Wf/xce08ttqOhEeUPXD+TG4ktnz3SKoJmzrJ+vQGKWiMkHprhMpHg5AEEq
uDKiU+eyz/+4CfPASzx4Npcv35cO2q55zsF/VSP987UYy6aq9XjFl3A8gFu/AKzKJqUvsjLZwVOE
6vxTHqpGdf+hvm86R/QLbJNV/DdKlOoZDCylbcwzTdIE2GQAkOvlsHq7te5o1wvjYw44JNuOh2hN
+boGTmV5DW6WI6bW4JdaPCplfAEEynNIow1QKSI9gIXCTUTMIOWZZnwlVPKyLyEkzd1ycOhdxGOS
MveQlHzZj4MDCxFM76AWJD8psyhmCRzDh5wWLC8rWjF1qn2+KxJzDfGTi7Oa2fXe8Zz8yNsqsBQC
5PgUX+wSkEt8Ic2Henz+i0VCsj+lMmhnPaQMgU7HnTsj5hKpbtcqJYgqoQiTRKHoPBfR0zvgTzTb
TAHMKKLKgyQ+FVf+jrJ5k1TYjPMuMRCE1FgXFvu/XRg8kTJEpywDO7vbt9xEKzN59rTyEIH8gY+9
wz05nbwQXDnqP7+0TKmnfq7iW64ieiBWWtOrL59ILj4BDCWth7eOHQJFqHTog995XJy0+ij4gOBX
xT86qwToxyletPxsHgf8nFhMs5BNDd/RogLbi2nqdu83k6kMDiDusTYIRFOaaEes2iW/n+pWXQZ3
Bljwu3aD0tdpsbQPcaBU9bvOvtrNs7J/Xnx63YyhBcI70r0Nowl6xMPbTGMDoNBtTO2re42inGpG
NgXoyTXB3qy8bXhnA8DsvJqVA6lPplQIgJarq7qfqgIdMfFjS73XigCvWTGvBPsI9snMxhOSfia3
oAxh1d6ajR2h3v0MLlxvGEY7TszEFx+NHQ4Ltsa0a92GZsYcbNlJZdSrGmWKsDrNnTAq/Cqyk47T
IaR9WIUygOla+JuNqdU1AabqtCo6bhHcoJLPKTson9WIOCwOc01ft2G1hHo2s+7kaYLJ4+HcLuTV
81uVJBzGrF1ryqjd+A0kVZCj3xiFZXOItdLG6Gm5ZV+n3gLonj4yE445ExSIFWYYSxiJk3SHK7ud
C7GWYjf/sV2iofk6ZKJMNysRtGzVXo4FYFVfKACT3avdE5rIIhm1ri2NwafdftHU8BkNGsRTbLuG
ZWI1RxAQYoRkA+nHZ90TyiyeXpZe3FpVxgyeI1wJcHEodbNzFAdLGh40qT2miIqQsafFITDbs556
KMBZhjRNLRL3F7ACb16zLTsXl/S+zdd+oPrqADol5x6bv106TUNwcKrTWfB6r2nyPTnRz85Qrpw1
0m3D9XvxH75ooujLqj7HWeA1ZF0ro2mKADFKd0kZK6h8SOr8xeq882UBGmhSjZ60+7d4UZFKX2nh
BbfG8yvODniD/PGOiVQWxXwpOJxNXqPxVpEuIOx51Awdm/lBux6vh1ilU6f50hrRaQH3LLcN5/yT
v53xFKNSbKsryAhx29aC1pR8WY/2yOYorgOofX9oqppO58f4wTjRS2euwSrVLKWqEf/4eDguxcZR
m145l+goNedwuse211CuTvZlAUkOn4yK4F2GOVqee1P1f4s5Mzf8Re0vTcDoG7/89gw/Qo8nHKzD
hwiyC5MYDZNZbD+qEBfMpEZlqFoLs7aVUC7xQgM2uz+637rHNkJtQPagbP/Ru8LpicxIZbf9tOUg
kvRdiPqsklP7s9kKAtir9YU3Q7Rd6lHto+HuiiwmOF9fjdEBTQk30SRCyroSoU34iEvVAc4Tz5fs
yVGZjBL0IKjsStJll1zodRQwtck4aHnDwnq88k/74rVK33i6sDyi7DMbmzayIyzlZT51BYVhJUAq
bXDhKYFsB8ittp3FWicv06j0WwtLaRYelBlIMhgkMXsoIpFAvof2pxq8Zr0PPYSw3gbjbyuri6bU
OLUlc506Qc3hWH9hj5PKmbt1otZ3go8H//PBuax7Kj4vSnpAdA6YGn3hPvKJgn/BXAgohg8NbWyi
9/SUu0x/mscfyifOsseyegnmfaHOiYKFjR8ACVqZ6riICLJRUVbIkzRxZ41ONIyUwyiG8h+hkqGu
UDNf78nFe/7GhXCG76IIEcur8LieviroVSIe6zhm3nFuQHnwcxqfN3a2qBImh3nl0Kl8Cys3LNH+
kGbI3qfx1JO98aJnRk54uzYCfq70Vs+N9nEjZpbyguoAhKxK5L5BT7Le+btM3nLUEg2KgQobZk/P
Nk8PlxvxR1YIRwB9/GFg2K4n8ugQxm8cuwlB2rFlrQpOlAEuTpgKRbzUkDntjGwx2ef7iKOMppk2
qCIO/jUhJuSVBaBAV3e+SrRXo4ppBnB2Xoys5SMuD0mWTv4eaPKGNh1hZzJsRzNFa6sg9HT9eYVr
vCetCd8HbYeRP8WZdD9f3rp70KX15M9ivJWx4/wqAiiLbNFvhruJ/j3CypsGGb8SM85vzGMXGKcR
7T2bQhdIFIOeXnKgKm9apfDftVAlMMqqk/4aLox4yn0uGbKtCeoZHoKL1kOOo5NALU6M9wHfyd4a
9L5p8Ra62BH99q1VJjSlK5NogouOqhshvQwVRL1n81DFYMv1+/UtJ76ed6eHWCV/MKH5bxDX0PDe
Kk8s9T8eO8MxgZzQUvX610QTySMR45psprsbCIkVv31HlcFsp3UNN02K1HYvvPIAb7XmVF5C4cKw
q5Rky5E+CQk7k4LbjTqgOkinrF+xsVPC1x+HYBSjB97B6blyMQghGZALPoZBHA5TaPx+NM4XR72J
TsQFRH6Q77f5R8UoN+xwqM7YXLETlLYcmnC6KBUHYAye1gWdHN1pL4AvPH1gTr27FWJN0JUb/DlP
ckZHnXulQdSwIVSQfvkmNP4ERcCqfcGK2D2zPqZcW/OtpqGSOApZKBkr4yBUfc9LIOpRr3Soe0Ry
xb5BjL2ysD3BEMg+mM/oZ7lnGD8s1tUYzFV1d+62UJU7wFQB8gcmPzkPgJt0EvVXielTwl5QFA7p
ZTxlGd0PxtutkOvDg3PQiEjFZCRfe6iG3SY5rL2Cr4U6JBmvT2+JAaESNv6zncbosUmkZPqmrGed
5ZUTqlP09EQ9LCcgppdctUybiAktg4P2s8SY8TePk3l7yD+4fdRapUS2oDRz4mfYiEEmUw2IhR7+
gRWa3eEjZtKv68GwnBOmfFlMTcPYBsOd1neHn1+kTLVDqXAovML3ThrV69T0KRW3PqZ7SoWkoMmE
ra0JON5R2uMJVc41vmDoN5jn4/reayL4ubJo9mUz0bf7iHzV0lyhKzAw6E3sSlN1alsfmlev4JKA
pB3RhXlJoO2Dh8jPIv5ybATlcFdD5KSjcQ6p9YDvlZS36g7yV+mdOYp2kg8HzVm9fcO81i9hpkMP
9CpJ3h1n3OrKWValxU3Krousgrah42c6IUnHTwiI+p9Ju6iMHrMpd2ws6jDy4BHaxKE8OwqmP4Kl
6L6fQ7H2KHJ6ZNMSNfdoRY3v76LFs5UN51h0Hr4djOdaWcUFI4ygHxJSuk+MLkfSiz7Gb9SxhX34
L+ifd6CJGv8HU9QE+SE098kRM7kU/c/bpw7Bp9mVHzd6FaHBG4n5FX//x1MBMc8Pc5yV/Y9BldTc
GXCzack3YkezIC/ZNTBhmM6DfBk2szYQUU4y72g3X07Jkom8U+hVKuAWZM+3L8jwy558RTwr2Xun
SSmUE6V0mw0Zmfc81BSUvFpMzplKDQSP95Ix94HUweB6KL8ZZdavaXfDTTJS3aOkcLdHO50NYWhz
jKFwA5ffNX7oqZiOioxRHiU5sN32/SiIl7XuUCGDJfflmJxu/3NYilsgNnVPb8R+NW5FWtJLKcsU
1raRxGfL8cE1oH+WkhicZ9kk8/HyF93kWt6ZkaYcYV4x4+zeisLSBIxTSuTrNhr2axW8edHuyGuc
6yJXv66he+hPVnmHTGBQD/AdwJnremWmhpbS2h1BKku8eUukYXEal8un7i0uihFASMLKf1Fjq7dM
JYj5ews/LXdKy+x8rdGwJ/Kn+mRaT187DR6z5wiMBf/q4b3HLS+jmbefqCt6ZJnByoVoO8hVa/3L
OPoB9oWZn5iP3R58N3ESWcUkVxXUAuGrxKbpeQjFXlDGS7Y2CvlYpx7gZPXqkYpm5QArXrfOM76U
UbT09Isds442+3lO07pIMuLS2ns2BrSQ1tK5BvxFzVAA3SUBLPN+ZWJiVB6N2hmvOng4SJKM5sLH
ht1XZrUUFGs1Yen6HQXkkZg+f4pxmdKdhXFX919B8wcPI/FZaA61br3V/oGsZFJd/05Kj90URRpG
PtsjNo+jbgIfvhx/6GmjmVc4EK0TzkGWNuP83Ig4yujunCh8277JhNdQoeKtRgCAvRHNTQc4m4fD
w5/ChOaicl7tXIltnHO6icaol9wyL+NR/qnaWgsn3HdBuHe3BiUWjY+9ija/e2vRnv6KeBAIL11X
rAJLc2A9HMDAwbIAnHDompPWHSLD7xy47+RW48bIVxSdNyxitRt/8liFV9JzoJriHpq8/z0fzT+C
/o6tZ/F74Cf4vVhwQVHXv/YCar9LJPODi7144gqEi86YScbbkWyavj71kcOAdEoQ3Fc/OAENi7ga
Zxr3jU0w4lWGTgxb5/jq0jEgejZ+lAiVxA5nzcyTISWVh/0luz5AVFMo1+E0aNkj1EdGgUWLFgxc
2IJeo5t06Ic7QB8vdjfLE+8cSug6a5btU6XdCYUTOnR0CN9StbLKInZlsB1tuu620PoTbwh5MIVK
z5n8xSKsL2b9iwcbTo30sRvdOSa3y02bNL5mI5zuiTsmHztwXaoUaTYRtROZa9ttTihMCd74BmLV
ejM1TU8ffb1iGokDxnaNF1n3MLg4nESt4H9ORR2Knah8WVcd9/Ffh1SnLkUgFXV56SzTJ8xHe5ZU
ETpVzSH1EsWPJowzPvngbkWIAYdFfqdgeEuFjys1td+nWGtbbm4Rmh0MEVumADDapFaX5FhVQZmS
jafbbbQr9idiURp8hN5dIzmRY5JqqQd8bH4ZN3o+92ISxlYjOPrj00jBG0zt5bxODfijyv1JpGPh
vu2UnKKFB8eWUHZD9K2okEdXn7DFrQ2lfEEOzNRnCmBAbITNV0YLEprGAyTkrJw7V+MtIpExXL2f
ps8bLCIepRnTzoXZrdHSJ7FOHZIF9tip3Bu0AAq1dW2QqA3zJBrcQpF8JlSYJgGvm9F7krWsjAp4
VlH+C0zrKxMVxZ6u4HZdYIqoxvi5XWDrTSGql05zR0ISPU+V62EXDUa7Ozn0ouU5uZnVbx79gks+
50Yvu+rHWrIIqq7DDY9FjcsNq1A2GiHl5Gu08/1Yenp6w6CssRHLlAg4ZbUN0Tjr4z5KgQFpJGUZ
EPVfcv1I8P/U/vQyOHswuGeKSDOAMWoceENdRtUDHCyAHZEd6ycc5qvTTTOG1vt+B/QJtegIXWYX
R4/N7FbCLCFQOhdKbaX/HJcRaCu9uK0ETx52qsWQOAWuGrM4JupfhfE5fxGN457XpVfnzE1lDZ2P
0YXXBPouQdaMifykimWJ0jzRwC+zuRY7CYn9VDZ6gLPmjG3jdctlP9iyDYNwVfehCaxAVGRzgSrX
0XWzIXH9NHsZuYvuVpbr3kduR9eORNXUHuSJK2elylEccsJBNnB9FE8obMQ/bVKB5q/r5yYyRUAk
p6pus2zbe2B9vXm8t5jlKWjfG2E1F1Sn1q26wGcwf7goqfSGRQCAtm6Ksq0sV3xJyR1JQ5BNSk84
UIyLuFKqFkIgKdxJvYc0rJBtCS5TX4j2AjG4WE9JdE5bT+nNTnNoHUHVivDVeB/VwvWj1B8cnWpU
v+tziC+HaMHDDw7GgdEXdWaw0g53d9kgIUdEkVFkBK6vq4MIv+BGtXylMXxIzZBcj8q9LSDq/lj4
vUt46mpx35EXAuIKUSyHuTAQnD6fsnrJiIVr3yLX1Dzfu6YM4NsngFk0KxndwUyI8hnfLTJaUS3E
QuOMvXXLn1bTvfHCdQouqE0P72zXA1bX4qchRbHnJObyH+6NTw8outn4k5n7toKE7lG+mjGfxphU
LYoiQ4Nv54sDSUYDUXQ92ievTFRPZNO6lmi2mXiAWHwubydXhqERzaqryHAjgVMRBliBfPL3E556
aup0d6tqBtzwKgo2335pjviBscqL/RG32YTXOBBduaWiYf1+kdxnSlZesTKtVF5otYdVOKugbrgz
ZCio9+qqRXN1nwAaDBL+kyAamqDJNb4hGua2JbxD8t5t1dmJQEtiA+WiI+pDwmTW4LAG8+WPcQaZ
N58z5wQalksqoul/G3kNOMWDN6dj9GDR1/k5EApr8+590vYs+p30o++nK9ZbVCKs99ie8ZjyCCmm
MpAd9gZ+Oe2FDXD/E+fQ4rcuTy5O35zZGo+oM34Q8GkziX6tw81cwBuvogX0wH3qUurVhcpEy623
iytkMsuws/AChSnn+GNV+xE0Zvat1JqTk9iGFWJSaU5Eq0uaijMnMoqWgv6fdJuFejfB1Psb0MMq
Y5YvJqahS44EWPP65tBSINMGOjzrudjy/hb3AHKxQGfXI1fZNJ/H4yCxhOte0bs6IJACJqfN+GcS
ukCjXUz5aP6aDxkHLuBx+mSadQPuF8zf4J/+nckR+7lNRXjbGak8ij+0JQZOfyIGh4KoFIraweYL
wJpADEAVMHXATauQ31OGFxYXolSPijgCsv4l9QD9uZP9FfJlbswb7RRNIKNp2jRF2MZ+4mVIEWHe
JyjI37gkNBCBkPJyPDTJSpDyTDxTEpuDy4iGeRddgiHLCFh47TPQ9G/IvkL6sX6pavurHSWyqlaR
KH2t4vCQhH7SFp9gJG69zVyYCHB74+DAWxhCRv6A8CyEX2wUD062ImPt6nwVHH6ega/pgqFUnriV
Ly2LuG0i66eP4kfYMxt0pNm9K6AeSPDf+etNS/nHKO34V0Lsz/q3+kF/fgRPoevoegJQ5MvK4JFi
UDDJTCIry3yG7f2FYBgUtGt26lqZRPUMmBV5YdogIXz1apJgLOZYcIHf3gcpNHRvtOfGV0B0Ntzh
thWnCxX8ldepNG9DJ+603SceOXC5yjjJBCtHHwEHeIe6uTt01962c2HEx3pCVryaiA9ulf+m0TpG
pEgW9MLPaVvQvQYkJC6O55etmp3NTHmozfylZmD/JkacpiMY4OBrd8/gl4RRsmr1y0gcfjeckiiA
sDnIUu6ogO9zW4oKDzI6CoPjty9egaWdlv+j2bRLL59pHdWfSg496goAnxAzeWajEkLRP6BntpIv
hxssGMk2dv/SRbG6p0OcExUNbInGxKzdtS+m56drrANeE61q1/l7IS7/HoFYXotmvgbDgeha4zTV
bWykeEyhqYZna+sE7P44RWQ921tFIsYM5WNjG29sXa7uOf9y6/ENS8Q6+zxSJbrnqrT3FChLZwEP
qRboauVAG2RGxYxGpR+va3jTS7N3geWIEB+kqeOEv1kv8rH25A5JjyrEHykKozPcXpXO28k9ywMN
sOdxg9krk1mGX64ETlP2LNpjupwuPDDFmYdflCPTq++jLET1Gs1R4xNjnhAqRf1OvXst7YJo9Vr3
FOqHXzJ/scsbfEWFhWpUxpPD5pbo9fpeRrAtt4CMRO6ob0tJ2xnizd4TaQUNneH9pzvrqm1EXDtH
MLrTckHONd16o8ZHhxPxtPBYZ81pUskcLYgbA4nhSP4usHb88S2m6z0ViYOTJEM6z4cbehDQe075
A/4l93iVIZW6Hcur8v5teECv0gb5TOkemZPO5WBmHfJFO83WitmkMA4DNb5HoJEM3L7XAJQhQ33S
FJT3/Ia2lnfNZ5HTsVtmxICy9Z8mVEcBr9NcMRNracSjDJt670GPcjiVSkiqmRw4oKFj9kLl5+ps
CzRKU0/UyJ4HBtz1TnAKJuepgs4hwsY7L1As5EDj/5fm6cn9iAfMG3i3XASXWX0gKye6fTbczHns
4bpOMZP0T8YtncEHm95xLDx7lc64pMi29Le5Z3sy5uluz0wMNYi1yM7c1lwQGXRhUJof3iHYTFCy
nhywbAB2Ezi8SXgSJy6pZGw6CyWUOpv5xsPG67K835yvfFL8dpp/BW1Xa7XfTARGhf81tesE+Vq2
g7ZYXE379ijKYCoInQvmWbSsa+xXrXM22OozNnY4r5E3rmMtbq3mo47kd7KnwDhL+BJIaInf2L8R
Y5LVEuH5i4VctrGzRYnY+9jMTJsxfPsIpTp4Vny7J8wSGngFJepKGIeQ199FGp+C1DzYnxRUwhMO
KJko3zl/XCw7UKMNQwus2KcRnIYX68/mOvbzWSpGWqyf2T+EkVJ7q9+NFVvyAfNxANa8uSgh1uLz
2UEfraySKDxq5Vud5hUZ34nO2IBTBkKstYEdVwek+/BcEyK4g68MNk/nx0R6K33oQswhq05Q7O10
EmmDKqSMYruMDZ9Ze/JgRRm7n6Ety3gVHyBl08a8oLrJxvFTszyGe+UEpT9AQMqQF7RSgCWJZl1y
eoskXP9Qv+VOyqN83V4JbqJrOP8+ZpNYfHuLyhtwn9u2+PzF3rv4lWJ45FbJ4qZiaWq/faHS5633
jMCDbz3qMezhE0nNtWOnpvhWJ3Vt3O1wMsS6jJ0LRUQh37AyZYk/UFmJ7/atpZ7ZVHVowDDM2o2D
ZGUTFW7UPBp1pv/CS/jav++mFAZJGDOYoBB5D3NTECmTUXvIT+1mRCsRN7KPfhVDaoGF6u23DN47
f8FshuRch2Jx3DAVCW8YII6sunFImFNTo4QhSGO0aBkWjgaiNyBOmQ4RryVRWqCkpbBvYJX660NU
lnFTjb6d7OeQqVwObvXNkbCZF87BPASB+zDVDKqFG8+ijRkEcwUD0U5il96zcIcuY7KX918cx6eE
ZuJASr1x0AkgTLDVstEgdb1BxjseId3u9hN03ubqwiZ0QVR4eiU0kbAp7S12Uy8hA+BxfGVrBNm7
nBIWafzmSM+uszcluoFi++eCi4BeJTrHXCNP7f9ctQqh6muUPGLN3NHCD5M3DMlODgTZkEsSKUOJ
SH+85956U79NJSMWpFdW6fzWWMQ7W1j8jV4fayOKcX6s3/M8BZhLH+oG9nKJbpL++8ktQbR+clEC
317ACM6dQkokF87hRvuvX2RywzLSiDHPpXfIIlVF8WBZFzNNX3IYbVOiKz6PMwytizvf/qh3axD+
6xrHxI0zG6M435lHI5j2M+S2RN0APesIVDQm2C0dWtw8JQcKpcOaB6EWuNAUMJFB1Kegord4kRMH
qXY8FI6w04nAQGLoqIoiFSQa2V1mnluyreRUtjB716BXn1wZkS3HCm99V6lnqxShlqFV1m82Ik4x
kVBfrsXfEFlStVCEJHoHugJ1xQjmei0pkjzKzdhTpX4vaN3cUm3PW3QbXbG4U2Ok1GDVKKUn8UZo
6MyfjUCcC/Ar5q9OjI1mgcfyPQmMa/SF7WnY8FRK/LS0tVyX8v5HOWuyNFM5Lqr6kxqqrJ1sgEh1
knXGDGfSwFgomqEw5Iy+9YTva1Ly8mCJZFPEYr+q91gcW/SgBBvk7U3DvoWjMmy30kM2GQhz+4jI
oX2WVQcZVpIxLmUbnV08tBZDtXb9q16bJorMJA6tTWFhYBT5Tye5kaX1umCNFk5YUKNQdnVrzlE5
cLWq8sPmpnIRjl3wCxPT8rYfBbHUOv51MxcGk2YqLITwvNixgE3rHjGcOuHOpSVqkizNmpDetWrV
P4Ca2dU4DOVQ3+2DWtBok/nekqEWeftIQYS8BisjuOur91Yz2T8mNIQRVn6euz87H7gBrDd534f9
eOJp+wqGcV7AJKOEecqE3t9gQmLhQ1Jf/eIeMt/lCiw3dQkR/niaYL75Lzb+I0ZL3pb7oHuqMul5
AteG2yTvnoClogAwD6fKh3Vxvfv/kxKO7kO+3xJvtw/LsRaKMsLknZk3gzl4V+fSVbhdJ5ZxLfuj
dRrq32UEohBHMxe2vy6fbJcJr5AFblJZe43XfolpNjaxGxPtnIbqB/HiQiX0dOlrdBGpFy1Lc4qu
W1AIDZBOYsqQ5gV5N6kCr6qx42ln+r1Q2R0BkwMpH7vxnMQS0mCh2ihqDO9exfDGuSneFWrs5wlV
FE+NEp1QWC4C2cvZ+bfK3WuC7iejuWbrgtZQzxnZtCeoArD2jGfbQPJxAz+5AdA5wVC34NkpRuSy
rEG0Wavwpme/jzTf1Nic4UR8wZgvPD+B5fJXNMD9ghsV9VeuElKkHr5a/Fh0QGYNnIgw/xYAW078
4HAifqTi3GFmokB0C4wUZvURwdYa3RGNA+I51E8NtekXG7oAfacsvh5rwYu7Jxr7ev80QGsLdT/E
QA22ZoBNvGBxeS6diF09mrJqTk2gsG5+b5DFhrf6p9EvS1/VPTVoOA/UUQoFKD0gdAsriXXhLxQO
/zjet7AHzrFEOGiGPPJIJ0tJ1Z8WK+uT7SyT+oVCgb4ASTj/ns6SwEMGI1A04igDooXdoV9A40MZ
mgqv/le8d5utg9/tGbcM0H0cjs/T2sQB9nYQ6v8THXvmxDbpGnuYd190NOLeGfit/6HR5DNek761
KwQj+pfg9+UYGVOC0WFEgTkrWCERtEuWLHOuQz5XAgb33Ks7PZfidXA3dJtju/2NNDNp/IJv0w/M
obrC62y+ZQWTwIL2wzkW1ISbhj7unAZYE6+P8h4z3xQZveb9U7rqvoEVV8Xmu7tUo154li27ddKi
ZPWPSCeWi/nsYz7x/8k0o8atlbwZxpKDSWlVTrZi86okwVBMmevrxKqsno72DF6ZrlbB71/CtwTA
aNZshK35KD12PAj8L+pyKeQrAoEIlxcLSuOpzvWceOQ3LAQiy2t1F9wFzy2oXUjQRXCaJ9+iXosJ
smwUy8bDEFs4f5+GahOq2qsohjxQMh5P/f8KjnTRxKJUe8RRpPO3Mh1Qe/yK6BpL4RRciDNDOSzk
rIkR5tuDXCaT7Qd58RuIk7NbEOCFMtsw3ELBoZwUBLfcOx9mVp3irhxlpap8STkV3SLTVJXivYTY
SDXC+BypYDEzB42KChJ+3hPcnP7LI9bPeD3UKd8EE3AwOvJx/PacNnRF5JHNOrGvPr9qByYH/iwc
21vKGcqPPSAhRr1RAXMwBZjOiV1oPKgwr6ybP1K4+mVJiZhiKX1PsVf1zS62qTYJS6h264UQX7Uc
9S9+fQkiTrE/ndfQV4bMONhyr0iW89ioMhgQE9vJFWABtsnQofiuuG1De0hBFUGjHi1nHDXLnKmw
KDfZAPrFHNnZy5hBWGkWAl3OCKgdeNSMQR0hzroXse263Cd2feSmbdMqEH6bShwYS18WS/LPpNHv
k1iF49WXMLE2TxDaidaEDYn+j91pjFtKza9698Qyi009XRm9ucKVjS0vFNTB59pYoNuJgez6ZiUZ
2CXcJ7r1ttd2JiQkay3lr0OghQrQ89WdPIqY3DohOARJwZTgxqQfyj6CZYUO3l7lq097oMbw9mNp
/ihj4+tEBcA70izmvPov5zGR/FA/N4N0HC+hmTrTw7hN5Ibsb646JJLrPFGjzAL2ueTun33cPD8O
T3L9rEpypx3dVnBbeGL/9EwpzMhAx49ZV7suO3utR0z5eIfiMBbYFk09rGCpsmB1MKBqAc3cXsPY
fb+85mAgbLLY0VqXAnoGsmdXAnZ+mYv2KGYL2vldWrCzKowuHflqfSusNZfHbs1F5Vm0e59qhhFq
Yw2+joWyw4dmVPhSnTFPRQBnSaTZiY2jLbeGw7DthVTDHKcT/YWr3ZqHcQTf/33jDb1sSI+VxMKX
PK906aBQiijtoLTJ28afHSQDz0TAJ2kUIw/87MGsx/ngTVJ7lyLn24tc7aiRr5sK3gcEfvmnSMm/
Y+n26Paqt24ALSd/DzEuriwqAlxV+h/f6n2Wq4qBoIZYc7bfoX8XnFApKg5dDH43e0DfToR4ako2
lWvE1HsVtZk/sXG3r3lWyfv/KtkVL2+b6w1wyew0sdeOlTpaiv//TrOuA4F4EDrPpBi7z+U2pJ5X
U/CW2VL63xD2omPs9hTlDyx7DPU8AdtLRxC3QgA2KNpUjnYPLf8kjOEAs662rWscje0u5t14j6zW
a1lD/zP+L5MMAC+P+AsHVdpgWaqgG5KYVGngI7EsmDUP254IUpi7lTRV42r8XhdC7pMDBQ0HrwbJ
Bt0ZYJTg84sDhYLMwcH9H7RbhGaz2/ni4HhL1+9Z6QNGSTwvgQdYiUz64kG2HJlB7cMvsuLcZUex
wc1S/VAta490gbF7ulsnz/XVjcfT6F4TZiG6uGqX4f00xsxyEtCXuUV+cyOQMKJ5WC1VTCHd30Kw
uycUpzA9yK10+zRriXPzRLVWo3QIfOof2NUyRDTtj1A9zX/gFfs08cQH0J3n7uBIrvKT3KpH1ptV
acWVoGh8C/72T9etbU7/esKtrnMnNdSkGvsbRtrb+Jjk/oEsHXwuYWCN+xfySaKPShXhzdM/uvIb
EgtDaycVtcBnjSgo/1qciB0FgA2kU3Yyp9rrDGIYV8HduH2Ni4MFhRaEYrjrTmPXoXAn9mGZe6fw
RsV3J5Dvrw4y4JUL5V6AriHxK9JLZ60a1upzNqYCJbnNmXi2WmZbTzZdnltvbnht9cwjHmwFcYCR
iBHsMS6v6kC3F028F/x24I99tj9CAhlcHekIZ6K9E1pOhCGt+tjnpjz8ofKo5dirOAEN9m2pImso
uqmaAuquGGB0a8Z9HIAcOz4zqRY5VbAtFCpIVZg6kByBLVYPDwusDpzp2o8C2QaebWgaNhuFPxKk
+kLMw3UqekC7aO3wBK2ODeDRgqC++85pq1SdgETw8hB+JqYW0GQAi4nfx/gxShuETjy2He1CoeGl
8kmKvnAJy6pkO/h6d8GBFqY66WWMNvdOwKJtSy1bs2TJs+e3j2+RwmCDPmlRDQeDh5g4gFq/vJfu
8OBNKImD92xq2L29w8e4WNHA3zH/Flo1BviKroEzO0/gab7tOYziSOpzj8pn1P5DlO2zWfFcjuzA
otEOU3uhwsovpJkACtSBKzD6OyLNUfyNr2+c5801lqPO6oKq1HD8Bs6vyAbnGaB2+5BziIfXvHM8
/VtBWLGowncy/5tHR1G2MncCLt9UCVv070O0H4aHcfO2kAlwPOlxn53LMF/C0QL3DYLkGrIyVZJi
u9D7Zh4lBqE1Jn5dffq3hJtTBY84nMczsf/DJARVfUTaa+/8IAQSVU2vtbLzAW0syvuuiPiBgrgq
k3BdKRAv3NZ26Db0k3fRPMD6rXtJ5sWwVW1O7+D5v301cNaDQN6Im5HrgbPfR++IEgp33uSED5H2
g+1fM03uGKHw+VXKCXimvfbUORFzw2W93J+La9yVJBPB2l4Qc7cSNSwJMHDW0UqXJLKAf1hwu4nX
lBpCrUTIM0Xd4/XHQWHXArhP5kMMIBIJhQdS9O2MBp2iEcrir6lAQJ1JSxppfv+Q8J+MSaCFPaQN
VfQSWlff2xMUv/5sV9tZMOM4HhBI1hHnnC3WvnLExCCjRxyYmvqDTGs7JlNR5Fr7nWH6CtkkKR0+
N1ejuQbd/kRnNMxWJauTmvNquLxmGJsPsUhV+BUSWrSEnJFc0tDp1D09zaj34XgoLYVbSCn7GfY/
hZ/uYPfN1H/4klFIvpT1L+/YZ5DXglC1wPRkAqlsQ13rGxtMjwlo0T8JoODlCAGxT9JHiTMuoQaE
XIno3UjxJF3LOG+ovMv18NFynd599028Xi+NNpVSj33dQfk+JDdykel3HsDT683uSUebCyfEKyxs
+Z3s/06VsEvsZQTLSSy6bpKpVQDdy8cM0lY6jJROsrgjKybGSFwSMqqFDLYXaZxAVBifKXDsJbNw
zdR5SbA+Gj+XNmU0N6bP1E4uBN/hjAIrwz6HSUOLlo3CDhMPUbl6D8xL0GSfIx1CjuvqUkvraQBG
Qvg8Gd/u1qopbHPS8st5f9gp3ADk4lFXo69VF/vG2A6+swJznlz5x+3OaYTlqgQP0067DD6VnQA7
dXcWBjcbUmXQMz9E1nNQ9lgXDrJdhXNYRH07gWJ1ko0FtTNW2Xd4bPoKLa+o4XK3xLbaXOliiOx9
NP0N4t8sG63V+bTwyytZf157+gx8v8fr+Jjl6l1zA7Ex+lZWP/d2n+MtW3LJdEX4NIndd4yMsy3L
F4kZH8wGhVp7eqgWVFOlGfDaHUU4DottZ3W3Ojfl2io1KYpYFh/aQc/CVu/cD0dMqWC/w5m+GObf
tt4Ozrfxby++SDmhRoY2iqyq8pKP8U0RR1DuTQUjQ2dsvmIcW/hS1iK0LTa567bbFIumn14ZP37w
ngkCoylavJm/vNataQpz/zUvTvCpbFdVudSZUfZuMvhJiMmGgmpi1w+Vi+AZ4rcwBN5sBrM/ha7U
OP7zBbrMR9PZP511iFtHw+E+ToTJbzWNVC+o4e1NzXiqFZC7pEe/vvKcGFN5VUxPR+fv5aOTgNpm
qL/UBARIyiSjzctld3Jhhh+pXnQ910uadP30FPj+AWs2DAbPoGy4Th0OFcmyIp0UrukxlGGIhJBe
fvit8n0Vw+IEQ9mr6EIYvs8MEp+BHNqWUD0q4MsGTirs3cMcyG0vY7T12P1guzuC6nByQBgV/cq8
BEzFJHbHbq3ywa+4dvamlPoCbo7LbNsF4Gp1CZiALL7AAFBrqwXBgDKO8yUeXa+VXkk83NcG4wBi
r9fG/7x/v/rPzgDRXorYEquVGmvG/9xs3UFU+4qqzD/4f7Vxp4DE9fWH7BqrixWezfgj2SzUwVw0
dq9Wm9pDSfwAH6biNU7zUADAZ7AmQTrQkUzT5F/Y7rKWMOLRx4WzJfeV41wcDnJyTjGIUlOV5X7B
VHmx11FVpFj1ZVdL75d6v4uCvKtwm35+P1a5ofXmoGlryE8PEIxYW6clZOG2P7e1/2ySpLegACq3
EgzQlXZ0wxz5cu2/oKZ7PAb4uPKpRRTGJbZbh+yILmCWS1wAN/4RX81M3VY3YQubfpezarMXWPSS
YncZ7yRfg3zG6cOiVzt3LloX8hWLcWB3hdsQTKXjd4DarjzYnf8EUmLYZ8UaX2TZHH/NKEy9nBJr
xsPnm6sOVz8nK4fNyyd3BNvjRchlM8w9ty0AWflCU8Og1Zw072k8qOF28UMtfdjssGHj+aqHi+Gp
89EqU9rOZUFwJGnVfa98HnvaydHQMpuNE1mY64d9VYLiwxxSNR7kMsiOYr8g/7x4Xj8xUmSmoo7B
0kghZWnPABag22xRn0H5RYG5CdjcRYVkmhwd4VXYyLcMeCo6av22VSu4OvKFLFuviH8PdHJjz4Qm
00Dcyg+foVzNRTMzcsRXW3RRSTJ5V91RHXUeDtkbxIqQexIFsXdNBjyqMLZKq3opbxfgVwb3f6tI
C9PKeQvZ819Dp3Whte+zuVR8X8DzP4DgnC4YRwgInb6n5+L7BQb9XG6I0sbH6jEzGuDwsT7Nqbnc
pBoJfevxk+XCcmfzcVVUlWK2GIaZ2JGkPsszkXgxn0ahOuCpjyG2kt9XSErNwvZSP0XIgM1mkszO
k8fkXEGWAd/Yqcjh8xJUwJ3RKl66wttDc1enbEiv31eRhzx/reZyaUBAogDBDbKhALFHWyciVi3f
ntd+k4f+6IuMXjSGc890xWHCFlla59E/tYXHo1VZIOE6RdH8p6Fr/nCoMI0RteoJ/IjDFzpQ80xg
McV04ZFfnRwKUgI79aOoGd9MB6dgy3vBCFH+7GYe/XoiBauE86OZaKulMAiGQxlnKzgqqlHZfIBd
MF/jUT+FrEi6u1N57H3ifzfWD/maw6nL22L/aJ/qZkfz936l0waz1UhOvYbap4Ikc9k0aql7J+/V
WOxBdbEkkKW+jrngCESFBbcsweS4hOKrHJS1ze3zeMqHYnweTT2oin9TxYgiJnZXcZRCC/9xLfuO
3M4eDgydYMHcSfAPorhbyyQapyiDtzI5vpbJuvqybCBhhIiF25QH59lPlrue/5BUn6OfUgl7NwhW
PDPazaU55/4LMneGm/T0E6V/atRANy5/mBrGHthg3z7SjtFCLxmAq11cbe9DL5sDiMk2CcL2wc7W
0Ekvz5SvS0YHlVgSHn2AXnloO5/KkrZmDXcUTISrHcuq9mQ2dXo++i5f/YWq6nI8HilQvdVCUdfl
7IjG3klWbUepB+tXr8QSh0rR/cIc6QNOEme5FmFlt9o1SYARVO/FIlnw+X+fFkf4nMNu9AYlzNVC
grAQp7ypLTtTm+KJGZg5V1zlAI+nLQ5+SlSEH9/XlH7terxLSv/cJC5qd6iv4CW+SvoHdgliD/gN
A2nP7AkFnA7EHjxDoMNtXr330vvSZ/HqqNpjB+nH7a+5wfY5gy6YJED4OHxgv5JI35HKs2ex19K7
ZWkorllFOQ3rAatrAPBzo3ehrU35Yg9HHFiPrQd6h0Dqcimxtl/bqm3PSligPhaqINHMuWbA1NIL
nho/40yS3764IW+EytdRfJDw/Y66RGCayxu6bF5s4WrnkP45eFLxk05hSegZHTYT/nNm3p/FrDgr
i+gcnTo+rQRcnTa6FNFmCwce6HJ6fXoJuaQJuBCpuNU4YRwiGUTkzqQyLD0yJproMTgo+ilbCAXm
VXsZifTTg7tSYH6PNCdmI1s61QIkymJgAiFtri1q/DbLB/Js1bT1UEr5UGxWGci8QABZJ7nAMQc7
Ob1R6XvRM0vfOYrqpP8EUFJvLd17XebQTe1YLQJQizy7n81u4z0wF7TQ2HcgloYp9XXkffVcQ6fM
x7i/yQynmQ7BICorCHMkkqakg1TlMkLVDSF06Y5ijCd18HY2XhDlCJqLmW1GNl2p/HN+38LyLeYa
Bkhf9wcO2Q9VCV19bdKwg4+7RIiwKyzA2Cf8FvOrlmXwOWH3ZOR6qD7SKutE5pufyBlS+Jh4SMN7
KEfJxCZuqdzI9q3dcA+xuSnfMDu1CzB0wPjSXYXsyqym6kryQwfxJ1mfjYTgcnHtdczrM0FIQTaI
DZXQAXnptmlbgK63sFJDoLQ4L1rH4XpV7VE7mrFO4WdVFjKnCUamFKiAush0+pH4XKGicxte0Amo
CZpfSM+11uh62NX6da+r+IPEbGG4HX2pcMt2W/SmqZaKDC9PsXLb3Z8VLzPs3LqeEuLIx/BlHaYM
9mLJUoci8vd3+7SWmWKKUR57iPOPXI+nGCf0eiLi1kKQhlWinrBE0UmRDzZaFdHVDWtS8fLzMDM2
VZlOePLRQxFRd8PHqs/h6o+Nsor8R75Hpc1B82Rj2dhZnPfo19UzgUis19Its797Z6cPhOfgdf1/
0oM+GdqE+Iw7wJ/OkTghDYzOG8wYx2N7GK0Fi/mwTvTnYUUW3lVgO9Mtikm5ROAcXsrjEJBkbY8l
tC+TBcNNwDiy8vkek49yeLhRlBHztZU2p9zTT0Ceo8AqxXuJTct3iy85MASbFwgJZK8uD8sx4pUV
2kVufsAVmHhqfktOK+yoZp9T1npsT5pdIsBznxDLpAqzytSXD14mnnhh7aO8bZxcgvjqMaymOLjG
OyZY4Vi7JEH3okdqxOXvAum9b8xfp5o5Xi/3CEgcWri+DbOvxLAx/OrMnD1gqm1ahFk8SrXA+EyG
FhF1yx5udrn1eyen4m1JhTGr8o3vMBBhPhJmx20ihENDOUeYFbUunLH1pg8b6dm2QS1z8vWrQdbZ
rLOG3bkj2h0eePb0aytbNSi4EI6b2VseXOTkyfOhFnpkrzg6ZZUTPzWNDKD8HqrJxqFCSDZZCPlp
VWX9A3Elf0x00tG/0fTZjLAUKq/VdqJAINFwruMBUvqULfnpES0f1MPt0ebipDt7Xsi1yUSxdw7l
wK6r0FXmXAPlkZfoESrJyKrIevHAHzv5Gqd+MT0/838VjbeMoiHyY2M56b4jjcSwx7StT1khWK9k
qqplo8811FJXuaIGoo3sR5p7t4n1cKwJ0Obmh3NHasl0GRMnvqjIUu7y3ORWBSqynCosrUzDCJKB
7U8dVzLcPcQ03n3HIhWXAYhfBLpB1O1fC+02oT6KPTiMYo9DmJWoXvBiiESxBtbGLun5j0CAkR5j
mVKG0/2Eqb2UD90Cwf/vkEij4R036u/9V5BoMowfFFSItgcKlQZJGomQZ0xmRkPe6o1bT8ioIbk4
YunP63W7XdPltgmpUaWs5W+sKS/LUjcjOnG8nNEQcLJHJH0CT1I4asPDcWP2a3MxDDV/ShHNaHCs
EbqZTspoNDx2OP57i/OoqK6FF2lYVvm8fCbAtacolo7FUtwYpXcDQ7Zk5XJDckaMjsZvOBGTOTMa
u5LiedFdb9pwF/sFnpRq6E9vI49X1mrNLS1KlBaqMM7fUDsKaZSPZLjdVpe/KVA+UO50RRLxfXIT
qiDIEM22Kj5yEfeDEm/RgNjYcWniiOZok+VOTl7WZf0pTnyywawz6vGA0FaWjdmBjRU2zDGpzgbi
/QsRdT2s8LJMC0vDu4SLgdqswdeqmS5mw1io2L/8GZ98MlrloZM1Gh9yId46UJue9Jipf+nERlmj
6jBqwKS49absl6t59U9M0EAVxk8Swq0Pne/qWMkvODvLJsZSeeYQwXzwgy4CIF4L43ZcolM2ud2K
kKV4SbFQ4EHpRqGxh1UPuK+gJgA7xM5QNESZN2aTK9WSqTrDS3gi3pA3Z1AXHs/p+e4XJx0uS7XW
jnf29pek63LWX0m9ihtG8Tm03xVJK737MyamIBrjn2I7lrAJ86GYbQkHj7PAmnK1veQbPustpwc0
yq9icCkOU6pj43De/GV8udm78KDmgpCJOveSpYp8Jn1ToLc0RGQdTGnL/X07r4EciMFptm7XJzhU
HKG9cPsDGQ4+2dCaeA4vG4pcfw9+I7XJNvTe68MV+XTHQqbqCTIVOSYS6ZUMpmeO1PngW49omJnw
YMkk0VyhQKgP3fgSYAHP2aHD4yd9hZp1FQ1LcDXdRmdCrd4w9Xjok5YJQMM3HcNASH46mFYxYrGC
hBQTzqz/DsiRkbOpe3adJ2S8zVcQCpkboE9tS+A11FduBXDN/8YDdDHIYWsP3MH7exeTfxfqNs33
ys5lR9WjZYMn23Y0Zs+Cfu/CpyopLMGK9EqBMuX4L7X67xxym5GNYgcJRDgUMR3lf7NoWCA7Y1hw
uQ5KaztYuYxDA4jElVb4mjCwQJbIVGfBQ1/uWtBzyn5KVPlkoR+bYHfiD7EFtmmIGiwS+ywJuSOY
9Mbp6nhwC5QbF0ttAEQOjcHCV60tiZdcnZyDI5dH5mP5yX9AueLaCG12H0u8XqTaTSzAJuN7XSTi
4fmD3RRYgbJPuxq+BmkgxlNmF5808ss4meuS1tP5J/idUBQTmPexyt60NpcMktDvGUq4R+OV7eTc
v152FcpWvUpJwv+NWQ5szyi779YEzMJ7ndORVH4vTOLPR0R9q1jrzBBf5Ed6xgbeMmCoNqPSIXe7
kRmSKtSnE1RAw1x6SCawBpHFtRaF2l4iuxHQL+sgIGhGOofD4Ufo3v9OHXluBLBs1+L6Zo6F839c
kKCOAwI9ys5QNzUlVPpWBGsm8llnC5iWEbu8pJDwXct4mlfKyY7ghDWp2bUBtQm0Qg4V559TArrc
6gm/1jEl5/SukF2SE50BLOA4bGX2UwMEHpUb/w8Br0OEvg7b6IRfRPROwOrqzYsYAuAqMxcvyLTS
eTAz/1BBAPMJ2GjYzSUAdIe3H8tdODz7cuS1k4fhOlYEt0FnxSY72EBmuZltzYpHo00psUKXvqRL
4cUDfMZD5WkznCPB5YoBdX04ajgeO4aoubTcBie+1R7TkZ3ZMlM2RZvVApHs4sQMri0QEW6Hps4Z
B4Xl1DnGHGDc78HjemKi20hKSp5ULQhnRRfKIdUoOYyyjYyCgyis7tAZJCEcAw+c6zXxtRqSiAbK
LmRuxg+bGowzgImdkuQHUnAxymZ/VYXNM25YgGcZpx9j7UFHpZK+cKSOQGZB2XOuUVD3Oc7geCRJ
o/NGCC+TbW+BQ+dY0RqQRY4ysnCdmWScGf9cl1Sv1Xe0Uq8E887ly+Y+4TMu/EHC02H1jnt1IcML
T3YSXaSJgQ3Sk0rFW8goFmWUMcPpZePiBVGcODI/Y1+mRpM4nOEVseySMSMuS24/aLrUAaxSO0DY
jqWQk9z48Go+E1Imy5ZBeOyPX6e6WhrDL+6kWiAocI887KsNe4F5Kb07nPz5tYhsdagmDZbLTaqv
hV4dpV8wqCLredZPeuAHSvMYWzQO6I1vCLd2YwH/lpGyXjJAnmMM8+ELEFIs8oOOHUvh0TzC0Hdd
gCyCiWhoqzS/2zOzDanB0zOHlcJi/C7g4L0NCixFSNY8E84kTLy5b+yNnMceQi4+Dt239n108NzQ
lgaqI8rt4I2HJYc3iTEsWW14ITZjx4liigvgIMCgXQqllBCTSmBX/4WOjiQKmvYN4eLxDwjcdkFC
aWvNte8tt+xR3PkzKJhYxW7kHdV7ivoBtOhrH6KZ3u8Yv3e3G6lGcF0HK8/4UAY4LiPYGSCMSmGh
GUw1DPd0FZ0C+bqLwEWTF7zuBroVSPGITLdNByLbVT+xWxoY0jWOteg0sEkeHqgUhPRH7qi0mmRU
JPGISvH7d6v2ccHpzWHprxpJla3yi0fZbeteXo1ECEzAYBiNI9uTnGy3F96aOD1/l94SUYLScksp
1xj6DfEaWA7LO8kfNVOfBO/pToXrGbgKD9Vs30cMPkwIbhLZuxWv+QDOp2FhxjoHwN7w9hmZ9mxa
beiYubBCyIE+9gCb2bc3FJ3BV9r6N9+K/g4nUBaun/0X3g5qw8I5zu4+TsegMogf0xi6WG18aYgn
XCIfzBfZP1loF6TUwR0zv1aL5p5NnkATU3u6G3PekiDMtWsL7KxDmTblJEdK53+8v15peSm4AOOm
//adQOSvWtCGMsbZZi1Q8Ouf0WqFEP7nuD+ujhkBi9uMpZUiXdCSowkghgF0UJtlN7ztL9oLceDU
qiXQS5nl9RZggDqhJe82codRIjNlahiWncEWKvZ620Mx05PkxUAMW70wHSZm4OAT9r2lhbj5ewyf
ZXg4mxb59gtmoxtdUMyMvNosFHPnT3+w0g1NOdeObPySQcZPuDbI0vPi4h0WHpZL4vFrz/WfEJBn
dUIYjdOYi75y/XjrOzsNK1F2eTlItxT+i47CaD4VVPo9TFfHm4yKqOKfh0eSDQNgnAkuw+mrH4N2
cciUs+yy/KN5S6LZgqZlTXk76UX+btum2QVvjgcljuyu4pOXkR7NZyXDr1QtjbmdRUAob7KPlDlQ
1bDKemuVsf6spgPbPdjoZ0JXbfgM8QqKmsBpZic5snKhAEogkkDCiEBvRc0CP5gjkaVoDeN3MONX
UcMFglls4fjFua8xiDXw0Nvsmz6N+PLmnBottOwTgXxkOw7AAzrHgRSSJj39BpWT97Q5YFFBLWQU
MALwbnAf3OlenR6lHOjKplXUnZp+2bYMt1W2NtcNJHTt/oTbqS1QVKaqLl9LVjRSQ9gXt9GG7m1V
SHE+badDXuYx8wbHUQCNvOsTTIyzfbMzfBWHiyi8Wz5/IVCM3FvfVtM9UyMFPx+Df0lawLgq9l8n
UVbUgZS2f2UqZujgZy+KiZhyR5Tdx3IrbmLIvANHVMVrYp0xRcz8uPY7YtFh02fvp1ImyEyseEhZ
ed39nHty7UYUU2uqmWAmXS9Ba3e+TJq+30HRq68PR4mEbdtoCx6XvyTk1R15zS8GDLt9AZIVKDiv
z7VpeeMJd1h5zYqzQBzyJS/pHFXLD3kBQvx4JpRWt0s1R/UPM5cyYhkr0uHHQKxh75zSuG2kx2y9
nyc1/ldtNOwhR63StQH+9Q0AMy1ZJTkafyTAoxHI7Ps5tZm7/diYRTvE1+vv9zi6b1EODOI81nT8
KDVgPa0JmQyN/XBiD3aSI9ubsFw8tyBZD6ApQ/aqjY5toDVmoR9QMFCZJ5BKRoMNX0EDUTplCVLB
CuB7F9VUJrYuuTgJPHpvb1j8ZLURG1iRlR5owhEJ7ix+yvqXCpsujxnkInDwcDaZ2yBiIUzdAybZ
kJ8TXuNE4ps7dUT7GM/NMs3Oos4cn6YVgE39A3wCVPfoPzGaM68yOYOoH43nRA1TBaDjFlj5hlIX
3lKwkkZcv+qo38/U7pBJmQNYgxWeM+rorictubNaZHo7zEJmU3YPmdV5v/Pt9+KCF8T3Q8URYKC0
n/ZZoHAX3rUfMFNiEJPMzAiVN600XMBH+LlVRlvRm37ck32q7IWGUANccJRnEHNkgTB8BsvTz1gv
ygxk6M/ctMsmnYVd1stufyRmLEunKeE4FSmXEDs5epwldRpRh4IM8SDGdvg73KofcpGh4nlS3fKS
Z9c5HeATGwMzEmtRS+yICdjHZemGutSk89wfMhvkjLt0mLFwwQ8ESAoxhw/c9+oGK7s1r/pDDfH6
BZKVq4/H2H3AeBH9F65BobALqxF56ZRgNl/pdZFk/ULStM34ALgh8C0nSRGqUnX3000Qkq75LiP5
GQB/rYr8M7GC0FjBbk5IihYdnzMwWrYcCYIsJkPydzsNWIhF99ErgmJrup4bXYqUHl+UxzsEno8M
zwF2qnvI9SOyowzz2dljMU+lXq6867PkkRWGKjsRI0WTyS2GlA0igk/3hJNDmjszMqMRdP6ZwxZW
xCUqEeX+MvEZfNR0N3P4sSbm6qYRKjdp/XBkUrhLGM/iCyak1VQS7kZtCb6N6VlQ3ub8muR5aBEq
IQ4xAXzxaUaQn3UbnLoz7tHQp8jySlK7059XwhGM91AtgF+rDRLYwW0byIw53FHoi32jox0Qwsnt
NmnMv9cpLg4oW2C/X20mEn2PG1iZpE9Je3WxLR2fueHuhLudjOl2DcmPtY8EKzNQZncMoZ/OuQEt
J3tsbVL5z0Cut1duVod2hU6yF3KkY1mtM6RNq9y7NY9+7O3wzT417TUjAq/Wy+JMmWgiiCu18Rgj
LYN+xtxaN4x8GUTAeFUULbhMdUFe/85IPhkTIQ6fTIsd+WFAvZbHJKn59zhrtS9Q2zKXUgEyCb16
/rEGtNEqagLsMLr2a7J+tEriWD0Zc/nu31+FOpYhPPWh94ZLgEs8OO85os35tcRAGRkBakulcJQn
0mQXF0R4yhO6OpvA+0ZqLCMzfcoQYBNm7sYsgHUqT7RuAkMnY0hpOSB28CUl1IQuv51ROEBul4ts
dMORd60eqChwU5RUeq5HwmyGkBdD1ha5ExhB0BD9N6zMA1FvlLnuUMpgei+emFfeQILiKJU1/zHm
Wbj9ZgdWeOtgUMFiqbe7DwTTw8rKQE3o4Ztyck8QhRhpPsUSN+B3K30cWSInX5KleYMrUF2jbCTw
la3c6SxkQAHBzSpIrOabUff6/QYgLDIf/auHJUnee5zEzMv7pxdipE/rq6Xgz+KbpxUpazMUdVuk
noT6xxy2CriklOSUDY4hLYnyQgcOCSEFNEGGcgHAglKGoHnCK3SPHPWl4cxogOotbAtuNvOvCSuR
11iUCBn7fL89dQsylKYxHtIxRraHWirVd95h7cC9qhBuSCqLOZibQDr6n5zyf1Rp083g4+vGpzUk
ux597g8S6N57SxtWZje7T2qyblwNPEYpUxZEkTvAIrpzhA7QyFcGkFAX8vN05AWzllef2uVnPj7t
BGLCYsqlQwOZ1L2f4U6yglXv7p1om1b9jBetolygLxk3rkZQZ0ddHV6NjYn8ljgahXH0ogPESfjg
u140/hDV3dZ7tBVPkvuJPC9/feRJl6KCXfaUgW2Gyr3VAh/kefLIBeQ5LLrGHSCDu3oTL4rwYQLL
RwMcEZHS2tflB3rqESOo5LDdO7qr3nkn02Fhl0MiJYKBnZym4q9mZo8OG+ieR/S/URko6OnWRXDr
WA7ZmRp2rv7unHpfXMDZRtHGdCw+hO7+LUzyZXA+TQu/JhFugvvMbhS79ZjjIsiCPBL576dfOgUQ
ibMGZhwgNk8B2gQqte0sPZsRXnM3UcK87eo2M7dzj3bjJGnnnOhtieoQ1y6/SEEIEhN1S4XSVkkF
vHkDEl3rvFuX0nl0l5bPI0VN8zTxZ1s2PD4q9uUYiwM11RF25sW/Cwlb24MVkbGqup9sUM7PB2VU
TQCA9rG/ZhJ6EjHBEl8sqRx8Bk27rYJLH+yZueMMD8Z/0yap12bpGvY8mIZb5EdSQriAGuqv89AY
dfKxOgvbdP5Wh5uspUZUBkbeKkFvAt1Krh3X2B0jmgx84eQUDwbhQyQxyvq8+urud1pujS/vKX3i
AqI2+/hzv1WnBM4fwF12jO1n1gVUecvMNTPfUYOVOgApJGUTJG7pPyRPrvRLl824zjMHCcVQsVlw
0am6VjGKgrLQVdDSlWeQKh9VnauPig3qpqL89imzGUctLiy923cVL39UwmMXgU3kiIB5/4yz4T6x
eXhyPz5Hfd3jdzRgCW14tcVHX8maCghqACIuYad66Z57xIxPwAenyeYd0xRdsqpeMpq18jOqS2zx
f2KhpYiwJo9ysXwI9Bl36625UrrAPcjEm6Qo/BPvvsCoqrKa4tRKUOh3empE2X+mhREFqZeTmYX9
QPjld36A0xxtgUngNWlVUi4c1oyZZ4ZF0KKN8RiIsgah25vHeOCthRgMM7bwrNkYzoxhEwToq21A
yTg+tWMAgLHFxAPsVDrGMoGgJUdE15/tZXemHpcmdFrMqUhHpqdQeQyHa1TGTxE8m576yjDP8/CP
t88cwgHlveEgzOQIfD7h6UHU443woL/A5f429MschnVnpB+lz7Kgmt1c63xdawP5H/KVZ3qsX70J
V85OM1SQfpQvxLZ6pJCjQREyjqHH8jAvX1R5/Tx+gATIloOW4t4ddUgNr4dz8k9mSzLiEI8zsWpZ
LqfDLZtGE/wkAzBP1HC/tsvw8bZXo8im5mEucpFyB3EpTsYFGbutI1dSHkeJMQ+OImOrDUTxcwoB
pBLn49LIaWoChWI/GxFwfikJwUadReAojlkHM5elwhALimQyuIYnzuQ4ROfJeF9H0255SBfPrOsA
zRkQMd241Samu4For4PL8ha96dIHPKHQoqO88m5sr8hpLH7ELPrTr5AbVV4wA+itB3Vm2GOo3hVW
Ccj3E9uvsDZT4XrZXvJTod6MmLxlFLEI20HXi/wb6Rbc6eLAMUGLH7yF8yqoIfRvL56aFS+04LJn
4fGscfbEYCa02a+HPX4O2M8E0tL9wJBtv8aoJP+jztPE0JbESRWA7vTJ7d+IFVOwI9tqZqU9gZbU
RvMZ2gxpTtmbnvZnBY9x2AvsztbbJ2CDU5z6+FjJQgX6PesCqfUT8NJGJhmoVY7y51i3kOoF/TjY
so++5JpWYTQBSQ4uK7a/SdgtAxgFGFQmilUsA5hUElRNY9rF8dbMZUzZ+ccxfWZemhIER4njXVAg
x6YH0hVVW/+xFE/2nxEUG/Y7FmEaQSwE4q0/0p4MMY+5nl+WIlKl4Ajhj9Ok7AAYUNen0b5y3G1y
VMhG7GuVxcLp2cl+K2VZtGNh+KAt7rVI1VvkUB3H1t64/POt/464iyU3d0WPZKvyDiCIU09D1b68
F+7KninPGm/7SOEHp36ALRj7cWSwXFtJhdKpMpYtqbyauuV3rm+bbLQyOb4jgQny4qzZIUWYeaY6
VUypT8DdVDlF5k1Y+/18p17atRX6ohKp2wkCDnrFSkyGV2W2bb57sc3moYHgVMHHbCuP920+Jnnt
aGOvNcx4psutdfljShScTwr8IkrQrsmVn8D9RkC+1ASXxLvNWjKjy+3KnOGNnXu2nSH+tvp5fTA4
4JOcIoh7V02YqImP6dbvLepsRFQJt4wz9U3pY1GxsxCyae3EBb7J90ZqX6DH5Y/3tNPNonnDLbRZ
V5Y9ujHE1iwivfSvW1rJshaZoY7uS2CwPJqJTKuge2GWrj/fH55neMEPL4MhL8RvmlcRh6LxSDsp
AOiNQSv3Vqdv7yFRH3ZWuya5CZBZ0MmhWw7Wk+cTacF0xUbkHh4s2mif8kaQj4/yaqhgoLJcCf2t
ro04urVzR2Th1FW6ngt5Ox8OoG1vf1oBawDeGauFNtdIkKYg6AOq5G+Y6uvPynt+c46K+UeGFWQ5
2RWEqCl1UWIFLgmkvTJl5yoFk/4kVLjMSeL6BaWqjlE+ma5SBTploBasphXAMXxECOzqkLlAi4LP
VXE/DOvwUEwY5UsudpXj8ZO9zO+uDVt/v7tF09iptun39zwMNqUZjGMhLidg+Zikp7Uf8sYtYRfz
zR5AYCsS8oQuNhM/oc5OfYN18Qg5y+SLoazi4XCO4u9pxZJ4sdORxiBe7rJJjdiQ6o8DfwzcdvN+
akKU6Y9mmvFzDW/pdUfeZFsN1aaSmUrc4/WogZnoSlb74Oi9FFx6uDpoLIBTLLIditaGnJtoVswb
6qvDwWdwO223EJbYKGDFpVWnJvWb46UofEsfYfpdRDMesK/p7+sk3VBvJ+4JjJ5QmrFNk856mwZ7
OR2AaV2JVrTzEg2ygzbLlOkY94Xq/xo9AcqSYLgdgrYyB3PhohwFp5iYmudT78zXHsFvHTzd3F59
GcEoPrOzZtTjTgJWXCE6gVudnG3YnNjPFjvK4GWuaEejhbHYvf7OHR2dxjn0yEM/fpvEVzCauhC2
OpKo+ymKkR1T0k40FFaDgb4Gm5rHhmUdiDvkhTo0fL1zXQj9yVVEDPKK6MbLp542CXNiArrQJ0x7
wNU+7YSG2IaSUp9QoFfW3LAm4+Aonj5UKX0RqdnVXwCuxjDdRFaB0WFKxbgSmmNupPWNJ8OahSNA
VRZBvOXM2VkFU9zcKQyGf2b47U4f4mhx2PtER1LeZnCi17UKKzYokb7S+V8ZKOK3Gx4jqWQT6PCP
XwsaGl3FC0dBQ8aULyK94GjFflSJ7qHotUvgwD/wMpLKG0PsTvKGbzvUx6OZKe09+zkHj8qAXnNa
02GbeeAsGeg9601rIV/qFUKJa9W5JxPfW1DXKlu/CGBxK0o/CZlQcyFzUMoWWUi3+QUidtLciXaN
PIC+8YziajTMDDMZCn3dpdKWQfBX3U+KQj99cMCzJXMFBiWpPFUVhprFtwDQFJazNtaw5DXx5w7E
2ZMHA1lUdwbJ9KDyzKlBRl41AuVmSCzidujBxBao7pnUZLxp/F3UBYE5JGD5gEshgtPmC2xm+Fjf
7tcs3KP5YesmmV+kkGe6sqfduC1VKm8m6dAEi7OVkBNGpLd2rnjZ4IdIQv6qTGkqlLR98md8Gzzx
oInRxCaUaXmDorwwZWTlg3+9IOsB9vK7uMiItBIGiylV1L3RY6W04lTsSA2SwX7Z3UMuONonqfjJ
uUCPDeRZXHCLrCDwcaxWS6qwotpGCtyI8M8kxRIUPQ3EV8TSL3Cv5wdChOmlqvi5RamanmHmJm2v
BfXMBwEay1iR1tSs2uCvTKPGxcki0Ijb2ye4wfAY2OeNsP0maW4R+rBt+f14VUm7Ot4I1M1kTwFj
Vi18T7Kb2ihhFwzkjU+bxADAArJBh4rbkAxsJNwR3Suuk/rvhxblqV18SGmTUXUTlgw2rIMo5XN/
yaeIOkcDvvWrwijBNYHNVbfpUWUq17A+fidreDFOGUuLZUW/1PJzv/Q4tp3czclWKNQTUrZ/oi/A
DdYUrV8mzSiApSZ3KxuMyt7wgiI05cxBvKzn9lMB6yx0xZb6eaRwj5CS/hOj8WtUCtnVgJ28v9BL
WGv+/dYW+45rgcjprsxUhKedVwz42CIRjyUuJim8Fo48aPC3QentsKFlMydFK/6cGhEbP+C2BSDj
uLCWwjRIat5UxttXvFVTm13Rit0WmsBUpgIn0r5DewkCHGNQZ0HvTJrFCHoa/Qo+hsM/JNZqmmLZ
pYc8qKEOoLAM1oMQMgLJnAMaN942we3XMJCn62iB+8aTd1ecjYjUSGYzcc6rusC84YnM6a4gzr3c
2edhWHbMsXQhaT8PF8b1wtW8rDogopg0eDqbwWvGFutjGUVpkUxf2Q7rKEjqM2wPecRIRfbXxw7u
uVIoFSzD70rONLInsMfmjThGKdqdqvfT/clyI/yja3NQTqhi66/xglZ+RM1FJDr43fXuKCoVS7rV
q0MXaDZwoJWRnTHsnfhFFw05jAcP0ZQtFwwSIdIGNeijM6MDEinLhPcPzMSU5O6pzFdyZT87F/KL
iF2Q+ojA6TpMK75kJthnIfNWs7/+3p2ZSYm9MTKP6fJggBIjy4SHLLn8DSlBC7MQ1qXx30RcY/eu
g0NLb1AArL/TWuA2Dq8cwr/VYrfRiLdzfaEOfuCsTuvxlImCoP5KK9CDIfAONJsl7PNTdk3DXEhk
RtuMz8Lc6zKDmdcVsuOpfGKHmu2CMvslWE7j+j8wQ8cy8RvXUVu069l+jHxcPIOSVU0gyGJmB3NS
Dut/3uzvOkCgDh2gHdIFA1dtVTOQRRQk3gbl5DnOcJIVS7Pv05uGFRbXYwT7P4WqpNsCTTILHObN
aBtEnF9DuCIs2dYgxeoLkWdN/GDuXaY3B80oaUu8vVSTd5yiqtPaY5ZfKCmCC7KgS4VSZGpDVR3z
B2M23nY+Ytb805p/nNcU90HqtQDEn/qhH9sxXay7TtBfmOyRfKuFsj5O9VnzLHilNkQ9C/535AAe
EyW94nNXldLixVqCktmPp3pF2LU9w7PBYu5kdRq4KarIhasKsEaaKr9zvgQ92TM/NZy7oqOi4blh
WkjjaH0xawcmX298FReSt5xPQ2oFrnkVtMNJaM3gflqxrlZ2jCcrYzE2Y+58P2glJyUTkiIJF4er
hJpiCgF2jlqccRftl7snzThplDD/+6RVb+GfRUDRW/5Im2sMsuJ1QE9rQ5ChvV1Q00/+BLMgw08S
68hHe8x9ZvmZSPdD2ZVQz27odUWgiOm5IcVOrRrVREqey/uiXIW76bWmRFivyGYiF3KPmVktopft
BRhRY1OqtcNYn4sc+GNie9iYWHUKJl7e5nYx6S+dXXv/EWVslUDPpfW3v/jpGRTczS4Wn6kVOSd7
QFo5xB6YD+p1t/wgdFRcNzy7Y/DxtZ83BrfBqQ+QGD2ya87RfOS4f1RUXE+wa4aEYyTIrZs2blqT
oj1aEFVYLZzl0vRDzjkR2yuYBItbzsWivufm2LChnfkoLkAxZRJ0rrAGqisq7GjZCuDujDasPvGG
dGuZg055I53vuwITU5GsgQ2C6/CbxA8Fxocz1UoDVZ0eJhBry0YaqyTwXrJPF1HSDU7KXj5EvM8k
EDmc2z/QFGFZsFdPDsCJbFiJ4J4WIuAzoKrHJvXsyZ79AGPeUfiERL2TLXktCGvkihPeVN55y3Nb
eytzb3/0Nnb42pt7oaIEjjHEstf75RxbGm2XRxfEi7LYBzLnViXZma/nDRaJgLdoRIG3fOGMPUkP
UCj7xBOH7mWTBkOXyczcDtlWci1H6XPSXqT6mnBWpK2lKDvMyWckn4UPQI8RQRBBSFaZWQCpGjzb
E9yqCcrCeHt9+OQ0UwFyHObBBrJgkZyUA64ErHf02TyjbG9mONgEbkkzAffdORpTAnJK88YsdUhQ
9tfm6+U9DFtTn9QE9KRO0RA8flJ/hsP8ZoA2jIx84UZZtKyGgRZVI9Uuz4WDiDOdlXVB4ybqehlb
TaPgRWliHRiTrwpKtoM64TRLl3FluSpzMTlpFob9gPrB+C1CqUdEGN77nELwgOB8Fn2+dNe13Ji7
lN4ZJcaeDhnl6aPZ0Z4uj3As3LKVKeFcyJG/2TxCZYrBeXeH7fIcDtr9P2Ziv4p2hyms3rRu+kGv
OC77BzZqmXx9dLWjiEY0xEf5MPhICc6XbeS29d3Enuin1h3umzKQcc681QItHkXP1AY4dLevg/rF
NqSoJ149zs9u6ZvQOZh7Sz7hoMnEJ2STKXFPHt90BUti/5+4rpgS2z0LQ5v6ngT65Q+RKzN3eRGg
PeYctfECg24KWtdEFvdpXP1TgfvmqKkdKbHE2igL3TaJLLYhsJLpbePcNbPZyRZoBprmiR27jVxk
aOcOcZHRcZSgUSbGwDJI3H61oN3VUCqTB9KW2blBL8w/oxRSnOzn0VHG12OpVThMFc91OH2sUFhD
9uSLY4om4E9SfBfYkCvLxK7a4EYdKbdt0l7OejtC+Gg2ekMaKgZQmoANGgiD5nn8D6vdzUmozWiR
0Z5ZR4MAjzw495sX8AA5dZnazFnvQ4WbLyE9VxEQbeA0S8gbnpLVDwBhPRMfoL4zBxcKa5vHW0yW
b5UwkdRZqATU0qKzrA48QPvM8jnZwSZtsr/tl2epXAek5+FG/LJ/nKwSaEPrFmlPxOcfk2l0097a
FQ8Cr/17bxy1mP5JLIGoRxzzYyoDx1O5k0R3xTi85X4ODPFeYBQzVg9hbIt7YvZwbFiVo+7gooS5
daBBFHxKYoNSEZiU4c+IM79zsmt9xk5MMkDykcL3oEgS/BD1CIvjrzyUA8o7bZKSN94dBIo/ecQc
KN/wklxlw01slbikCEaJbVnHlFf7tHecfBFIwFjlMZXLmfRRZHN+bMqnIbKIt6kUmqpPLJ332fLG
HfkhNzxfJWMu1peKDAxFQysdfVBlOQsLp9qZWWwFwu8ynYE/f7lhq8LRFw28O6VTQXAsPPy3Mggj
LALb0pXUY2/6pzEZ9aCsGNjZQqUtUT7aZyjqPNVXVErxeBjFQUxtNgYZCexKD2VwpC65/JKTaW47
ofiRjRFGfQ71ykTBoLxvpjweuVVpvm8pKRetql2X5Oc35rXOQLRi6HXzlD8XFSOmaewwEUpblAal
acg5CuI+RPj6TiVImV2ui5795drAoyxNPKGMsEphGKEa2q3JTZUqRA6Ix1Ci2aadnrtDg3smSBbK
hBWTvFG8btwdkveLmDms/01M/dL/5YYmCD0QTeRg74Q09/EyUIssibamvvilZWFiC6k41DxiRp2o
O6KmuSQLr70XWeVnaST/E+2Qf2TzPX2+bNm0UxKkXip6VQx+rTez4Iswk/jsTLWb6B6J3qciUfwj
HVPB/lLjbQzfA6B6tgssaeW9Bz2glZuGi9U5dJQPLWSvO0ElxLnEew2o2/HHDeqm6yveSxLTVrvW
KnOMST/jklVLW3Xv+VxfColWkhuYmA51cWOaL0pQ79s+a0JMSQxemIKp5rWVcReRR4v415+XNSZA
wjMZkYjcDhF4N5/8OJfYqKVGDxjIrifIe2AP62J/c4yOLavQNG4t24q9QuYbDtPGNxQvsGi33nD/
4+DK/Y4EWd08kk3+7ykgKVcXGWg3xOD7nnuQetkWo6u8AOZLZAoSs6O1pwNTFdFrpYExaIfEni92
vBI1kT+3Uv7yObJe+80FwzIA+hXGofhZEDYqKlmgGAMX0cA1ybUnYlwpyvK5kQVKaqUL8NGLVv8K
YnomXjMpAUdO0SDZkA3Fjsc1Cy0tg7UmUBxdggPDawgZdJGRrgNuCchKiiJ4BFUZccVE73ID9KIF
w9GblTrvasIutaftTyMNcpSBvn20Eut2Ha1iD9ZwuOr82zNaGUxEb28Llap/cO3t+pLudinXA1Zc
e5XF8LiIl94JngGGoCumrWQMHEvy+UeuwfGAaakRMxwY9zNcUqYDWjcGP6BfZcSzyqopWhIz8jFD
a+bixAWBwOvEbgNRFdwdyCV+RnOa//gh+ARrwbNbo2njulBg9pTlNHBn54hRwCA6DqMrtarTTQLl
c5nE0RQi5tIYOFskvZU1hsyi/6VSBruq5NUHoza6lXbRlrmNTQfno7hyQdvIK/tm/DUaMvr6S3OU
QpJ848UMQP5U09bwpR7Hcr7ed1mZe57qfKeoKGMSRSEXGBq1w3arUx+sKMc+FUOyb+O/wrIZFI1g
p6+NoWPn7OtU5tYRcLKQre5iULYSBxwWT0wj68aGFYU64WbBCpKthgnMQdRw0s72m8/B6yK3TkvO
XcslNO4DokFV8kcPDZYxxz4emtZhaYZlhsy23LMRLjyQ+2e+wFa1GVEDUfITI7/IlbkfohF87/MW
KXasJiOkcqlOJjLssGbfV1CkTDtwIhMA7eMzUMRhPJVGLL4fIWpkmxO8aPQSMwBOpw63cfLY7fdb
NTc9mTu7Xqu0ZoxAQoUmDc401AkbuYsyIZ+QIXwKIlwQO9JhR1IGpc6J3BiKOSXreVW9VpDN9Lqh
5o6Z5JODsyr+bJH9cGsGeCQ+xJpQh7FzKLDEiN773aNe8FOHwOx+ToLeO5/LWs3tJu4issC7zLa8
81Q+R3nWULmFlB+S0VPsrkK/LAiWe2Z4F69kJ469irc8roBES9xCQS9kUwOZScZZg8gJI0SmMax/
u3XeO2vR92JHrrRUrD7DnHBgZhYU94/wgSBI/DIaStsiwM4hYvz9zGTNwK0RKpYGv3jjCZDwtsGS
Fqs9nQ4Wez+IIupnuHtdCRFBbbZVWO4W+HKVnEjApIM7sB2jPplxiuOVICKg0mJu5RaZMYgBx9KL
/FhPP7d/vSqVNuX3cLQ9oOZAM8O+ZjtTPbafP6UPvplnKOpihie+uiCRX2Nb87erC/Yj/0EcMfT3
q0rE3qXoPq+V0WjYdIhdZE0jc2BI2SAGfIZdUxpyIvP7WZiRWdl1N+WTfA2/315G8WHcmxFNH4GJ
vzn6yQzzoBBGxqx4XrZeQOqdLVABQEscC32yPIkCEY/Hn4X9XjgvEB/Gxg/unDqJvbeVZJxr9VrG
gZ92LglyXdv3n9fGuc64yy8uvGyZsbWL4Uys1XNfgZXTFeosXHajE1wMVrNRLYlG+LS4cwXBB4lt
z1gu/bQWAe1iMRz+XFC/D0IN4uOE/cWw7Kf0uK4VL7wCBW4g4ufYCusrFZbNyjpukmv1t5kKIfy3
gyVsekmnTsrFOPStJoUXOLqrrf0+sMflD4tEah+9FJvqLYHwywXZj6GFZztNztIJKjcuI58syOMB
BxNuTpBPC9AlGkWFGOM8tVXmDuhoAR91Pr+W8Jt8T1/zH28aU10D5tMA8ndwBfO5enUXf13J9Tq8
QZa3sRNNNZIkyJSmXzoUKpnD1VQHKSfrtU/gMomFHary0rBYjv1bnZGjBRRXUIgiYo4oEAGR/9zU
/Kcl/RblaDKIOe1yhLjkAOgp1n9KrZyTkJynghqmZX0H/BXP+ofz0BQI6Ce4iXfIcxQZARIxVVzQ
xBxGq0EmthS764/yhVaL5daSF36MjYLLFPnyqA2BHrLWnP8N145dvpvbdmcuzirOWSZBB297Ppw9
sgQxy/ZYC01u+aerqpbzGwbWXckTf6SAiYgZBfhq2vyqf/MXlD6BQj4EaaY83ezsECPi95aPgbxp
M9z5ZIZj/YI5bwtUpGrKARbgfZAV6gzWVWHn/8QsswmD34Uv6AZkZnF4Ls9kJsrWmArdk0dDxQQ6
6385XSbMaNdLFFt3M2r2ublAnk4iXuhQY48b01pB2mUNn2LwngJKzT2sxN2/DgOkU7gqLaNrCv7c
B9m6Udw3xIAp909EmLGDwV0b8MedIVwWuL3PYknE4D29TSkUxfXlWSOa5rCqkV5EHVSZ0teJ2C/D
05cGCn89+YpaTUb1+GpHgP0RT/XhfQcycZE7XkstyKanOp12qU7qVrvjttXh4er3d9FVgCeZhE/K
ph1xb3Hp+F00Eo51HN4B5hZbQZl5TMlDvFoAsec2Q5R3KaojOc55V95CV2Nl/edzzUoRFzgxSos2
JRrof1SycEGIcwyoAtt9GKl158mdfhDfQwt6A9j0GOduEPHJsr2IKb4w2V5RMejv+KFsQbKwGLyO
RFE9ekD33mTrr5+UBBxy676qRVYTxveiUSme0CC0xmZvnN/85eWH/xV4aUXoKbDf3ZbnEafSFM/q
f6qAMB0qhWE8atLaVVQpv8TCAf/KXo4dxo5/5qJ2lpyJBPCjkoszldejE7VB8Tyg36E+AQYPKk9P
MBhIhfGh1UIpH6iCL8k8EvCAaSjrw+kwtWYalvCdQBxr3nYWg24mFyt6oinwzZPyEA1aSu9ERZUY
ow/Jrcz90P8upBPxOc2I6pDcl1KE1SWpf1evdnCYlX+EMGtAtZlTUl6skVCbwDNI6ARG0JLiKDiu
yrHcBoEurlLfzJlycfx7ioeLMH+5y3g6UuVDxSh5FOGwErixcn5wNMolWO66aTnbardPaSTeTwR6
SbAngh6BwofpEMT9YteXmpM242G43Gzf4q7tUEOV0WkLA7gC1ifbTtfDsGCTEING1C0ZdbJSH96B
BwltK24qX5MW7ZHC89Io81OvYZocdASWO56wgWK/PLkrnZQ86LWT2LbejALiQj/VLHUpRd5+Lrt4
VDe5NTNN6bVyIF9mFVQWUCX/DnOxXd1qCcsTqrAxoAcFgyC4jVkkt67hr5C9IEZuIrD+yizsyRkl
h2019+Beup30m63b7J5NRPlwOSf8cl2QT/NuJCi5QA2WtNOVL6kQWu/Vkm6+WzqCUvyB3kkyviix
heY+jMS2aDAnL1T0BdJ+wcb8Rklat2ugcpkQaLNe39u2amTSrDnF69mAzGVqYQb6SESqIFAAIqkV
L/kEzmO4gYlJ4ty+ja6hfHBzGBpNJ0wrlYMwTfEMMqAYl/clJ5AlNJ/LRLdYfTpa+M8LUsujBflW
pVzINuqZNnb1iOSVV2vWaVa9GrwTyS1Kl2qEz8p1s5Qb4KhJVsOYMTmr0LbHvKc+smzdqJGYFNVn
9dHQiAbIX/oz+KE7gdrzhi0wtGW+EsPmLTzCbwHM9KNvSvV4OeQQ0vTGB8XvsXDi8ufGajO/cjb0
qJAKI2o9sr5cjk3X6AcmC6RASHHa4KyX6Zr2VqT3Sl/I4CHvPBVfKPqycEgDdZc9J9CZHLq+5V2E
BexbB/nQ/wCKDxGrPgpPTcFUqCPcLYJPggnN47x0s97zOHJ6/+wq4JZK87YkMi4vKfWU0reDkfqp
TjVbYQVCRYXxrniUXMQtRmbmQUA3+gWvfLdlaxr87A8EbSaTF8kgkC6/kHrz0C9XXj1x6+UkDtAC
BqY++HIBdnulPoM3P8atylxH6emW+Am/Myes0wDsPUGSCZHne/aik0NX2F7VmWnOp/BEMqe1pmVj
odhrT+w/EPMuWXTMUdVZ1ERLSFG0pEAL/QhIIAZMluwJeTgok/c6mqGLTpR52w+lDOJ0v9SS93jT
b6m0n98fh3P/pgC9l4xTBr9S1LK06PWkqJnyw3+UsQ5ijuXEZMvOU5afLLhDps17nUPIc528b2/L
FXnVzF5rugAEoXsL7FlDoM9iMonlSBubs7wu88hjqKc4TeTP5Q6PF5a0F65iY71o5w5dqiPSJq88
kYqSG5aENjoadzrEpT3cX3MaQWSDOONcVrA0gVc3n+1407ONJTEU2ZUbVN1wnuXOunaWrzmqZ/CU
Vn7TXeI48bgYU8cR/S7J7E6ePeKZz9LsCXdlsrf1QPeUA6e44SXlhB9xrVSPH/gLD07MmMMr60wj
kuD2GH8T0sAQ2kvIwNrjvruekzpyjo6h3py4r6dZHRpDsX2pet96Pa/y4UKn+HLZnjoiN2zt7PoC
MuWBXjqTa8YhBEOvmmKTdwpfurLDmRCsQ/CO9mqtCXvlT2P/EW1cE6mFcOY6u9Kn7fUxr5yKYu45
30NIFRaA2/wZW6+Jt6dJAI6JgCuTV5gIsGUZSF4SNvxWIqAW5fjCTQ34eFU2JK4sWkXLzEvDOmEM
E3Wci+ZrVoAjJ3YEgcZMhGkI1E5d2lGu1jx+4ohVASTTWZ8X8jn0YA1WdIaqMrvCKfvL6dsJ3Mty
0GgvJVEX8YcHxzNFg1lk772vqEzUvwA9M4JQgFud4PGvNQWoBVno9TbFN9+6f7ffNQK1tEovH8Je
+zGNF1t6USxvog5pcSK7q7nsUo+EMdheNMn6jbZHVXd/W6PEPuItMiqEi4tcUc+Aq/g18fFMmlFx
5Y9/ZZYhpDNK6olypvjwhrxXP4T+BkU1V0Il7ow4penfmnTKD0vbPOkBdeu1KUCE+u4tyxFJsbLu
D0CeXzkRFK5IWImjZ9I3tdWkkfp2M5jfjHks6fJj8SnDdgWw+8+X751SJL1yt+Isd8EVFQ0d5uHU
elAgHukTfEF/K8MJRF9LxwILHDW209boe9SFhsmefC+rIRZRrvlr9Nv72m2Jy8/TjFtHgXJho/o8
eMAwUqQ7FRjw5CwIn3vsB77ZyY0QX9z+gohe8RBTsaTszVJESCk5VkCqxBzOKx7TaGT7Z+DgHWGL
smK8sEaiXeeRlMfdyG0vwsjt4EhutiRAipEEn7D72+24nnyHPgcE1uWhBpvuOxEYPULAELv8sExU
fTAgWtSXNDF0hWfBkvjCAeU1d5l9ptuMqKadGe9aUHI5wV53XeBcy0Y4JXk+O+CJI1svBJ5LQ/VD
P7S3xeZx7gsMJuKDVkci6BqdZ2Wm+Jdse4JmrmO7n9IFYHd8grD8hCAlJDnYVdWtydMlXvETc2PP
6qLslLTfFKBZWodecW6i7fByGG7X1LLeywnCeB6KlwGgvUT8I3ju1PCgd4h8vrCGTaAhjdqUIyHC
bm6sRDKS1VEATZrxnjFrN2Xk/9Xo09DLf7/4Blsea9+Ow/oGhA3CvYlMoutdFucUo04txJtjRRqr
rx81S3lTtmXPfyB+D9/r/IxebIPHr0pkZiKZVFb3uPZzc3Jrh7UsQH56dsWn5dpYFdcPyAe1Bzt3
nQlXcA9BM/6yA9/uxY8M52DmrZNh+pekD/3lupX/XCvo4S4BDzaSU2M8b8RRouaSfBKD/qfuZ1uj
ZZoYS5xEmei5+jTKlB+AnU0pAG3gLK9zNefbYRPQ6VPDkvzzhpUe6WVtW/Y0H38sqSA2v3xsm3F7
GPdwhteJb3rj5DqZ+tPE9WpgeyFz0v31K2++85Xd+wI+K4WDhIAtUXX6qkuAdyQAjE16SGOB9sDi
8SWEWONMQNMrxzVh/AbqkZCIzDn9qYUmXwBR/gNiiy9+WE/TUQJ2AgX68YFWVrDeQidAxDG98vhq
wPqjoZHgQiXjC+aC4jKLMgiRfDG+EqDqWiAeZP+lmwv7vZaePSs5f1VjBRFNiiDWtIXc2YSrE/Ev
faBE26acacSNwZCL5yT+rn0Gbr9Vls3cUlZ8rG0PxBRBNkNd5YKjcuqCXL3CeMSdnf/N/kP7F2Sg
JuJLwWLp5d7DBbCLv1wHJOqbBjy33sc6h3NNEbiZK98WxN1xb1XQy9TBbLI4n09LIBbHZcYdJbcj
g3GFy+3y3/C5YaKCZ+qGCNhsCoV3i6cXUzNYbihAd0PaN9elOnBn0wAaLtQ5k3840kxuPCTGqCWX
pRgSkVNWj5ed6z9193CCKAe8+pH81BmvUkqnvp/OK59wHnh/g05o0O9Y6bEuLDADRAcJ8Uph6RBF
FUg3RHsrvRoUQqlDAt2W6Zdeixzo8BhGZoDFRFmHWQxrm+S7401QZE+Ktk4g2PwxGUqz0Axy/Iqd
vfn0Wk7NrMOfi5Hxeb2RvpFRHmGvwCTvzy+gjVcWmvnU6y8WcbuphaETQ8x/AAAMsVsWIB0lK9tK
VOjbaZu3VWAY5VZyimon11VvauWo6mKffioVQQc+vrFgfrhIEMkO96NXcRJ46vFiTbX8H5E1ACt7
vAT7Klc0m2zuNnQuw21YhgslUt5wv8L4jYwnoDn6kY3WLq2TMtEDtttM1VRrlJXaS4oMT9o/uXKg
leK7hZ9r2/uP/Hk5+a/mDVTxAar+pwIcFWxKvd+fxj5J+Q3hLltMkZu8fKRSeIJlEslsXgzwzXrI
tS1Kfe+a+jWOZXA2lfK5LL13LRjXWj2OrGGuYjetSqdTUs92Qb8kw0zElfPnhqoJGtDPIjNlxMS2
Epek/1Aksta6NXUrmH3+GgNfy4JTkb8xO5aQMTuq2ikZCNIdp0DtIsmyEErKm8BE7qGyzJL6L/22
89QcRtt/H6Kk7/8y7DmSCxL8m3mdXzxwl7SkukYSr5hgGlEdlXKuNFOGyTbT/lLjdS95fMob87zu
J84qzvDWCvIszfDuyrlbxi7oirfYmTg+IfGiWbj1Q6QH7UI9sph/Ml40j2Z/3imS6YnLv0CpWpO1
S7NmfHuXqaSnL9wRodiPqNSl8+cdqouLDVqGgfSyu4VcpfLYY/4+2Ky4HTzAjktgexXgHZwcadup
19KJXVc0AygG/PhnPAkdzCAiprKg2xNQOjW99bGyCfrqsM99OYtCf089Nfx7aRBQXnkJFzSZONMF
DYzTz8opjf12lgOG6ScWuY4/hUcKlbBT67iUlScsmhNeanFScp0xzPMGfJdmWJ2mpUn1aqPhDIua
D4Ahf9fgXY8bjPGlvylSoQ/38Yi6ae7PQX/LgbXiBXS5ZYoOWAkianxqmUDCIPUdfbIGuITJEfCx
xNECN5i50pTN4eFaQ/gIko3EMOqIBttGXWo1sjVN0BqM2hyOZivmpKqXV/hXYhtK6uDxRtspcfk6
/A78IRDYkV0sJBT4cxYpSdF2U9x72JTbcAbOjIcvxScgAOPWyw7Uepm0itLoM3cbhLDSNQ4gs4vf
279kGjt+JbnKu+3UL5HmjfysjV1MhrW6ael1iy7cx8PzsFl+P/mFZcUapwDowEh6qMXPjxmgyAie
afw+cVgNBzv4euVEnrLIv6hD0H4HjA3Q/PCQVvXhnprmxg5ZR9KJjqDohJ4bsQwlvCNeAjQWlF1i
Xbv8JXtjHnG2UjqnQU5NmqaUUY5KF3a4Y6DlE83c9FhntPm5JCcTJjl6ZV7S6H0CtHunY5BisKde
GFoqh4V1ClPqOez5mZ8JvkONEBVKtLeM3bFB+z6jDPd3fEOxoN4NqrIT6693rf9R2vBzc59/7TCW
lifJQOM5yQbNJdv2QvHjH0LcurcVWxMxNhQnNTwC6JLIKlajH0KN5Cj7ATx7K/deP1w3ElvhDeRg
A82f6XNMFnsA/khpZJBAeCOQ7aNeqn2xtEI8t7SqLR51zbf4Uwm5I7coUrOv8QoBMHAd2SbOcgUi
PBsbS256YTQ55rjFQVU/jz0McyAqs+hpUFopidTr4ztLAeDDJn6WOeJ/3UQaxX4M5PEwDOb6CJQo
o2Vfun/RZUH4mivKPz6d5t58lOAt9Q0rXOxUj1adMnlBHH81myPS3mN4nQrEURNikAMYOFxl2s59
fqyH9HPG8En9O7leCn28/xndmgHm3TpsamoDKgjQvtIbBb+Ff5lmc0nt5HjGpMIwdi0Xkp7X5UQA
H6Whd4dzFhPCe5wlb2yz0LEJAs2l8ubHQt9i1JKDaYtg2b5p69vsbtLSi/NGdKpdlNung50+6doX
+DVyRnemC8pzIqxQ4dN86zm0av3fP8AEhLPNXQeuBUDqJhDFJvBE7VRKomASdLUCvlgqPchCay4g
O/7Iq+4Gqn6OFy9BCuRN1NxlDtd7CdnicyREOhwkSoV84JhZlOs2FDy4xTivt9FIjYTk+1LkWtHC
kI6VKBxiLSc2WuGdetcSQirE186P1KU7waigq9J7papuJ1RmK0hOf3cN4iQwwBokiIVpxtULmuNb
X0JzS9DJ4MIBL7WiBRwWFCfDH2cuJ48U1MiLKzvC46H36EP0qWkF31kG6i9UmQLL/esyKpV3tT6Y
rhyWSdhqv76eghGGIPMwVuvToFcnuJ9mYXD2NYAns5E+g3pFLSG7T3AI6yAkysCPb6KZq6Mx/ku3
dmqc4awGkYl3kA//IhjfzNHgVszdVxRtC704akNgAxkAx/n5GUf1EDEhxwGAR7GvyN2nk1cCg0ih
L8rLiw+mmY8oUDuqTGMtyDIN6gG/QHe7b+vgESM3M7s+vYMaZiGtN8PINBDROfpmggud1foLxRh6
vEsA+IYwQppp80D7zSvxtLg3dW7goqmUPFeD0UQVO5Xo9+RSLKNOVDOG1p3Jr+YBAYJScKV1aPNw
LeCk4RkixuXbd1bq+SHUW14lixlUTAs4WXFg46MkXx9jBla+OhDYiH6Ovmc9EZOAdw+H5XHpT+HO
egwqkNja+dfSjaOPLFNEL8CfJfuYigtUgGTjOgEC3MeJj20hqfsyzXK8MY/kf1HRu9/rk/O8f3vc
RPlyHoW3VpjgTgqan7zR0P85dSaHGgI1mtvK7F7CnDXc3IzNDclozrFE38ctg7cTosQTzN3r/DJh
oW+indyr23n2YiaR32NApa3RQrpWAJ6wfkYbT6122OWy6UY73CMLoRUWBpgXsRYwXHSegMVybTQ8
R95yzirykQceNggGWnA+Z7/NAadzPL1VSqs2vETBkWaBQ3gjTU7j9A57gURfhCPCkkAJZP96w8Yz
GRrpS9ubJUqn6cyzxnFlsAralJA1gHRJTRVGM37VJbNe46sKjGEoHopUMXcyoUGU5A3GXMOc6FTo
nnaYT6psL+mXdl3ZI0cNpJ5DOSIEgxciEpOLc+4jdeZjnFaARsU+Hws6Xc7349WFqEpvSxvdYQb4
AQByeWSaZe5VNMSxz0S/GSy44C6BY9c5du6QwuoE8QtUX4ihUpKX+IiHQ0JW+B8tGmBS/eyxS9st
4+c+jg9DN6TBgqwSLY3jsNICeteiGFusA58nj5XML3N6RgxGdhpUTnuRnPmTFoafUGuy+AxP3n4U
aKVx260jO/HAm0GHOQhNgujfaMHKNkTgbCuRQSJaehJIvfpAkG8ztmPff/c2uhOsJ0GZH/Awtj1J
Oi6F5jiwCMRg93Yh0sTSneI87q1wayfbcGZHUXOtYXbcl7Moq0H+8ybhWICjEfvneY94QV/hhin/
FvKTeiTK0Is15eQXOupMdSSZ6BnnDXlcB98hhHYzmCZXbP5jCRfIQZTiyqSoIQ7460L8Fg5upMVX
WOmoc58ycDkAg304qJ34MJalXYu0CcaqVwltUmupUuahpL2KAw/yIe61C1YouU9tVWqkEdTa01li
DVahL/WFgyemAgIRxLzS9QXqC40P2hWYhbrf+q4mxdddMQ2+rqdESVzugdSRQzNDVrKtZoJqqHBi
apGQv1egOMqf+9wLYXRYocn72aRSyOZpj9JtG9WEczn4EzEDbvDFbI1I/kRm8DkyFJPogokzhZ29
VOp6/2KEFindl+XKiQRrzHm68Qaz9GfP+e5d7tzKVyuWr2XuJSnIMcEHRAdCbiOZ9MzqpMMRFRlx
I6l8pA4B/pMbXpnCw5eh2I/k+iYhEWKa/k/iwUua1uwCXP6kI/ljE+HnSRXYGSEMrg2DVXRfkhYc
Avwbrg1x4PXZ+Er28WkU6J00gZ/Cm8uQXd1Tyf9bD7usgAzgtTBc26pIAeasnE4NGl5qGonEOAQw
PMQRRCm0I8HgxBBZ6tOOCpTe/wUs/fvqZ0nmE9/02kqBmg4bQl6fNqd7YeupydHiY8qudTcj/8S5
yFC+Rj1/PJHD/y0+XclZpKsCNTi2ymmsfhV/8G1eP840AlC5cx27CBY9JDgHVfVSTvPI3tev49SU
n9VIhrM4Lx6VXgkIAC0+ZOo6ILX3eodeJAIrWefbkkOa1Jp3UVo3I7hyw5QhqfisqaMP+WRi8fTY
OUsTHsKPlnBj3OTaazAfe2C4uC5CULy6wRCdNmvLl/YiU6xmAkiaZBgFfX/3y0esiJpwchVlpA0r
MEKbrQcjkiYIzc2hEJXFOQSPMamo36XIzNuddetWF7AbA/weLbDaBWKveNvkSRG/UyHyOVrJahWM
2fT4Ouw24Pbww4Bpd9h4sD9PTtd8XInQDRNhzNw5+sh7Hlrkd2rXtpESQ4Nwb5yjlMKisyPhamvW
06NW2m+DNtlzEMFoty3Yr/ewd4JbpNCzJrazEe0mCqGm09pxUEdDqyo4TOgLCT8mytQiDCSe39YO
JjaI0zsmu8nhgzuNxpENZp/qtNPyz26d3eiMRXgFFGwFJkJWASjg69jHqRzmlwsS7SsTGBY2CsfG
QErLfQth9yC8NPAG1Qcn6Glox9hTlPHiwnJD2gh8vjr/5qzzU2rnoKBNbFC30SwDD+rA3x+aJYPn
/522/FBRW5swpfHl4EsqIDXANC8WxZ9zxuMJf6PENZVpQnpKAv07kfybbkLruliZ9rWecgUwfda9
xnUb7dyze/74zV9z3EgSxgjOMNnFpS45r3ymkyVYvM/3pjPs2ca5+ycN58WfJNzC4AFhJDyBYnha
3FFqCv1jRhpLr3bLXcW4O3JMaaNDfsCiffU9VLlPmi6o9YQ8GpAzoDnHUfXqC78tlttTuzKS4Y/l
3ds/4D/MEcRVrtcQDxa4rprEAKw6hF7b+kvPc+lNFC3BJaR6HdNPPV/Cra8qA9XpXZQl6Pa7RykV
On8Palq3ljRKWRhPiBedIF+LOPJoUyh0dwNDrtd62psC9cOChV+Xv/Xf8vCEfngPplOBtZacgaJE
EDk86+CvcgMDAeAiTtyZwPsEHHtnMrsTxO85AlFWa0Wi5xBMz5/Sr1IpSjP9tPiVsevMZ6ijuOHR
mZq1gVDI4dgitNaP/TAoL3FNSYsSEq1ctjg3o9Nl2oXtxLrGV1u723sZxHGxwb4ZjFxvXGoyybih
o3TrXKzaqbmlVl8Iya+3NcYJQp17Il8vMa5jRsOxfOnuwR79tTVVuXm8MRuPHbwyRW+OpSUfV/HV
sdbTaU5ltUaUWxIxIdbYLAfOof+1c9sYJCEi0z57ScxIm6V4lBxN92dm3qI0lJgTPtIwkEul6MhI
hrltSOeX0qkoDkKjpo2ezguIpn/EfTD3Bq8cBTvKsoLbLG2s3tS3d3V9iqXiAfj3akZBBJamSYIZ
+lOwKKMfeaJjfTPMb9PDBV5zhpZcQmWJ44mIfLngLoLK8QTeGFVB59dg0ESUTIk1IMle0M1Eyxsy
DaBkpvDgi4Unwhlj6t4YNSfCW7E6ntP4Xv5198d4PT6Y/2sEA1yJoXNT7PlY6q05AMBia90oOTD1
qmIzu0sS03+Ez6JUheSmWb8DXp9W4Ta3191LLeYHey3dQW5Cn18qnOH0f+aTeSbTWbsKvWN+fZXS
w8tc8YjcuZAUm00RJstTKdLIuDG2lrqoh2YK+5mMqAO7KHoDZlDuDduTLRAx+qnEoUbU/g/7QdwZ
NT1izXT191yCk16UEJDiysvcrZ6om28fVzxvn2PLVwWQO9rTPHcugCCUdId8x+WT94pNcLv1WOsY
G5fyzEtu/ZdIyM5VUB83xxIDebNNtd0QkIQiAmB8bRt4YrBBqBQQHGPlVBwuj2YGiQcuJPUHGyOA
sPY0Rot+LuivnkA3YuKSdw5RC+G+yoY0POq6E0U/Gptst+Tl4wUZScn8bEGrpMioHNjpu9GomLoj
sp/wacD8NfYgm+2ZWY7K61KKdAHq3nDRXOJGPgux3wnTZ/xzZ2nD2OyqY6ue/BdN5OeFsRRQ0skv
lnXNwiaxJcsNMw5EXyezMIhsDBUetHSOqfTiE6gSHRM32hiuXdmXk18fJG8xvURLE817hKigXAZ2
App4lkNxQETqYqBM+KPXwlyPfNoI2ZURb79Uy/A8pDmnUM4jYM8Ipm7Mw+bZOuU5a3B3H9MgjG4v
wBSQ6eiF2iskyPgfReHfqnu8wZi2ybUA+MVUjA6+9Dx7EtX5RXdE/t4X9Llzkiy2i/ltg4yqejYH
j+uBMwqqCqZUbCDZ4W1Vb+ubGXbfLkPJ4sv+2s9mXAH3qAZ/W2FerUYMZaguXNk2JfqIPqcb/7c2
A/55ucoycz/3NbQrfGWP2XQ4qJjSL1PUduPYLqnZqVxoh7chFRMg5DvmPXNjF1v0tUkthD+chlvg
y+wxKDOblT+FzlNPj2EuSX9vnpvvw9Aw5h/mFsemUDS1gy6NsyS1+1OJwFJsHxlpRvcwbD77G7tg
9NyJP79UgR1bfb1QyEhf+yuZN+mV3jKQo3JVb5Lu4jq005tK7OXPMlCieW1k8lbl7YkbzoHoWuc4
PjfEpLmR52uFJc0+DOKwaRkmC6AP5hmPYNiOCew/d/XcVHqhGcObN3rOFLr5mSPQgeuSZPq0P0vh
Evqncj1yNZEvmo/f76HniXT3C/30Jm0HfU7dJN/efyDRvANeQ7WDPoalSCsNf6PEJCgfmL1VT/mb
Rgn2yoZrF2thfRIL7h+KCqht03gdTJ0Ly5t0zO8+HlXPRPyOnbSvHBXsj2XuLNOnWyK/neqpTl1e
LDigEuixIP4g8eVjJhUKH7TGoctzmrVUjyun4AGEsLT0CoNMjDZ4lfoMYwIptp47qGDHPcJjs1Ix
6VMe8FlRC+P6BlfgJVZcCgW0kuh7K1cFE053jpR3yJrZYQ0CjytcqCi73lUKYHQao9Poiv2QHBat
r/2DAL557M397iv00IKnkooDQbYl857itxSpr6C1S3Uvizw4CPxZumBjARvss9DWLJZdZyj3XanI
tlPPiax1Pzvzl3LzGJ4Zj7byWlhDpuv5Y7k0A1kyUvZbZqLeBz2eVs6wjviOY6qcEtomaJObDh7a
NCjRkY3f2RFEgAt3JvRKUzgiFeVUC4zhxEfvfqOZPgxM3nwLBRMwss+lwWLUGNu3UF19EoGZScXc
2jagAx7hVzPcqVrpoXnLRVJpNnZIOmWk7Cmfau08/bBZKLXZ2SwODnlBuhkcj9NUu4U5VZFoUdU9
xmAFTJZjWmpZ68yQ6lZPfWfZlUq+GD/lzTgNXBHf4bgqTOQq9fpQMwE/7S/uKqrzOps0OpJiLzyG
GnJ+qU+6PDXjxFFOxMDNnRQBLdegENCmYdiSLGMpsSD5/K0h+QL4pEAbxG989eqnoNG18+5LzZn1
5eH5/wq+eaLx/HtKnsv9vYY6Swgi8D4tl06Z28hGs6rMHDVtw6pVYjUNQ23vQY8G+t+HddymuCN8
QOjgbZIEqOGI0eQl2s1ncz+XXdK+qv+5fPl+xNxYbf6iuEiqr8aK+KV9gYq2ckfkOX60OQ/Vtls1
4sVXNHK/J0u44XBrxMAOFR98vZFm5JFKFTJX4Y8/1Spc3Df7FlLSrkQmV9KV0Rw11xAzD0PsAbxV
YmBTl62ZG9YMSfb9DGzLFarZsYdDJLCd57lYzZcvzB9W0H1o/bAI1pWLHEjVC/7Spcmer0rj/Ew2
8MHxymP34NslBeNHhKaDJig60FpQFag8IYQ1mPjktzhxxRLjLDLJ0OX/rnOWCh8yccN3CUFO9Cgv
OfRztoMuqVI+m5zjErH5OH/SrWNFe20zLx3DBAhlWh/06AfvUcyapNeoST16pVOl1yc+S346EQUc
qq4kU5ac3N0KBuJ+//0WUjfyn5TXqEcMTRW5D2JB0LmBOGErhGdiRx36WnBvcZW6bxhZRXiwn4aX
Pvd2Ydxu/Jqher9I8zQfpVyQIWIBKOJuSESKqvIj4vzo8XUIIX9v+9pFS4+wP/KwW/J5+dafw6Dg
OFcXXIEii5nE6QZie4sIk76JqbaXpKxBzanqp9GPVcdZROxcznwVymqntBagZp7kApX5+h4XYFd4
nXCOJUKmmr/6hkOisajTOkCwc4nvfx/wye9IYyaIypU0Rq4P6WhKwRkN//hKk8wGUI2c8tkoEML/
7uY5V5NNeMwx2WR47pIcN/+VNkFYKwkj1lV6sL4eGMcTWToCk/x5Y6gcRYqv9OgwW3D3QEYbO+Sc
Hm9DFore0RSqayJiujQY9MfMZZ0/PEgb2TF1mFxk1vo3UGxPcUvrUpQ43tD8eIoQn5jwEHq5rQy7
9ai71NTJ4MIDEI/22KUduTS2QjnG7QMhwaFqNh2s7Fwyigz8BhSVP8cL6r9N/3GQvRNhlbIMwkve
KgljojkD67F+6rWr4iFFvuoX97KHvpeIEo3DYAcubNfGGHDTjZlmcT/fR8sJgEVj7IhHfGlq2wkk
jW6586v3HrrorPxYl30i3iYrovw/XYKgBz8EVE0gbkZTyb9jbPW94wz5bVumeY5x/QawdrP4biiO
y8M1gXMKOCcXvz/6CdkDN16UMIZxP/oxvRm+Q6xxUYY66iyOZQjFlCt2Y270pYzYW5oYPyAOh7Yp
RxqZIEoKbOdPdPYFf5kaHD0cZnmc10ldwldQswpeV20WPxsrQfZy+235a+Ki9vcJmPfUCUUrgmMK
qxS1f4nJjfAVPijNrVDlfvYJOxjiV2ciZQS8NdW0gdYN6YYUV3nHESTuIGETcRQjvSabnMNzNPN2
SaZjojgnr89Sv51ex6RhJ3fgNlmZNMiAEaBRG+RM3p783pYGgduaJ+t2H6aw4N/+8mK/1CjcH8Gj
74pH4bRsj5el6gMsnlZTsJYu+YTNHPe+JF0qjKeTu5/P9ohgB4Tyz4/vBYhdMbNkS69Nr7AestRU
ijc7PxshZZdnnt4E155OyJruoeFWDuSqXlwGdTHw43YMhLYFQ3D9QLoXljjp5coktOmYhmfA23Pb
yEA0P4AR19ynFgV5k89EEgzO00wjdfIpIlvkSFFxgFVHMS8tNZZp6wf1Zdv4uXy8FVuHS9tf6aqX
eA1VjrHYXyUGGmUm7Pz5XZhQbDZXj3gMII4eGUIITcLlBE9hxe2ZhMOu65okKS191ElQYrwCC9gA
j/wmN/P5rX+xnctX9l+w8OnJFAPViYqLBPNQ2u5qbTQkUyL9XA8stQpz9sfOj9DZIhYyPBX9UMRX
h3yUZVfA2zNeMmNdeV7jzCCLi4VW+Zj4+Ttn5y0F/iTRuz6hU3zYjWDU5/0feptvjzOr84/LbP64
C3Am9T8bLfmFn9OQkV98RWpaYz5L/89MBz5qup94ozzP9GOf7AhWFb0Y/fKNNAh+puUb8EDtZG2F
hs+37aTSSVwLuMIwSKDWsNTJCGn77+/F3VVO0uCxUKUeXKT3ROaoCdzXIUyW4zG/M1gX6Fyr32s+
fwHFmCOxoEkhA2PLsG98SROCI9Zy1UZukpdGughnau9/dTxIeKogpxk4YgFp0kvdfZygiTYSdeks
cEjyB5OLyM0x8hFjXNxDUv8HHZsDtM/F99x4Q6CxlNa+Y6JqGKCA99mfL45Z8e/gVwixSM4wsuGX
MMJhBNnAPA3O29moKahWuyV0pZciDOemKQUdFKjTbUMGnv0okIm2tlVucQEVcTJAK+LnikowH0wA
2HpDcBMKaxuJjKUPtIEXh/YiKw9gWyzeZAx7yamXWw7BS/Zub7BbDw6dr9cYUFHzVkLig/wyGvvB
CD5nf2zvMwt6PY3Oy9R7z1yNmOgNaKF+KGQfRAOwRE/W39Ur6/rIZDpXbQz2IlIlQUTjTBG5KXWc
tLGBg+/4gneFK9SQfPFj/QKklm/3m+ViINYHFZJiBnJMuzj+pdGGiApJUNlMNMAogKvg7CrrMUnt
0YGJ9OahlXQdZBavRuNsur7flgQO57wg+JD/7+QYqhercZ8TSBFB4AoacCvoK6DPwlKRud9CY9Ue
JdQD6CEuNVyWh53LFZjpB6U2m2XbUJV+FZAH1cs45nNwN1xBXssJgo64tCJ4giHMBQve+zO4Shll
UKbz2uOZC7ufWzemfGGvBCBK3VbUteHau9RazCHw8RysI3k5F5t7zTKaUNraXI5LNoJjKAoMIQr2
D0yfwk9Nf6HaeWeIS/v1bgMp8qhBp/+08h+NFGieNR9Pnoo4s2E+KP/XmQofllzrLSlqzaTV+Jae
5ZfkbZlH3KC99SWakN23TEHcXgS0U+Wjt8wKJZ4fEczhb53M8hTn1FWLrXfJyhxEb/aDHWsSYXgG
/Pm4f993hrOud0mk0v2ZAdGMGF0BSTbydh7O6iVnnOZt5R7dMJDufRwdSb5cu66PAKo43ODMv/c6
gcHXuG0M1IlgdNBnuzI+Q1VIYThl/tORaJWFYBZfutLJoXk8VGuY2/YutBbJR4Xo3vcTelr14MjU
EWYX1ElJCodESUdZmHyVpYpd1+K3aib0m6ewCjOdX4UanBH1tZojk5xCNmzrd3xwTE/EUL/fPK0V
pM63RTQHgx3u7vwZj87tVnin8eKWoIMak4in3h6tNso/i0Jen1fH1Kd82jojSevh2kGDd604Ze9c
FsoOV1Dwv6fcLEWSxXSd7ICJCJAwlS0QV33czuyLagqKCr513XPkTEohMHb+95laj2xPg9FI4r/I
1iP40bEfOXXKhIDEAwJ567taJLJlTsNtgMD1h5Wdo64Iicbseo/LFo7KbWtitStYrsZHaQ8w8OPt
X/iGPLylyNvm0VT/7cx4bImkQ3nm4KuVkOQIUG5z0CmuyumibUFlSmGpjPpAlJF7KoZtbqt7KAnl
DPiKrQ0sOkfo3ym1o+yQLwOvRlgKxMirBknreh5XFx30h5jcTTuXofVOREN7fIUmrwTs0rahVwnd
wpgoaomgy0wgE3ss0IdBK7hxc4DWp35doy57fd9Dxr+TdGxN04gwABCNccK+dDsXnfcZ3+1Q5cax
2iyLmRIBgXuBCRxmIfN2QOS3oIhJAnvNCpSX9DD0UMjI3p/7SF9urpZtogmMozkj2F448gZETHxz
Azb1lkNK8ic7ijAkfj3Kaxha0mwc0hg6I2yp20dI1s3oC/NE3kq52yjJeOsiYN4BCeKtm0SzJUJr
y/goIkGovK/3N789uXSDM/cuE/9j1YfAInogjcnK0Onwin3VxHOW4/nz6Fgl1WYwP8SFTduooYO4
hjV6WH542c2zhlgbghx93fjInpDBrSTPyh++nTl9yfB/JZ9QMzlRrT1rHM47BfTUACZ0boM7m0H3
0BCCu+yEVJChy86UuYNeKbL9+VTfXpjGdxZDk1Ze1mulMWJX+gbGprp4Lj8/SYtYRHphxicPRvLL
uj5bi7DfVw3jUvGdYNIbrbu68IcIgWvjWd9apwVFy88nDnuCCzWMbEFmLYceYE8i2OAaAITASPZD
c7sRNMYShw9+UU4pbRBAxudbMBSUU9CxGqamYLd0w2ZCDrrOATCypf/DbPIem/N5gwCr+5P0d8ss
9Ocvm95BWA8W0X0RJVx9dLVjjkKW4g1dUfN/48HdGIa73V6vhJvY2CpeMPw6bgt6NtL16FaVTROC
4+AF/DPz7O8queDjz9p9b4Xz1xjo0XVbaVtczxRmPB7kUg6UHXnTGX2W49dHfyRH+BXqz/aDQGFv
HD2KVb3KpBaWBApubGRNiV0gKvio19Ac5cGltZrEZZ1ZvQ0j3ojvsXaWz5P83QEa/dRzQTISfUia
ALsu+G26ZU/lDXzeAO5PiogLfL+wc2udOJErr83mZuMM80xromGHlIO/r57yUK0n04jgyxHoGCOL
j9vnxZ4tU5xCpnvwuDPa49cmr0Qb0s2nyivqgerfjNL8Mnb4S3ZjsGN13NDolgRu9OfBZMOuMCTe
JmiuUwSti7ScP9Kmc56dI5hZgMuLpnlVEvT/tjKxoAlOah00PtwuahsDwLWlodPnX4QlXz21M8X5
54ND9IgokUucYCqb32SSuuVMFun6kiuWqA2cTNE+dUINOo9g5cIBlpELf9xCtT9yB95x0uETT4mZ
aISiDa57nBmO6WASixoFSzf9UnTfcMSW4ruj/EbkjdmQ9u1LusOAgFkR6YOS6M2MT5rtRBStrhqR
qkrW67NiKPOjBdt5Qp6vXp/VkzX4C8kvklxdVEZg1JvZRF2A5jY1lBQ8Bp59sgClsgiWeEhnvOPn
Fh2VUnT/kfsTuU4FioQLSaW/Ezs/1C9feLUYTxaVv+DvTSI2nXjg4WH+HKHxQImWNmXbtr4QJszy
lZ/OIOtkV4GZGwkfgFbK8E9OPIzfigdhddCnLb4KHovfubrZIFavDAxMNHIYGkx4r03aSaqHm7/q
P3IlAbdSpMie1TQ5rK7rqTzBDZaDaRAw0DSB2FBkz2JCMVFz8yrbA9O5VriXA/ykeuk9P0KhKAna
2+bUm67RIV23ijkJXlpz3/JpCnF9qM2sHWu826Q4zaQ/xtWsBcLqTmRTqCOh6p9y13FfTxU00vxd
Frx8EB/1PILCyG2iISrHcx/TEQSZs8W+5YD4DJ8ne4KkUpdjGXaMQhr8rvsuh3LsmPjkWow9pW3k
TCdhTeN3MnXU7TkmpJrk3XArpI/pUeszy2t8D4c1KE70WBjivsuxvwEPAK9N57mgS4LIWXbyIGjQ
RNWJM2MklccMnGuEFA2ROs9loVf6B4I7miIgVxYOFHPLtu1lh8Yq/PicdLW3EzPi78hJptVTtT/4
J4u6XLuL6whVLSM4kvawHcZu0qOdTAiIJZj30Zk7N0QmulIiYIpHAhHjeTHVaAPR/My5wMp6JRAI
gchS9lL9Rf8vCVbf37I3Vs4LdNtbjVIytfMyWm0RUvNrZWDa5tkEsGkXXJfMmUauqijuRFH0rhOJ
EgxHUU1iPHZJG1Uba55weQXi6D1Vto9++CtunfFzV89bJGGe+vGBWpZc9KdtZ0pWyjkAJTvxkffo
q195arHzSQ4K/DsZPPmixNJG7kGSJYN9c2Gf4JoRN8CNriUwSWThqXvnV/JZLf0RiCZjZOdg/xUa
0vw5GE77dk8M8Jstc5kWD3K2ILzMKuIPe0N22SiLN+5PV/pEUHWpCx/jbbvX2FZKtVt0/mPJ8m2A
zblvF5h+bEipQq95KMytfIWQUJAnNNjfTucsRlw7K3IQA2N6xzUZ1SdlUZ8cmCOzXqM1EHHtWuW5
0603zhgYyMIy0ww3/LeQrMVkI0mqVBW7b2RZi5WJkAWmBneQP8pdR9/ug3qVam7QUqHwp+Yy2UNI
gkzAtcWMJ5lkMu0FvuINPoqqi47RIhvHk76QB4osb45j86C8IbQjF6g9JJAxqqLpDP72VIqhL5gd
hK3xFWys5flfq+tp196/jnzlbe6DpA1QiFriwcL4d5AE6EQ/KF4wCzH1zKGhmFC5VDPq5CdsYqfT
PXTBmDvKrl8i1GU3xB0M4kz2z4CN+4HLKTMvzG6k3KZf2poJxmX/NpHYOftlCv/As6X7b2p+PoyV
EH1jvXjw+m7HBQ7LUnUtEkYHAhSjF11L6I2uFIK+lswERXoWwo4kXVup20p8IMJePuBf43Om3EkG
mUSy4Tt9eSDHxu0Zm+E00Ap1iGghDIGnkzRwhiNgQ5wq3lruzFLcUIydhc4kQ0QSRWrskbznUdMP
+zV9qWxtyNzVJQFBvG2aqwRUysUByd9e/fwaPmS1X0NjDkBTMll1JsA3VzOZuJdSJ2v3wWDcg5Ol
hFvcemVM7AXuIyVDJ89caqUW4XY/c3opPt7WDLZ7YUCkuWybUaBCfUmd5nog+/Cyp/NqIHkqS0aj
BDWIS4Cv5jk4tiKDWUY/NLVxzK289d70U7mgkXWEyDganJGtJs7yu5ttPAOtVX0kv3505hTwLwJe
E0y9KYnIiIwHEgPbrWfx8Mxg+tYQXBZ6bnu4480t79qzghJeuhIT1Nr38YZ4zeO3oeKmsr9a24YS
Cn50SwPNjd49bH3I2nHYMiQKwZsIoWrPbQ56pBnDgo2jR6+qJrqn3hh8y1CKd7E3M4I9ZIPOhzsj
jga+VuCkA0f1XPTuorl4Sasv1nNfWjbDhyJMW7Xqu36uJ0vOXN0bOgFttOItvU/nYOfJJacwrOgF
35iub2rHUBpQU+6nX28r012QaytcP5sF3e/fV+A/vA1Uzfx8Q0KnMJzEq/8ZJq4vm6rZBBJ8+TUN
dE0kohH1rIugs3P7zSxUz4jtN9FInelaLHoiuKPHqTBb7jX+3aPx+uFmIvvQRE8aKqKNnbs4D64O
9TnmQbjNh3uwV1v8FsiFpigJKtmyyfSsscxh6qXv4y1HxK2p3bWWj7CC4ieR1u/5r/i28O71tX5Y
SxTM7ZT1ZfhLfFB2YJoqT1Rd6VQ4LLMyPkSEcBofy0ynTSw00fLeQJ+3793/bl1FBTUYFQJrMpQw
Mo9zC5u435327YN5Q0ZfrR11NhFLN0BeFQJPTz1NjVV5UGMO8k2AGo4KZQao/dcKoHUyJTZ2E6t0
gO1LyRB6RS4ond1Jnq5VEhaR0rIlmUBlneH7526OT5I274a/FLZ3wn6AEU8A7m5Hi0gFH0WPX2ei
tQa7AX+jQjT/j21hZK+ZDIX/iKV7alavO6Fonhk1/ECnCbPMumgP5AylAbu1Hju4H66NF3X0mZrn
9lx0GeclBAv9FmoMLXtyOKiUsVmtPPQpZyu6A/gMMYEi0hQ/bdtnz4mk4wMe7PPdiGDjuXL8Lrxw
EvY7fWTf2XUOzh+dHrBQUGAzWKtBt3YODSTWqbEY0Ueo+iIcmsW3Hcgyy+29pkHmwGrLMuTuR/YV
9FEMmbBmdAFuGNnnhcu4kj0/S2JYxbODsTgV0D0tRnpsJyqh8ZQQNBVXo5sI59dwiNmwhpyI8/EJ
Wxdv9JvD+oFiR72rwgrwLaViHIQY92kDmQrEJKVIbR+AgzYY2XT6n3CEt/g0/FlqyHk1yGffkv86
HIw4uApyRHZU7GoJkeBohMHD8xRzsYWx6wa4k/BAfP6Gnr8IIUy0LMH/VOgZGzf+rzyYnjB85AU4
C097CrUsMPvCv+HXL6WXaS4XsZ2LgAeuZM3pK5ElrU7pk3h6/uqyKIX7/6o//93UNIQz7nUzC087
rTrQfJfduSYGFKt8hAIx/4ILz4Ek3q3eN2PG1+WgkpxZMK78fuY6DLzSXfwPfbaz86he8w+rlgzt
L89nFOzvh1dE1ADf3Bw6UdhsvEZBrg/5KsNoTumqjNY7VGYwODcnJMid9cZ296XkeQXwG++FTdHN
JlUO7mLSrWwP4DqAIXDJlDu4Hz4zA9dKXPePzFCNB3paavX623xdfDVCp5VDfExZS6O5yl1KNZ/4
nzSMckdeQdYQ9qrRyE+k8M2dWRc3Y2wbBKzya8t0swJJtjyOzr+Uq4gx5axQ29oKraICnLNOOqib
zD5QAAa4ECdLaAMB0egznfLbQ3935U+2bNqyxf1pLYzmUuH3YJ/Zdoz56ZjJd+yW2y4nfQ2xAmLe
B3DSMDCCj8gsz12KMbhZX3vy64yOyO7hUp37kup/a737nOFSzbYiSXSxrOLq1XbNDl6eFbI5fxgm
0mBNxxagCH94d8KilXZ2Pq1qC7AAK08V4ogdmnb0FvW/Iw2DyNJlnKSNUFhXnyfQuOqRNRyD2Wee
A8pe2IurfggZOMpVnJLp3sEMmE8XrVd6gpzsOoQClXBDmaNd8raJIJ/AoR17wS3p/OqkZ8U06kUi
dRT/xMyf1z9yer0vJ1riShTYtWBYVoSxPkwofBqvwIByyk5e3/QIbDeBrSqmnN5P1oyAu27ue9Ch
m79PcFFQyrDvzYDlWJCtAtSKDBpBJi8o0Wfp7EDWSYfEXy050xhKEbiGLusu1MI5/89p/z3HteLc
IpRxdcclJsPykXrSpTCUCHQE/UtK49koE8K/0h6WJd4o55iX1rLmJPsMR/qpzD8wdLNnoFrjNbYu
CHztIAin0qHsrMEhgZM4VfbBPKLH9S8n09X+1l7PHqlI/wtbBGKqZ8JqdTas3tjZSb3RGYZoAgbY
tIU+WSKFBgEeYFRVYlDvpMtcH6ETEURmjvQsU9z6px8izvgxZRY7zS8kNbLsCSC9VIVoXhtY5svM
8ZtUZDeXPAP2/MwyjE8mA84wgr4xnmUDLtxU+QJ22emNIia26CA7mjixZ2eLcXVsJqjEPCMg9TeS
328lnhpTN8RMUGjF3Hv+z0Vp6jeT2g61mXzRBIq0okH64zZDGl9uJorxEHnI9/uBFCpIVkNqNE25
DZm5c5YmeFDCXll+pL5LT2HNFWXXfrMv8R5GRJETHyfCguHCDQ/pdiKINb1WFSAChRbWDlhFBBfU
LQH2IpQ4hFQ44bg2cp69aEqq+FNSDwwlwERXG45/cnlkeKCFcdUQf1yRkUOD3oFeWpyW0BAMUlsm
VOvqyPa6b1Wz09qrR0Gnt1G8QpEtgjDQYPUaDsjtS/6zT0MLZm1VHBzZLUMpg8jA1wb834t9UyF5
Q+FDL3fVB7xDcqMM6qx6W4Su9Zomnlq4mBSa/vJ6aXzpgucEn1Wl3why/RoC6vcOJqGHXM5777G2
dn6xNvuah3C3Gys7MCScQJVKtxJEQQJ+J82WQCo75NdPLgP7Ak7wonU0xguFrcePaH70x3e3tDgs
Uo7dZnVWr2AmgA++Dx3Bs7ILRaze/Xg/jz/vL8osp7GfjcQHHrLlzR/uOOC1yYgfF9i7Bs516lH1
yJmqO7Mv5NbCLfsLmUzfEsp2f9TF5VSgOsieBm4k898FRNGe8rO1qAmtf7ZYj9WmjO8zlFQwSvzM
ONSko2EwCLsHi41xNXbQkp+shW1/gKIS8v6MsPpPBRgeRmePISKcyotiSvIocAhOirCzqooY9ErJ
fDZRTb03BYFEoYRCEFqDoInzpaVVR+phOynwm7Haa+Uriov965ijepJGLtJDQM0CC3f6qxKpPE6z
kjl/csSJr/pU/vwHC4jeKIRngFRB1l3Y1eqa5ixNdf9GVz0geZ7pyvWI47lOMX52Fdw+5bVOjY+t
fb7FXjX4uQvWD9AbsAyZEKMwU8rIEY78Q09XpbDigSQKGgT775dsR4jGpZ2kXg8EFyluHTv3PVXF
cDTUgBornOjlxddSup2hKaglrGJFVKne7psdgOL8oEL3x8d96iJPd7dUvLESZwBNAQGqeh4zMYso
QhnfN8nkQu4iJS4mrBnj3/fgzknQLJ7OSdRxoF2S7rUWyR3is0FeTekDM3GB9OHX0jy2/iGsA4UM
/x+YZtrtMMDFxOcvyYnOTtQfvw7l1iqXKHZvF8nZ/Odk1jLKxM5Nxv4Ph8TX6ILlDMToIOvJQwmo
VWzBnvZtyNvkOENU8so6gix7RC1Nbp9+DAJjLTc0zMokI4zBYYbi9OLhTHDBT3UooBxNkxy0KPdZ
SXm1YeaG+I9XlEoxANBplmuI5MdpOn8nkzSseeY3Xt76FDrgXHRgHZHtbmdCw0kVngznYMFsNX4D
zt6XRG8u0V0wzPIwNJeYccAhv200EF3sES8whreDsyOdHmpxIa0ffpeL06z+qRd06QP+w7jLLJRN
Y1w6Rnl37u18yXQ5kVOJ/lu+f3IbeoeeEPjN3u/a0YRBU3YZ/mpvv3Oa4gbtVYjghcL0+XnoNAUy
86qMWjU9l/MdSEOXTYGMW4KbfJNNVhTuUwWEY0tAVfDIfdHKGjUlLg6UIOAXaehX8spk86VdSH8C
46DxViM+sD8ACcoevTibwv5dhHi0lvd2Kc4FiyI8VYRXi31dvpuvq/+eu+KjR0brm6Vwom314Ytl
U0TtZnKMicUZI7kVI4yW2BXEBSbqvtsVNJeyYGRj7TZkvN5RaI7jVPE/olWT4jLVI4Phptp+K9wc
Gnmz7Tm7m7cCDzgVYGGGeMuqQHTgtkU4SFshbwn9Ejy9CvqvaaLf0/FVp7nBkZ3zgoQ/tiobYif1
eYCIbcxZoukX9XHSEIN9cf/DjqBHZZEu0V9z1TMv6QuobDbOylS9RCvHOtPF6jO0xfWiLt/zc6bZ
2L2OGKvgJd7P4RUfL9hfcrW1ZwnGe0n3yOeRzMSbeColgxvNPj9Yh27X9wmB2DGeRxOGj+PBy6bR
wBDvRIAj39AP2Coz1v3lCF6aAFYtuZpAB4YzjyJ6Ya8oUliv18A3XerloUy42HnAxAcdDrFHew7R
t4dbzFqmvcuft8aHRXNJFCWvWi23Ev0sf2Ae9UP3cPtnaJeyP4GfEksdUjWSLmg964tb9QaCZjp6
ZmJT5rG5lTnclXr22p2c+ugImFC19Y8NXFKWWhvvYYg7hgPXuDQdlsxCjFtLx9Ohefu1QvYur0Df
rl62O8UWZBz6+IAhGikv6d10hdNNVZfQI4GMZe7FqU8Ik5XiGNOTfXZt2FOPP8fMztvN1V8a63cm
qJfYLY3/p6uhcZMyT1qmjiyPR0n6+QGGLgdWRndxt49u10Sp9ECxzTIKbms28/CC+8esd5EkSFYQ
bMcVHAAcXZvj87gxG12bxJ6pFlsThoiaR3IjSEdiYZJI7BRIKf3/GQupqyjmdb2nSDvKJss/Ka9l
yy5+rZgvlaM0cjkYmPZSgjbzmQQNXiL6Yn5gS16OZJIii5XEoKfY5q6LpHRdnKRJ5ecIMeQJmQSJ
uLxqhXKUss+mdTetntVr/MmkLx3WzZQviiKOqdnXp6ZffoIbkcQhecEHOTkKpNuf7kvNLQk+7JCE
AKuYkdgiattFcbZR5UaXCDodDsIuk8osgFyfxoOH7TK+PiCZDdVOkC1FlLmgNGbmS/e0pL0Cu5wv
NHjN7N26Hdfcf6ZmudmoNN0qVv8fi8w9S6cqFBhKCc348sDBWuAhZO1+u1qsJDLszcYNATvDbcZ1
XBQWmitUXxR3oqQ7FQ0uMLkLJr9FAEN7MBXqP2+f1zVEx/mdkY9ERtx/uJ8lWsnE/UBJDH1T5u7I
hSYZiqH4n3I5p9I784WbWPlvzPhDN6pcUcee0fSR+Anfp+gD9kF6j9lx3e+QRI36zDi8Ca/OVAxU
QxRCGO+iN2VdjJGRbT3q/kHKt4QaHez777titvd0804owqo6PXcw+hiFoGhogK/SiKXPvY4UyCux
O8RFQv1TPG1xPTcCuV36XkrejVeswWcbxeKktWX2TxZizEdBeEMMe6ORO1voihsg38U8DzDR1U10
XH1lMn1aT8QZlimXJaDbl+lOH46V+jHGjeQLjYaZiAGMaXKOxv/fhW9YelnB8TN/tGzR/9Tyv8jU
WXeBtQHtZ9754bdhTVbvfQ3drj4Rc9NhJIqEJmjosD3ZDu9Jdth9eHFTNTkNADJBfSXKm+lviXzL
N5pIhT8j9FRRJ/ql0EbGSLtqCZi/mSBk00Zst/VmPzwrKr2KFOY2c3cS7B9fOgvHvZ7qFDPHmxXm
t+MPwVr/V/jSERPj8VhJn+v3u+KP9iHuqH9XbEDKZsDWMstZUbVQWYpXmqbkof+Hi5iowTDQGkQ3
jQjq+qRJLk9VRPQd7/JXyrZjBPHX3yopi5ayT4hK2wqtYAFHXd3tENA8IQPQOA7SPIKb7k+qGKkB
Jqr7SBHh1bpQVseeF4KAYXI6jtXFgK7ZX4um8V7asLZoSfTB7K6XDff3d2wpXFzqfd5hemQ89UdE
TKLukPSyVKk8JsovTLcJ787RWmOsynzlmbmSyeFzdfFYOCuvHrApsRg9W2yZIDBjKg90RKsRqSSm
tjMWeo1bQsaiMR7zAf0B3cMjnYK0s4rXIjHGOkumY+5VTeovZs9OY74Ws9IrJl4BMmoC5i651ab3
zEfmql8ykHIaai+neZZNVhngwDm7HVETWIMO0p5NEA6mGf8cmJtaMHmHL0jcZYxPll4PbDxEprHI
s8crMX6uYEXYK62nd2DKIoR0R6i4RbzKol330tHPIYnq1dUhvxZeZCVS2wWJbAz7IgTqPgm5Y8xR
xQt01uPjiPvFvzskcrE+pl7fQeTDsC7MjJfCioAB2Q2jcS/hokfRemIBVEzzQWxWyqel8df8bKM/
/u1snZDz589YE6dG9F9jWzTXh1RwPAFN3LOD4+eSnUO2htb7uX9u3DVNqTJVFjDny2qVhYHXtCC/
GIrtIkUIKYNRem4i0+COMHh2OG9VH1xaxn2htpZHjg2nAYh4Wmxs9lPLBV5xXIatVlUtT4rLKziV
D/tmOJUBVUTRf+LKfJyL6YofCxUNpRxtau/p/eHvojuCERQP+36kHOotM3jB+YwCK4PzhLODL6d7
gloqI091W038uxcMr01QjOavVIkuSWHxxK1O7kiXC9AZ1xVqj0mKKbqebwrJVqDvmg5PErk6pwiQ
u/+bV0WYszEhLH8aThmgLd61OZAStFDQEm1qzSCUT+fXvWmARCeVg4nInRcOXCR1OLd/xcs+LjVA
sOnjQld5864w2FJnZzxJlSzKvYqKYUiYY/GzSywWD+XJdNaspVDxapplU0RtjLu7GSC9lbPyn6Gz
SMeQNQj0WUcFXm7mN+Lcjn4u2yd1wvJqBSIBlUI2zkCX5qFQyZqfDehNcwVZWvsFcf+ZRtXyXOT7
w+SVMk6rEVwTzNWqM1ZGkKfxI+x5MWLVSJKVOJYyRkcb0pS8hUIgO8VQ2NV9QgI9O3P0JJOK9g4g
GrYYvIFUCMbAHZls0wYOSto5NbOzIidbavnPKdT45Oob4JMWa3bh+LScEnVHQfFs2K8kU9icxAAY
IVi0sooNXVLobp6roie8p9OE5RAICnk2YxGiWHlEK+UUr3YIkWYrGaH215EFT2/8ZYVjUzuXkybe
Ic2pnr1LM01mGRZUq4f49iZr+2+74Iqjvinr3FBaOLWEcab/5ThUC6FTOj0UDTukon7Pmb0KsSGW
q/ufU3gcu6VpSaOQqPv8+3ODEc9gRIp+vc6b8nlb6U6XAr8DD4po0roaaK1xFEKBmUlFEwqY2687
NAshcca46db8ZhFwvv9v6LgJABo0Vmg44aXq3PPaXmB1DKgxWChQoXiXrO3z40Y8uV2BWyn7/Ngl
c3gQf+enNxGIMN6iqlgl0AKKri0dqT4lOrgTbkeMV3HHGrp3YjlP65A4fjf8I4ZQTGMhSZQOSOgH
U5vS4Gdp5Bf4UFO73/xHAoOZNCBOaZYpziT1EISLvwsWUbKouCUJSCtY2jJhQ7t3MUETFhr6QqL7
kko49r7nIb7saAP88CuvoDcINImG9IlzeCiVZj2HUscwFx32fnzicz3Ln+XXuz83xuoToCm1QQy4
5vXjPJdiDsQn0EoJsb3xtjT9pAcqJKX3w9D4SpwiE+kFDKTwJHv0dJ7wMsV3AVHCJIh+dh0AMFcP
CiYjhAKJRvsQMyqHTUu9GvaoR8UB2loNdbW99Qv/JUJFJYgA0z1AfWD+kdatehlUgDnkr2AiBf5w
zX9BXdC8T/tecWlPXO5uo/RolsSbeu59mz/z8fkJNe0cXFebLaiiUosVyDYnzK+qpQIbY5T8mh1p
VHdouRE4UHesohp8nEXadh1LfGBYvGZuU4P1ia9QTkK7ASyrz6WX8wABAztnEJUd33vBOL7s1od8
N9hSa0vx0jgnefc0jMdSW6C8OggL0C1y/f94YqbtpPpHmiKilzzVsaa8Yb5zQnxxBqqdNufg2ZAH
q1CJ0NdD3wDiNxfKhRMtDKvf4POwb+99TiGuWXTkoYL81ZeFB8OKiXhwDaMzQedPRa5+Y+T+g2g/
HQIv4JjLYX5kPm/5ODDAoKkWEwT0tUxuuSol+XtlDj4+8P5L/VE6cjUrT1ccseOcHnAGtUMN/aHW
L8hjhISmXqauMkAtUR2hY1AFcnsJNoenoJod7DBIVmkO2iOXPWdUutZGPmHLtSSYelgQKBzLnTg1
ntQkSQzwQN2p6iRDwER7VLUmSJaiBstGl/jz+UUMFqGl0TF6IREqJaRvT1KpPNRsUgKlm1GDZ4bz
l2YwsJazU9mxKe6GgpPORnVBa6pURuknhgyOKyMLi2qwxqbMLd22FFo5slkzRdfLcUWzCB0dhhtN
FNAr2XgMn6aU4zJojbIyNhNNeO2OGqwVHnESVewxD+SZR23czCXdM+kGhqCYGBoGSKTyJP77t+Ye
XDuf2JVdbbvNAAUupqDolJ9//RIsD4vF8LSMl9g/DtdiC4BIbsNU1HZt5LSD+wj9e/sxP2ziqGOy
gChgDJbeSgSlcseAUCL7Z/MRhFlsZVjP5YiSg+vineRl3Xg2BqzwckVgAlmaIQFETU8iCePvk35x
vvtpTCItSp6jKCUhhWFYeHijDWFgzOfDH7/RngIZEHFk+w6qXf6EYOXGcMuc7qkMiKBftJy4poqv
WTwDYHUQjb4Son672VkhcaIHcTPZYo64gm2fWJiTZvErinvFEgFFgfy+Zctjz7C+kEi0bre4phhd
2sj62o/iDo/Z3Nniekhe3T7WH5M1v95f2VmGXYOidhvUXleiTkVnr+NLZlR25ZQjjg+URTv3b/bM
T4SVdCy0LrHCtWU0Cp0IDtPe3X0aOcQUJdx1hOMysVzmOOqsb8lPTsp1spWvG/tO2/i3i2jCmU1x
cZrp9B5W25On51E0DwGXCxgO9P8xeFO1SgmtcyOrh/fcY+iPheRB+PljvBOMafHR1dVaKnkYj5Jq
CovdW3vdZtUaarSAuB/UFGg9jnSqVWV9enEhe3kId4FEP4Rf+N4AveAq4SIATJ+qy4+4JLocg+MT
DyW2ux81Y+LlJoq8GUFyT0gQT9SqMwm2JlfeuTsPSGPy2J5jRLqH4PO9acWkJ2dm/tCP8MgNTWBR
sEkfI4qbjKR8B5pMCH7zsb80WhULxzMQhXyqqMAiF2fzFRf5/bg9AbOUhyRhCRZ1ns1IEWAQJhOf
u625bLTPrSvQKPpajwurRvXu8O8t+SHkiG84CjUcC3R7L+qOZbrAkmiicqVwDJIO5my1BG1QSRY8
VxbdK+RsMuGFmX3vr5MNWa+I8gWUjtRBh8COvAbSwHUnt0TrFfYVnrBlBEmjXjQoG76W9AvlAtE4
kZJ2TR9gU9QQ4t4+Zu81ya/4rLpyk526a0YFCSiUnVnns3sRFOeYb5tIt2f/ASFRD83s16oRRwZ0
/P1o/+wRMHj0TnmEL10IQ2VknH953OoUVwCefc/79ejtzkbbQ7unNYaAWfHAgCLU8TsN6RGjiw5e
ZMf/UA9Rwz2U55KM0BDUSQVRYfoUMNKlDdCfrQQN9+r53u2eHZsHhlZiAV3YxL4L4SkftACJS62M
+ki507+KJO6HcATrFQN5iJ7JzbDdtBawpMDa5oXU23Ht3JnnfuB65yvo+b0shqZKbtL2QXHiZIZz
sUXJu48IA0xchGovtjLAqTKAPLmqM1uN8kLlG1C3UK/Cp792J24uqI5cXtTWkYWk/mwqNI++RXrg
7SGumjoqrY4Ro+pKV4KKA8T4pvvic+NA3+GSk3YS8nerdgjZWDjgQbobo6fgZB29b4EBWaDtKoDi
uyEEzzBnz6kRDU8J4gWDqiMDNn5l4A9aKMUOsgeh8p596TFw2c0KK8eN1C12AGgclZGr96Z5ONG9
vANX2zfDErkAMyqYnu7gKWrdpwZc4e2SyCUSw2ISlJLdfcdXsHoxCLAvwu7xotxsre43SszWL1N/
Q/tDJrnTnz35VVnPYZciz8gYIrXmvROKueEDL0SvBTDDqe5GwP77lrIHtibmM5XTjLnIEdGe6lKs
/97pxhywR0S81HLfMKaIYyEhv81YcaauKz31gyW2eP55WqHB1ntv9B0+fGrCFPYASsn6MwmtqCFP
o+umLpI6GNo99lxj+jKnzwRLuTDp7HazxHBJKe4tnkNWz3vQ2pkrYJJqOcF2HticptHqR5/ABgu0
i6FKo6AmuIm67UPnMo3UNXGGfKKuVtU91COmU7z7E58CnXZYc9VYdTyEpM9CJbU19qu+JilgRBmh
PEidBf0y6SpUUrcdmDTu5i8kYoINLa+SpqbQFenZSha6vHbLnm8HaRLqDVrgvy4wcuVgb0rQk2by
peepqUahU1HFp1KS3ABlaMUxNDgM992C3iLHyVaIpxlI3jUkSJ8rVxpDD1/Kue8+WRIv94zOtdco
dpjZiWfmWHozLsKNRTEFJyzj9smwFjBgrSTOh3jgzI7xhbZXpq9PhNdP0LrfFBAawZX9219M2Jma
pb1pcXbXeOgUeM8iPg3VxiupMb96TwF617zC2Kdk18Wc0vRgQRz4guNVtjz+T/rdMVMF1Ml53Eei
WYghHu4fApm7WgKCM5zFEs7WRbt/iI4lpUTY5DlBXrxEmrzmbyVMN5X0pWlp/9FwhuolSzvHSkYs
t+tljjrb8GuPREjIx9wjfHsErKFXByUI9wtSrDlCZ8wvld6xYiIVloByAmdTODdefDg5Udh4d1nv
5To+vPKv2RA/oYcTrlGOw4L2ZEWz9NaFLHYGpt9SSKNEYqqL+e4vqiU/CkUjmpDZkuia+eKDTRZE
H296PI+VRA4Pu3eb+ba6HGFdLYIg42VlcrjGuWkFEQ8Pyk8y3NKBe6RlZCrArP0EOlGeurLlqStE
GKQEhNukc6BiTNBP0hBvtVCS4pLx+QoQKgdn0jMCenQBT/63mHPloe5cNCMyJatQeKXS8surOuAI
4F26iljVYZuDO0pSQSK3DOT7acmQIvwYhSHoOGZz8nrrkrOdCn9GrtnnVCNEKxr/AeagFy6AbNND
c+hHWYAYSe6RzeAQt7zRIncs6DCzcMSTia6uslprZV7y06KvLUOBi2iiCR0Hbc3HD7/0oDz3n7be
6a4kV/7YUkCTnqeLY7R9lQaUnEhj/ggb5YXUjIVD9lpzGXz0wo4n9MEzI3zJpBbe8HFfkZiRhQYv
LIsi8UtfuwkfkfvHC7C+x3LT8S6WsEvttw4b1OzTN8BZQNS001dkI/2p9azjKHrTFczr6Jz/3K1h
lfkb5eA6RWgs2LBlmkfI9nxrDQqrk11wBr10/ghM9fr92b67RaOPmZwhLRk4c4JWH/EdfYKWoVGT
+6aI4eyxOmx9rsLKtgnLOT7J47XFGEcCelS1IqEb/LaJgcxtEQy25cfVpNmQ+KOXTwgJAEhJAMXb
bAq0B+fiAxPVNUzl0B4j8J+eRwFecdQyPdHA8Z5Lw46hSBIycdtPTlR8eYpb6uSMlyzK5wUtQmcH
xZSGLcRKepGSswMMPclpQ8xk6BNx1r7iJ/YkZDF7EB2vCYwqzt13CKKYpaG5W/bW0XBK4OJham7q
YLj+TCskCtf/8mTm1c0MdTl919+bs+97ZrboOblHGhsTBJYDB3vNYiJl1ipOglRvxPI0mL+nxTXw
y9JELYqjEBtdOAbUJBTPUW/sPPSvC5SSglPm7fesQLHbWjrp+Ne0/2shwVejRNm40gN0BeJzfLHP
EH1iNhWrkw4xPrIYBLUMtX1Q93vvuSAsDlrZfWAJpYti6poge1pOEPRzkIY8nWDdjIq4JJtyBoJg
eaUiqK2Di2RUF9HURsE/6qnHiz11uq4syod54xvfzoGPD+NnooswdjFBWKNRBN0h1FhGwLWfhVvb
faiek7+BgzMWdYed9iA4Uok0nfEh1yVQ1cVeozXJM+0Jb2H5lUPuARPnS/esgOlpjNx0XIksRR3b
o0wd8lAOksvQnH9V7QHkvFdYxmk9SGNL+WiihKb3EYh9vp9hopZMmxDJp9OhwHRk5rslAfyYikUF
+oKmz5eu9V9PZpjO0vn1mnfj+A2OnlPP2ztL8uQu/RR/hHtN0zA+3J7/M+5S4WDOcnYCcdiwN1Rr
XcvxfN7k5Lx9vZWDN83rN1USZI/SSBjiQoXRJmXOg0Yc9EQ7RQAK+aZCUEvt81eNta4h5mUUqpTh
eDnapVABii0rIWNL8FhC09Ra5fWATfl7kfp2tlcHhIm2SnDKCxaF2W4rMWvO8otcFLMU3RL62lcp
nGdoGrlF/6J3ZK8rw7K/jLcndeDKfxJGSKNCIbmx91vVfXSj2db3Z9mSsHH05R7pUQH+CaKMyQzq
0bWhX6vcrDLstGpCeyY5vOCYjQ/wk1Uke0F7RoLXaohl5OiXyUs40Whn/CvnO6hKYi285N8NbJzG
B8SEhykRf7rTfJzZ+rfb6LXHNsYwUzdC2HnQKMh4QPB0B0OAmgFzTdya1U1yYu9KH+HM7S3udOgh
xxhEM3SJnAapFZ5I1S72WBOH+P9egKK8LKHA7bBOZ+NZbLr9lJkdkUmVD6OW6+6rS27Ufr4h7jFW
zKLqu1R9yBVPExWwWz9c6WUE1i4OV8FeTAYgmuJ5521DK31OHIBXouk9PxpAfdXT2bZhz4eoj/2Z
DYhJMeOeVGXAN15EtuQz76J+1GFjrEKKAh1SrilV03PD6IUspU0Tf8dJPk+MILpGhXH0sN1z1utW
XDq7qwK/8CscSDxauLXi4P63O0aQZrkBx3zvVZ89gtf1cnMcuiK1p185e0OFTz9BTt38kjof22nA
Stn8aIsi4yNkrpDUfXOcnfC1YUSXIWxRuXc27jmoQW4nAXiPdbvEbGDngxFCzFcidmeoYN278tt2
BE4ogEdWIddka3izztpYumP6PCa8DFaNEhF18BEMmxpIuJvpz4iVEmtIC96KaG6AR5Wks951H5SM
ZtapmQawnXgUAx9h2HdEk4YNT4/iv2wMOM5dx0i4NGFKBS76VMoshq34oF9sjZYdLEofdnq2qke2
9mG4FZvJglPYUtrdzjIMbGsmvnwIdrCvrkPhmtn3sO8wg1hkV4GmHcxUjJIv+WGsRhXCYKmbNupi
iVnkGQ0ZNmXjIxL1Pwomdxf4t6nUP/d9+iPDbvH0l8bcUa9IyVBU/BsDmgPD2XQAX91HykEhNHoi
oDRrw56X20t/Pbpqkh7DcOgZx6ZD8vEZyPPKHh6IAxg0EzMkE1+/nL6xYqBXvqgXUQuFefFTdSDN
ZAL10mGrelsVJh3UnrMI61tPBT5J2X/NZLUk0EBLfOpMFN7hSqqQgTw+O86BpedjwcFIHcR8gYGJ
vzPmzxI1mSL7bj6t1SXZ8NI+QyZp4QyD8Aog6joytTewtwCfbsuFrIVCdBnIWq2I351WRwp/5zKo
JrAHiY+D/pgpgnHjXS3mBTDDRB5Db4g4hL6Y07n57tTUGVhn+3d0I2gLvvHOOMgfLC0BFt3FwNOn
VpSEg3HRwaNp4WtYsqToV8DPKQdIIg7YMmiJhiryCzkPp+c0MtOP7FJbrJ4Jd6F/hZZlVKxQK6DQ
PxDdpgs4+iUGdeuU9jt0qz5Wkfl22xOAY7e97xDKYgTX5OkT9EWNYRaahEoj2ZPBmTIfsEcyNr5+
zJu890XaEpUZTNvv3SlPZOXn5wr98/wjrK/e7RdafFSgL3ze14XdJtEumBmk/bdhHh7hLo5nhLG8
a0ruTi6oCBIi8UKtgby+qoA5gGthA9Od/X9uO7TRneftWQzmZdN184twz/xo5Cx/XnC+qajLwSMD
YwuPFnr09nzU8cUHUbR6JxUD5hF349fh/R9L70rJE4gfcuyucocexqSA/EEe5+Re3I5zI72SeJZI
sFRXD44tgMNnJrJ6FE+onBXpvjcD28PT2OzbA7rqa0hI48iVL//IVfXGCNPf3s9vVf8YyycU+5hh
52mnBUnnwN4RjgqPS2AA/6K7YQ8qXAw9tr6bBMrQo2ZMzHCBfrsnhY+JSo+iGrH3CsGblEbAfMbn
empqqZoQrOOdbXACxLnQAuWXGRLM05Wb0uluriCiT72lfltrl1upunwnv3KNEQAvfeSmc0R/V9BU
sTm/bJww1327BbKvGmVDfTtJV/asaqr/5fL73CpMMTwH9bqx75pNTyVRcc8c8u6kIrcj6kfgW5Xw
Qk+XmIWjeZeAmTJExkN0Fd87EFbWYLC0VILQKwt83DkC7nTjSrXIpktDYWH0XS7i9BFH6/Ovnrts
pfPkBD1z1opTVyW5FqQ4QhVHQXsGKG7IH9UaViMRV4UC6/GEH6iozN6eZSsBUcSeTWqumLoLFsoG
VapRVQl8f0x/2j4+7BT69Qicv4EFyQVy996J6pOtdJ4owXvyWOdhMS7wWEkkfgi9LcNMN6rktrD+
yosV6XP3B3zr3SNXGp6haxkCHeEjDhAVqFOr+TgqBlrM1EgU1dSwXi6dWJT3iZq/f89Zz5+FqBco
xsLnzq45SOgeUOJtz6Tw75cKbGT30kgnILxWfaRw374Pn9LoRDATKmqGZ067Vwj1uclPv/KT43dI
wxJ8vx7XJAHus91T3yTFEEwCC5A9AKVNvLlNizHlDdUi57jWRVd6wolsiJTOUl4LG2oYim8IMtuh
j8LAzwd5Fu0K1U/StdHj4tdDfv+GgY7wWmFN9D3ZexL6SDMggHjZg0mb+lAKAKOyj9+c7E5Jymua
iXZ3juwj1vQUeGA2Qg16zHOzOZbv9juSrr4mUfZktVpmyVERd8PlSKNOB2wnwO6DALKFHBAN9UGZ
64LHJZI7GcwOKSQbjLto6HEBbvcbmIiycMjSTCks+OjmM7k70Y9OfQi0upwMfOLW3z9KlvWTjdSu
BLWp6CAe1vD8LiwjH9dRjF+fBQ6wbAHudBvhtff1JNSa9gsgP7DTXPDcJi4wEBbCGYJzBB2MR3oi
QYn57mOA5fpxHlacMQTellPDvNCD7xar6yAz6UalcuellJGSXPc7sCp6qxSjsf5uIFqdY2+9NeBP
93JO9xiVUKaXLZm/wFBlbaU3tYmZBagVEmw5bMuTRaI2hZBhD59UdXU6gnbsg1r9IOy0YY2Z8Mcz
1Hc3q8/1FsNv3JgLrXw7LyB5xt19ODTTzg7sPOL8CU+xFDcSMXU+qgdfIssjTYm2t/PESYeRa2o0
Im7wUbif+s2kW27QspA0kO5XBzLaueEPEv4PRjFvf8X/20guXHn1jQOAMBFpIT6Q0I4DiG6LiWfk
AdDgMVusCQD2uxbtFMZSa127DKSf2dApuO4nbUUwv9O+VBoEuTS8vSZCzGd6tJwFgeXtl7BDRDNt
wBJR8o/x72y1fHXyRZ4ZaIRdPW67klh+2JGeF/KsEPxy5Us4FtVENFrdu4plFaSJ6/wsfm4kRwGS
lnxU2eAdxbYdDKZrLSucjZKzbJQMm6ifi2eZJ2hhslTHe+fSl7eLU7fqBgWminHup4b/ObuB4atP
Y4s4j7JWvh8Ijkg6sfTFkaxB4yJ09UPJel+QBYfbZC4dmEodP2Tei0qeACFmEsu86LVPBaGj2jzV
iusUHi1xPt/P4JW7IHVQhmMHQWXmPHavm4FkGW1YWo41KuxzSjy+1zExpVDwIhT6VP+0onT2HXVi
+O2PlvIFmnVuCrmiupjZ0yOPQE2CrhZ0HNKBdq0E+wqL++jTAt51ZBVL4A6QjeTdyA7HCcFpQY8Y
406x7REysLtxaeAvdcMVqwXM3dW2/mfaP2TYI1CJURvmG5e987L4QccUmDQSyneoENVwV3DzEvzQ
YW/yE3oeSv+yF70Fvwy3772vJ0XPsqjAE1wmhkTMszvpHR4UmARwoaL+nZoYfIKjgvbhZFITQ+Sc
zKLE7SFD+7HmL6mlU7Lybn1p4Kh5cHs8zEdyhIzoK0xco7sIXf+PzqPAztfvO26BH50UammSoMkI
RB9AhoMtLB63wD7SWnaSgx4HC8ret2IMGEoCvDTF0AHbrUeWJVSuhHEpD06agdQAOpHbLhyqItWQ
fogsW9tHqDL0LGKWgVSIpHyhAwp1FVIwGDBMXRQuCEaczm0YvMECyUh7qWF5R/NP3BOhJXuQaaJY
6fcB0qlwUZsoq5yzfCW3TNwrIMdAKBDtaTgamU8uqYeWf6K0wMGNuRZLIlFORydZj79HraoJFA6N
exd3uZGvSA0ZwSM0+4v6WU4+JgOxITbNTiBaaxd5fZPcb7Wv+SBlHi27wvoZCg2Zew/hxmyXvYxC
RFrBKDFJNkp3lIf8+S+icrP8hgwNEeuRGEnamiVYES6HGAl3kkPkSQJWJ2MiHWnh1OMHO+nJNaeW
eEUB8gtZjzGKkBgIzVExrPS3HBxm1hauKNNavJTC127giR255lbycauNfGdpg1VZfsJ8/6h3jAtq
wAsZ2cH3ZEK5AFa9+eTcMx7jmWyhqT3i+BMAxlDCcUJlHM0fDcAI8wmtCiPtE7PldzwTCWdTo+Tc
MF6n0vk9lXADP1yXEQ5fdNU60kPCMOW2qA/ZNf5CYCawkR+JepCXW4kQacRbYs2WD5IWE7tp8ViA
jwllW//Jnp+YdI8JXlhhoJhJORA7AfwVibStZ4TL664f6ZXkDjVJ/gDuB1gGcMdEelXTCe7xKn+w
YUyAQ29NVZs9zdSLXyzpszTlDhmBCod0GuLL3B7zRCFX8ZnbSKz23c2349uKN7qfG85ztUyWGv3Y
maZdQ0x+t7ZqqSDOEtNfSJoKHFqTeAFMohhyCcOiM4P3ZOJCbbKzOsp3LnTf32wcuTGXo3/yBVKO
BCKmtaBQMxyeE5KOesBcowSnKmJqnxh4TE1RvkU92iCd8G4gOQnXUe62brL8mftClGezqTC5N3Bt
zQz4lIr6ZPQB4rLaD7luyaLwHSfvT0GK2gOhPb1IHOxH7QduM6yfpo+jcwhnWEcz1mswIiI6YPhy
Cam7PhPo5KQIsz91FAz0vDlVqXS/hZitWXInmhizFUz1ln/M7BXd39chaXnYSfTrtvtCPbwODPzy
xvHbebucPS7vyk9yXLufJYP/cjencOEPtGbH2a0uLoFxSXx2rbSrCJMWsAGHuP4DhZcWmW6M4FEf
7p53XkqxASWZ065VYy9OCdUCwQdSd+WJ9SQxqg9T1HxO5I6EAO6Kzm+/Fzi6wxmiGLGN6gH4Tqxk
oJQlq+PfiyHyuDJKdz4oJZFx+Ct+XRvwE4h6DrWYSK3VQNaUu3vjzjNdS8BKgElfnVvW7ylGvaIJ
0hYjEHWKtwPzr+7zYiGSISEQ8afXB5l4soUeGV2g1RfVSZX6CeiQe0iGTBF8b8Czua936ZR8ldXP
Ho9nOM8haAR/LkwCWBYngRjoXhJlVn4XUg1BGlqZ1pD246aUlSAXmjo4Pm13q0pkPzAt5TSgNzwz
hxTF0jxI+8Lvs1Aw5i6ohK8lLvmnpI5lD37PJ7K5V8WbFHHcoJx0aoptSb/cXfOjjEiGKhWU0UGO
E3g8HoSAr6II7YxbgJwNNCSIXdLlu3E7qU+LsLc1cIASZzRgrwYke0LPhe5Bt50lvMvEYbTJJ7ZC
7sucgqeJ7niarfOhVvORbz6lauvBbONLMeh4K6u+xSEODVh86E0gyYpwl8qboX3CI6wqEOG5HpoB
eRJoFKJCDiqh9KwAEs7XeFqVIeKYL0fr0YUKZU+WukmAokN7mrGkonhc2bv3J43zIbVIWD4r+QJH
mEtQC3iF9P//ue+7Mhz2C/Tcv+9xhE/3C4SnGGOd60FEg8X/epDVTeT0lmZ5WGG/omze3jSkqC0J
hl6BOwbWgWVET4XEAOMwao2QkvIfAnw2Zx2nxG8FhyPBVSbAzXmy8UX8Dv7NbNsWVFf+ZJJb2TGx
F7/jUyrv7D/aSupfAfojlPzK8EHad63ez0Iyqx6kX2Y/iONC5frOpZOu6f8Qt1Jkgrvs794ekFze
o4gBqc0Q+r7jTzKRVDqy37hXGanZAEDA5g7xt0Oc68LTVyJUci3Q9UXUNINdClPBqFWWlXC24Eyh
xbM+a0AKjj5ZjW8TwZCE3OX1GG/Whv3OPBZA8Z1AunQ7cEtxlaCBFeo07eElqTWcYpQZHg04LbZ9
wUuQRGqXeEnB91vcGzTrx6e9MkRNQkBldpihsRYLme5ycDTM7psdzrhdWJKp3lFuuk/GF8sIsjYz
VkbEUOzEtfFOenRkWDDBp9FBx1JhiEQA8jrjdxbcPSjYiMCvSfRk3R8tCE52VEg4Ee3piB+GqZ2y
K9K+LiG+fBA9GD2yF37ri/Ms0fhKLEJMZ4tabC+eHCx4SbglEHdGflezIMAEW7RdHHGCIErq8QIC
Pb7bAapeSV23KLtQiI8UwkICY61dtXIEVASNL5L/ref1QOz33Bff6eqRYrzVv/aoNz1Ogp2xpq3e
gCvciZHNVTUz7N7TbTwgM51wAaz8a8lIi91kNih/btspNewyqwqTMgW6PhgVL5MLyA95Hpy7q8qI
+4yMa2hmrMV0hY+mHaDZotdxqmXRQuzm11qoZmhfkHpfz3aAWuiYFzo2ZLR2ySuB/NEi0JExu9l5
T8SrsF3Q+KXg5GLtozpM+fEUJ/+IQRglFHkpEozgdxm1EiiV74rW4h6oJyRnBFOVX6wvacn3ygad
BvhXbpoWGfk996QkPl1ULo7R2VRapIxC0gU5PU3tJ14LnM3maOUaPc+RKHkc4r+GUcfwjMwiNpzz
LFj9eiUwwq7jY7c0IFy2sFAgNvPWezL1XwIvgdhJ3NXAwnHf532wcqkBmvp4dsAXGiNLb8phr1ok
7TXYerBLn0GDBF2QBD/bwbCj8vD78GcO9vUxe/ZS4K20ZfzS4zg9TpBcNHBWxJhQW/x5vmcgOMot
mwGHo1AKVpXc2E0trtu9TYln0m8SR7Ey7kF8IjN2iRunGH4dnSgSqiJEJ1i57xuUymRaE4Vt4BiH
e+i2Rd6B6mhbs2AVxEJKKmKk+lmBhxtDqBjmjRd1eu0YAHgOdKM0TLEgN/7irl2XWZQiQ69s9Yub
NQVuQ5HZoYEO0edZ+SduWvsBi3eS+urLIkVObbLCrF9j2Om2zfNrPfVcMz01vSy7Te5cU+gr78Bw
UFLddVmvdp1kgzmkaPBzRFwrPHRmnLl/e/rhV+irPVujoX50El3vXCy5ggNA3emR2EKmgi8X/scE
87cvIZmgbRZPEdaJstSMEy4qC0tKnbQQ6lrK1txe2iCLLjPBSqJg0A+ZHTXMrZny/u5UbnaOa8Yz
14khGON5OJwRgw15qqMhWPkCW0GqUNmH5M95h1dDntXhMTTPGuEzT7HUYVCyBtKDBs3Eiy5Pn4Rl
pryiXVLLp3PGi6vpV8QtZ1dsO08Xuo8fmfTXH6Wacj7bC6YuEsqxL7BG0ngCn9fPcXeFpkf8Zlt8
HgOpm4Uwtuac++yPJsuOlD5ixXf1MpsQ1Uq+G9DR9lN/gYUEg2ZMAZ/pukWKeMf8G9TwKG8kNHqK
Tf2frHcVidlG6WINt9cxmnipAB85dudGdqMO4L8Mq5Lg8wtRO/Ev6PDFBas3/UZqsvP34o2tbD56
vJKkBLhqcDausbJ90vh5s4nxgNSEbXEpbIZfwS2o60D88sUgExlR21H9c9G34F4p1yUWcTWoohv0
wL0rd6SEngK1OTsJByMU/dKG9c0+DP9RAPC1a8IaDfmGHXEn3Ps+soGrV2U+O40EF4R/ERYE7Gqw
2BU5UscKza4COs25Xv34J4Y8MiHQYC4z7NVxgBxC6eXpAS2d3nSHEpAsffAAymCKLk350XSHaYMT
RhFI7vqRhxy9tgysUK3w4jBTFkVO06PnD6oiDKbBopIIbrfOjKfOGQF61DC09ACqgTz+rmcwx9tZ
ws3wwOLTvBjfyTrp0epUbC395FKUF0oExtIafjUM7F2NSDYVLWF9Z/RguO7O3IO0fuoSkhgI1k0L
L3cYGJq3IIPLf8LV+Y2gz8WTFlbB8/KyJBtEUwyQuF8Wch/rABYP2WnRZ5aPa4haaRN2Nx40ka55
8upepGG3c4sD4Dh/zZzgEaoncXx9TpGgnPKycV52TLUJL1rPDCQTjC6w7hMf8YacCUbfTcwF7Ux9
wccaingOFyHo/3y9fYcREto2UiiniSGnpWxCaoT48SeLOPD/QCdHNgqPpRlB5sMwcdEd/QFIbMXO
FjOMPI0OkNBH+NGL8vMtyO4VsNmw7t9OkQh4d4ZPK66Nim1o8c23hHj/YB4vutMZHM/rxXVr+smP
3UH9fETZUEhrW0fwpG35JpFNf3joEyj2KcFhp+uJVnyJ6XmQF6sBoohDsFuhRqAgxJGdZD2NpN8n
WIJfTF04qePEGbfx8yjagMpdpbM1+wgviSpNb4ojnUvaUWTo9acv9NGRGY23ETXdVpPVlahtLbSn
iP0HWwqZ7Dd+yAcsuivQv39fQmUgYroZ0u7g+MT4pUKHV/4MBvnzjbEA0WU7T5k98iS1EWmKXMmI
jnyPmMr/uyrPlduvTBYgtFGKNcV0NV/JW4mjTwq2qq0LWmpCdJrge8tQPSryZzPMnYSmiC69KWyO
MnE9pP5w5EWf1swxbtvL3XrIfjNyz8YFPEx+WdBsCngyhHISm2Ibw5QbNYe3U/0dS3xbTuQ5IMOa
4LcISbk7If3c2rrt+iVH7ukXMl2JCUlpOFx1euc9VsDAv+DVxBDDxPdRsrBTLUeP3ajg3wRcWB0t
TbZJZSF/PrPEhrDYuNGo78TDsZ5oNqXRCCajDTbWpse9SXcjJhIQfxJhDBsr8XvR0W0ZulvUnmR5
wdr0l+/Y7pNHRnIQ4Omq7AW58iLhL4N8KA1G4uzhyHCwGOcP4bWyZlLSmtF6DNpeSK8uDPQ6Eai7
CnJHEzKM3v1Ih6O3lWK9RaylGn8cL6kiIR223ZmutuFxNYbI9pBgUXj3mL0VYkLuRxBodaFu5ENm
8j0kCUgwNfZMSl4l395MK+jam4Df0O+3+uyKsfAbhdNbSIXUiPUzLo3HN7fpL6cE6i3T3phDcr2W
j0YvIRD2oSei4YVZsUGa0+Z3DtnI1bir9MLYX7LVCGYac1ZL+Y/Z/gQo9jkg64Sif/GpOGHr2Ic9
zPFS9jrOtoHwavNlK8DoCya10yDZ37Rw8pRH2UzJm7/z2M1UAZJylUu2y6GVXvc3DqPxxRsOE0td
Q/3dYH220PJmsc8LZX+P2FeSITFstI7p8NKY+J3Cdrjisu+7nuQ3Vi4Phxgvm/To56oOqT9ck1rS
Uj9cy/I1pDPtfFJGhTG+3AVRN1qfgSyI6gguvhK4d7OMB6IfbCZtoSY/lRvXgD2OvGpMIQjWbxv2
ZgNmacW7aVzKtA7uxk4LD3/ILwFdh86b3IY5Xu/lXuBcqV9UBvUziNdaiW94bs7kw8akY8PCvkmm
+4Cb7a5B9CbKOI99su5bpEYps6lUwO1sk4DJMuKAdOolshX/4c83iITDknYGrNlOBPMuUNRRT6Cy
ThSOfyjnYilcSJDHQqKmop8J3ArIn3hGobxGCv0AfAOeORRf/s5LpGm2sqYvBVvicP8+r4+Tbgk6
dbxRyh/HN3aZm5dNWw31ZGDZuQcpqPwtzAsnO1AJWzTAE1jx/TAqlMGDYih0QZJFMZLbd1cH4yIN
hZFQKenqTsGSHDyZ1rG843sJRss6BOPp01wrgq7vHKUD0ZBEef4lBG+bA9vUeqDLa+9L7/EZqcBA
yW/ZoDSAOGK1PpBqwzorvjRGMoAzWmc1UOOLQSdO5plArNve/jzsnIgsyx2/NnHnNPfiY7JKkH3Y
i+WN0EhD1jWU8mjtenn1cpx77NXajvs4Ffgflh//tzZYzCiM/Uv9HG3OLCJ4SQjyflJDyucSeJIO
bovQVEtr4YJQ/bMbfC8MI0pgh1NgyoDAvjr/cJCxjBsGWKY8HWHq3HVlpWRvfFu8ySbVd6Al0DNc
NUPWXhF0DENh/h9FLEhXLGBBQxWk1MC0S34x54QZZLWjurkNSongDtl/QdODbG3cQjfuvw1FXnok
IDQUYOn6Y9Gig4bpTaOyQQ6YmQCAI+NBtRfCrCthf38rEmFSHKtiN6ahThuo6uFDvusjnSnqPEG5
vawD+cYGXP6S+mxKduYTyax/FwYF4C461EuNvAiL6xnLemnhBExXLKzGuRb+cX7mdnMO6Jw+qNvI
J2zpMBXbg1QOwhAQHHHy9lRlHUMmFfROwcaQowVguttSHMUlCpcXWAlinMDyPNMQ4eowiiPpLFdK
tgr45IvGIlss1skdcFPOWd/BunSzFdjWXlMh06285scZzAUuIaruhZadg/9uYfdw51IQ+AphG7j9
nHwUCBNE1wAvVynYbs54So7BeslotpnnonXn9I3PbliRlDx1IMCYBZPnRCoWkj6uRR8V2QNfcMr4
uR2PpgKYjEAu8RdMaBWC2qpLs0iUw2o6Cx7tnurPsOH3PZSXCtdfu2KNdBXmhyqgiV6eQLa64jf1
Tf6HOO4lF3HuTI+78DI5DRdZg650QLliIeQKdiCH5EwDTQnwaTde7tGTtkweUOcPBg9RAZv2GQmw
yYewrFNR/RgFWHyzbvlUh7bVl2qjTyRYOmxV3MbORdB3Q64QOtFANmplPFbFU15cTLMGhj+oilqF
D8+prUrfWaT45xZ0PkWGEckqZgkIRwGWd549pxboEmph7rGzcQ/SxLjCbEfbEJQ/xpQxFdeDezHt
xGT9y2kdmrF7YOBqZ78ett7bezQ2QLX1rhJFjf3ZORiaRp3v4+ohdyZmfFIAHWlI9uzJLtMwA2WF
YUTmvYDcD2EIkpKwSSRzLEhsPoPHPiIhycmQukPtUKE54fHh0ctOSvicTEk/QkQjjNhUWFH5wfby
MwjpNuNTIDwW8R2FLE2qlPjnMoghj60HsTmxa94XyVvyGeqsCRWKbgVxnJo8t49e7pZ3+adKaXGn
9Yewd+GzEngeRlIFpfaOliw+NbhviOvhK34nX3DhuXjGPWKkC38q8ZlH7tbu/yC+sr80LcF9Uuk8
XH6LNNgrk8IreY7J/lCVW89FVuldHZSYxsvXb9qsQ/e0IjV6L4mPQOQAWXJRoJ3tVIb03HQM+iwN
pZjc+nLHlnKMVFCc9tl4mHDweP3FySzgHC+efGRhMuczepeaB+VTUsbgfv5rPgoqT2iYyIudHRrh
0w5aT7JVMeDCyG7qp6J56H+57gNKFGTNK8AK761JGnC6zhkCNMVZozOd6nW+nZS9cWXX1XpaJAeG
H+v0fBiRPXZMlQrQEaSjjYOrkmqPUtYvEzHHLL7fukOWDXqh3bZj34kGed6sPqF5OK6vQf66tAkM
nm8+XPddzxZ8n5dp37+539qn/5WyhSxocrFlCNlsjdTHEKkPU4DuBgY4fyMimmi4Sf0APEaudSaz
1QZ6tEFz23lFVwI/alpXZ64/ZoRKqodjyYNT0XeGNgAD1L355E9VOrp+PdIVXzLkqWEqaUtyNuGz
SQgV6Sh/o0e4+95HIuTHBpDjbsS6ePTOcql+nz3oOF8VM7jFi1L6e1DEd5GxHBz1fQ/n8p+qHkkA
t09hfpoXP/XP66NlfxJ4lmwjnUil3x8CmQfDG4dNFZXocD8FUkndwex8WcSUUEURXw8oPlWzNzLl
0ex4t8OguYpY50ZL7Nnsa37mX8aH0VjEL310BtKTaI1c8fNxaaQfLX6XE5+ASfIbt4nLD2oUv0lH
NKk3p77MFlov7u/spjycdCbvAJ7yyXYC0cwwC+dzjQjKfTnl5Q36hxjJB9YxyJGbxhvS82cJ54Iz
LllK9i33Xb6Q7jjzQ3HK7kU8Ah1EicarUkytNSYprP4DM4T8M2XXTWff65t2pLD72J+FyByXC2Ig
R5bJSjnTZ9pPHGIHzLRVzXOxc4lFu7l8xEfOxKDbBA/seveP3oNAV8gZTp3Re/Am7NSAqQxcBQLq
Zo/3sME/O7txmKaXjvtYQQlzYPyNTL+hAdq4Q1DPcTpIW4tVJNlDxd7oH8WjOcGMSLxxETjvEqNd
jMsGZJkDKgq8xHplU3Q6eyEKxvjWI1LgwEs4a/BpKpjeGyl4iWOOJVIY7L70TiPF6XxwRV64iH/i
LlaMcHc3/ExKLXORf6WLVSZcrNDJbXGIX7LKtrZEKufxaSsca1TzOvK0vCH2arVoZe2w4GMcCvOc
aYva5IPsGyDbXe7cFFMjuSxDYt5JzTdD2Fhc0TicApFrbUDqTZ8MXvELMus8OUXluUWwEn7CaSSm
2mnd7TT+afI4Mak8eFUoKaw90XhWHyiZeG5m5dQ1mj+ftMzuJpUtIh49sTPdQ00NjNm/Cug+fqqq
gXNhmDChWvnH6L/U8w6qbZgjRuUPlBraJZKIhTNJNeoBva3xooooHuoZVdMpVmMwLwITvObzR3gJ
vs1ZjWlyg43iIW9Sg9+tgIK4X+gjC07dwTf6DAkUFTZIfO3jT8cjdgsNoMt0Pyk3vEirUNxyutJB
QB/RZluo78MRrEEeDm8HVKNZd6HCjdpL4G88rkFJC4qiKT47I4JfUwCjnIz2GevD1+XwdmSxmhjy
SPAbtg0um+oR8cnxAhOSA5+mcrqpRXKi1q8sYR8SWjkQXfd0zVnwIAFny5++DGB+5NteCVhjdd2F
7zCqLWfDHsLHQ+eSQKXbIstmPLlpyytgXY+7SHJaEyDYyY50q5d+fHvyAvMuBDeXT7pjUv4Hvwbd
sih9hgbBmAfu1C/BMWVOAcmL8gj22H+6EB2/p04YC7/1yphtidxC/fHQuJu6gdLjjaGlyt6m2jTd
rrunuhhZTWPhhJ6RTrzLEjJOXldZuOkQoM7rY7Zko5qCfT3VICTjgCIAV/9OhqM5/FXy0fJp/uJr
wQLATKWKTOYiPQYvAelaB5MvyK7auIZSay/qEdwtRHNa15h9k2GxTKQTAV2e4O9NlnkghQlyyKu4
nYulmkIf/6hhEgGjArH4H+pLMptXkOwll2SofySz+zapB0gNvJqU6BVUiBvRrclv4xH/Pk6lISQJ
XQDxHp0h1tFyDdStTb7XCfn7+7F5VbfPE2PGE2wQlwEd61D41IYUJXq6cxf3mhVOoZzCJA6uY930
2Fsg2nHswAMOnFb0PLu1VIrUEvYOUjBLOO7twv5RikHd2rU92bWUnpspbV0VfhMe9fX5u8YzdHs4
N0xSgBTmxYz5X2MtQzRIHcNlfBxvh78wgRN8/yFEXhXiqL4ZT236V4WAaBHSTaH5TCZh3Qc2hZy2
DaYY4Iv8W90ViTI5JY//K5521pM2PLzXdHgv6mVfY/5v+MtO88KMNC5pOvkB1JplVwI9qP4zvjx4
EgUUgSQmRLCV3Zt+r9ugpoqgh2lB76+BSnRZzAYIdygbD3K3eyKAwcoVTYo+W+Dz0GnwbyoZE3hZ
Nqy64d6PxtiOaEZ6dNXBFAaH7IuT71WJoqfuYAQ/ges5LyffDwt923TUZ5UP6dNEY1ZgG6CUKheH
pP0l71VSYSZxgNGw4d1LVBhLfFzkf9mB1HHmL8UHCU0qfBdBze2EefXP/BpmZiDVElBlSMyZElnv
2Q88CDFioksJN6lOWsX2sgaldizvCtRSXCqOAI/rSAG/6c62z4z5rS4r3Ya4Z6MrdO7qMmW0sWlp
Fl6Rycqvxdv+g0GCMkYhS+Eq8OIbQCpJfjLIHCrCFR9wSgI4nJj2W0pibcVeC0WxiRgikphQijni
i6WShM0kPo51fi8I1yDpPaZ5AEoWI/onwgAkis30yqnAp3pmbj7I/I52v1YUh+ZUEjHXypgh+DbR
agOHv0HEgXUzChrpq4hSk0C6erabL8yz1fU9XpKOEflPGVvjJvBu4y1zcA145uIrd1tpiuoDWVs0
IOZFlnqf3NaWj/FvzzsMDlB0RM76vgw0RwxMX+1oQe7hjWlNn76Mx29zDCYj6CfJgI0de20/z9/O
VWn1250RM7jeVKFUu6yFtiPRKX8UrrO5ZG73f2Y9ZG03ztrX1RyfHYE7HoVabsvyxkv7r1bsxcg+
51SPgSSeAD+y9rgUE0h/o9PLZm4qmkMcn5S1+s+iQpbWDfZB55KXiTxEkQEGwUdCc1RLqpaPofog
pfAg2Sxcbbkz4cT1cl6g56nYtRyjQSrwxL6uXfR/Hsrzcabisw3u2wNM27pBGllw/tAk45UUngQI
dCyT9rlG8Tal+J1KDaFSmVkSunnB+n6Pb1OzgkWlwiexCnftusq0reMkrfoir32G5DhXHhqaNEqi
xZWsi5REHyXjPiPaB64lLi0PxKGrTODkiDskDvgkSMNgFDClT1FX2WM9u9eBLba3VOE7jHUT8RSf
eeI3Z5D02mZLsV0QBQrgZ5+5jpVY6BKlDg08VjsP0JAlBG2aC2AeUFiYWCwNfSs7wqxjrftC7Lio
/Ko/ImOXbn8DXu/2htQdv6kdV9udR6ojJEVbB3dkUjAUk53ZWxmsCI4Og21JuF2aaoTiiPXkCQei
3HX5VtlSdHPCaZ6UPh3aICYDeDE7GmTZ1hCWR1b+fGZUmjaxMqFPuKHD71PamZ5lL2+LTRieqb/e
u0KS55Ee37SayVvxzmzaWpoRBebzfv7wLilwMrZ4Sph0B6b5BNFIBw1beSm7iS366+CuZPHUqFY/
9ejq8JKQPilR5h6udhWWY5vyWmEMhMVVxFDyyNke59CGrtO6S3XoVEun/95GjAFlfGjOOjG0haeP
nmJVoRYcVMKsxtd3KmPD87C6y/03eVSNKcju63yPNA0KVVL0R7C1JYHAnrNeT9vjsRLo/GBzoZeN
QDL/Cu+C/77Lsv1+NPXyStEnjr7LlZvrA4IzyUKQipwyHkB4DiPmJzcp6UBBZRG00t71SLous1d5
NXbkFVbt+ttM4HFaxjSg6xFx6esbEaDru3s9Mgtv5ofkA8WLsLTsFgoiOnaMkx5WXh3mjIrqf5MK
k+pCQoEmde/Obg52BD2L6dtcuAGcYSqG+/6JUWFNn08kDMQsdj46fMmS0rpFgNVJ1cdTMYPetd8w
GAusumGKEjrJ2wwJhTIFOPaYRqOX7NSuAKRALm3dE+VWBdXBofuRDEBIXFdxjvITZpRkVRRs6LK+
YApN7TGcW38iNxv3nzuKK4TDjL087D+nc6P21UeW8KD74hS5ONzmbJsAO1CZZ7+ikgTIcXi1tlmh
HVhSmw74yt69h4biJyRB+HuD6aaceEb6M5uFpu3tY6JUgq8nWzoErQQYRgpQp9ZaXquzw+MXq8RI
2dLM3xEZ4bxd60CvD5kmjLNuCyn7sDH3VG6TmD7H+tBWw2LNtJgzFcGauVz8XsrDeACQEkhH7WAp
2bM5kJzOF8w8FiiGRndTz4kPL5BBrRiuQ+G8P4x2jjVGAN1jWOp6MLFhBLLTMh2hzmC/FOvxa7Rd
/4WSIqnR78w0I1iaKbsDYs3Lqu2yh/06LykkmAKelb/AogEfuir1i9n10U/LIvZLNCHfUmiBY9+m
AdorpgJNNGe4Fin1bXDx78a1jyx4lDzOZGDWPs03o9m41wzfkQDVzCERjDfvyvNRg7cT19BojMp0
Oe/3tkUoAXHBzyX4ZiGkjiH6UvhOBencMeNc4RurI6N3QPXfK8BZJsxh2BVxRzdD0beOu1LRn8wi
T5vSvEPsVGtU/LXvmavEilpE46T5UgdAk7LcjjxMRmPXrRfD6/0FD0fyg4Z7KixDWsB57PnknrNB
an1gS1aUq9zkMe+lSCYDmRhTrikBw45B0TBWcoRhW2s0z48oa0gZz+NFORzl+YhOWr8COaccYrF5
SxLVe2atO61KmGKR6Okeviaq8i22c+rQ8Uu3MOxy4sj89nqegilIMGN9jEP1V4yza8J7tZ+vIcoB
YTlkUASZgNcER12LBRCQCM6zVD/yT3SSxV4C4BNPMwe7L2Rec7WZBZhXQj06q+wqmDDV/qmBieNl
VjvKHSTl2gLzzkL6JsJAI1P0oNzIRGrFnUwVhTsCToUAANRnVy9hSViI+HNPt6orccDhmBEhvFAw
xY0fmcsJpRNbGJhcILungnU1n9S7npRMYfBab+b5HeGwG/5oo1p08TK9IFA0qmG/PNvCb45Z3YGN
WWb4KjBsQl3MJN1c3v7EHSbUqU3+894L3aXxfxiRganmH+5Ouf7c875nM8fpdaqjlTf+D/a2hFNO
yQuClecQHCLGeS3JNLbBYWPpcAqaUdSuxKD2ul4bRYVSEdKlBd9CT2S5cuLkJiWgmO4+eAsVPlE5
vOsDBLeNTfhxuC3jirGt6HNu7xJtBqg7xqxC+pI7701Yx+3zIf2wH+qJ93wCZtLc1x57KMY4/+rj
eVvSntvbHf5fl3mmSkxm2i0H7aoU8Yc0Sv9yIRQl5aJL35I3mOAQzM1PwLSfoFXHS0Tkb/hx6vxO
/ZbTLYmjcSmgG368kQLGVy/hLVik+11+JkvNmm1H3pKj7U6Aalrh8QsqcB+9JB+ohxACGiKogCPB
N5lAHyfMJ3nBCUUtG61jiM5jQV8oShlZStWYbbacPZKP6F1AebRfCw0nIthuuPairdQlMg5DPgeG
du6b3rMsciFpqLZPV8BYmoChKBMjSR0mxSvMArfuKLBdyq3h2nPEat4iAfYV0ryfnxtoa1VXJ460
HkJWlXk+vwqenlgtyqXhMjom/wLStogG8Duc3UaTuidZy02CokJcN02lO+ASpLOX1r1nVF2uBRxo
AQLPtZ02oMEEFfMrb5i47n7EmAhWH2sl5vaTtBBWiTr9n5FE3spSpRIG0gNSl61k7cSs8lzbgEYw
gyebM0G58bJysGjTJ2xJNAWK0Wq4xdvgMyw9WCDT9tbxVbzUAnj76a6PVXgeNBBf3hpIIqf4d8A8
0xSeH3HGEQEXqn2zP/S6niYaOKD1cfuDkAwOJK1MSEDx+VJWvwXhslPaxE0/W9tEzgSTqwqZCY5W
68fk7sHkJkkvDqvxCzqgEQoN+0HwfMS050QG2oZIfc8OqoOqpzjE326ENj+EcxwpxB8fuj6oHKUu
Y5tAuEKATlZJUu2OzjQHLc1RVE7fXxLLh7XCAceqD3w1YbZNDP8AnIu9u9B4Ehv3So32Y7Qt+BNc
BpuID4szUyNNVSPZxKvbKfO56ESNZTiSs9tHNy79qccNcqMB16AU+nvx7Sp7g2Bwfthd5iqHEirO
p2cH/HUunQVQBGsLLwqRHlhppJWquYBDRBal4vgyvTDiJ02Zpm+qYWQ37DRYqzaWy1wG+R7aMxn0
uoFRh9KDYgPKT32UZRI4lh97vXjX8ZR8H89lGlCqrxYZn4nmVrTr6Gznut+u32aP3i46/blPSiG2
AHa66TeiDySYwG4TPE70OLU+tqbKzYJAY17KXlEOmeAYQSVVtl4W8L9BJlOVFO6/5CHmcuvKhLWA
sN3P5DZBzH0LpfP4Bgz6LYVa2GBKOfxrVZGXaTJl0fabMPBTUun1vJANpdFeeTpHRJw7JAsVWPsf
flDHAHY7M4QKzP5YK0zLYCP8pJ27X4QE6V8GNbajRCCi0IXpRax7Xyu/QdqjzcMfa6yaduUU5/Nz
6cvZJRnGf5VXLuLWhWAJ5769bNebWUZws5X7zdwkmqnvo8NDaxsK6L2NPjf9XJ/HjfEjpgPZmBrG
qtj8DBsRQylYgjNQ0xunrutTkR3Uu9xptFX21ff0O2As4s5FDfcW19S+//kDQGjvm9tFRFLocUoc
qLVrqb3ygdWoUM9xx0+YccBb+JIaZ0coaVNU/gdQPn2G2fxRUTlnNVArvDa+NQHkbkPJQek8t45i
Ong4JdymUpNZWV8Hsp7NY2bQAEpq/nL4LfkkUTk/coR45LrehXxnZpQnamgmJrcy3lsztajN5437
iOCVAviPm7p43pMNRhxh+r4QgR7djrXOaufR/B6VACWfTSMUFuueTkSdIu2uM9xBx+G9mbhCBmV7
f1afXZrgfKgcGU87lgedM5LU0hPXfz9JvtOJdwkgEKV1iM/6LU3cfBAPKt8ciL0mkwBiKDQDrgDU
XOPPjdoFwCpR0r/rx+HkMOe8J2G57SNIJiTQb+gb8yhtbc2K5+Ok+Z7eNF3E63AZXzLQkXRTinGy
ad+pygMmAMR5DzneCp1fSurLlpW2fvtKh0cY1+59wmaHMdfj7kdC2I9FsqLPjudIWI6t+Q1uhjld
kNv1uRqibqJGboiMA+MydrNedMeRVB4a7CpqWFjxhkTiI5CKmzN7WN0c1D5zJH4T+6WhxuX8ySNR
ihrwcLWkiz4oQrTj2bP0qZeeAq/YNeLniiq30yG61qoUWIzvzzScL+/sptr5SSUa2ZHeZqilzX6A
dk2Mg0b9zblaKW1uDKrSEUTPmRdGRK9dArXPZpubrC041KKslGxaROywWEnfRsaDsHRZ5+tmgCkA
orNvz1VI7chZJv9SQ0Spjj9BtQe+b+NFahofaU3T41QE6eIzVa6cPwvPfQEkdyVVMu4YvLNGLcjL
OH0y9erRTVek+4KlGvHNL5chS8vHzwiZUlXMDfsOdQg4b939spxggdJKcNxVyHWoPePcjgPcyumH
XSBXbKuUtdZ9ih5UOVElsSKZ6QS4V9Cs5S8wjoUxCZOIaEFr0tB2G/h198zUnUUSvC1yAOCNHWFR
N0GGec1Sw4x6P16OAZvzIJZTxuEFpHWEQgNzS386iAxQlM9y9NohSzcQapqvSDs+hzEPRluA6AFc
v6LD2Z17oTlWVaaagnE/6gnub/P/QV/s3zgZ5f3K9T/Z2XUZr5MpoIKU76dDKqNhu5UK0BENzFVp
waJVqrngr1J4bafS4wz1v3eRqAgrUq+G99RaFHyITrX2uyPoIrpg2OXCtCA7G/NSFsRbOHw1jgxB
7K/S3lrRF3bzEW5U1xsRVxs0z6UCAnHeNiUrgSyEZHLw7RN41n+BRdxBcRceU2gFPexv9Eok9ioz
woPvsBmAANZR7y/ESGvEATx2+rPuGAo+Ub/skTxVZr+Cj5yXDNOuJyKthHW5SgW/4Z4oWeJ/w+Id
KSZxE1sM4KXJhtzwv/OzhTwOL+vkRtOqK/WYyKk9n3eGKd4REkySzIBeh8hXfYZchoHfkatVONbG
UL+S2KkfoCOrtMg7sYsLAd6UhwOJsmh0h5Hojv2KkPDsZZIabRAeZJrKolDb91t6UvkekU0uVzcJ
2bkUTq1DCh3RBhjxCX7ks7hIaLblg75yaBqbXgQu39MyNzCgIDz93V9yarBptkmfJUzzfR0FgzjB
1UYCDJ5NZ2nbsGod+BmnZpMg2OnvIJhqCmSlAyZMqFYiVNoYwLhItRlYuM/TE0C/voC7w4kSOucE
CnW2rqEUr3AflkR2BgTPxv/RKgWxItZ47RoBGbkTM5HM2BDU8AlOv0DaO1i2Dw5UQLUltl4PyutT
cHfA9QqcxMhAwfTA05PT9AeWo74FMfwQEkM8YvNgVzX2KyW5QaoymgnqErtq4d9SrTZUpBgG4SYc
YJg+DCAaDEmmqYyGTMnrc8COX/G6GdV8extNyi7W6jv6pqewyLEDJorIS+yqpaJJbb+hzi7TwWN5
+2jSz8ZasbTEOYgThmLR3/2aUwWGlmkK/Yjw6NvLtn+A7pdWrLpjmxlRB1LUwGmPSjKP216MjPYn
5A7P61ls5ec3nm36xYCV3RiN0jZX7XyCJULmSl6MEmpAA5coKZvY5u78siavgOJ9c9GHGRVJxixy
mGvxThHArbwG+vGRIwJsDk+NRs7s+ux6QZcQm3bHt1H8mNellGkMzoVnVGxiQMEREvBLHGz4IMWN
P3bAKlGPhkhI6irCqv1Hk8ToK7GwCcLGa0yFUiXuQaSdI82zzflNLfYJO19JI9yX7kVVanBt3M97
rgb88+Bg4L8OUQGerqKRHMWP3aEMH27eGPMAl+hpB1AVx592RbTUvhhYFVZb7QFEjYo/2rrP4/qr
0YMiObt0TPi+691gQuTgWzYJzMJEmRpjrheu1ii6sO5yUa8lq73022JqLlEiS9PqZ6K2dIqzP0ee
PGYHtmX1/WL/jZKG0LZLdZrd3gJzVoAlAg7QTMhpKzElWYCbdznFYe5qN3P5bdIypuIHiGqWySpc
LwCszz3lDZzVue0q4VNzLbrokcgSz7TMHeds6vyV4KBJMofUR2lfR90iqPbsnkyPi5+Ry+i2aZil
5S7zLGqEmJ8n/RyWJdQ+bLsINcnMak+zUvaHZu0fqAC1z0jVDK5iECyTqS+MeF32+iYXqWygcZco
f5/hvo3kTBJTT4AaYOOTL1o6vn0Jaea04XXTXOABSYrbR02BXnd/r79I7w2M2A5C0ibyo8FGOUwq
mltYkG9o2a2cIDvsQ7ecWyoEpgOrOAUIKGdZWnUy4PEm6nhUJmp4l/v8lw3SV1ou+Jh+FWNDKih0
WuJCewUMNK70D+gKN0fx3jCnqQm3oLOBtjhu+rZyjqLJw+l2LMv2z6YeOKtXsQJWi73NZ1nM47MB
dtzVg27BUSeq2XCkSdb621m4iQ1XC1pIcSjauF9pgeX+TwN78+RhrrD+bmLsgYS4Zyl2q7qXgzeZ
DVtGKB2tIn8KI4nGmvrHwPFr2ZxOgxwIXgI/YxwaaRZRKcXxtRMr4BQw0AKisScBwVNbTSFWZtpg
cY1ysnxiiFRgO62vFVL6M9ejnPxPs7ConOgmIKfM/8j4oupud5ptpPc6Dw8kG0MfzDnt5Hyen1CI
csC37t925/XnX6aND5QpQb0vTSITmVOlnAp8ttoB3XyBs2jhKb1rFQXcs6oQ2Mt8LmwZdkX1Q8Tz
aXyJUP6NXfTb7nel8mETbbHCIZGTso/vbSFPa24sBvJZgmJNm8tS4UUqRDCVVD/BNzo4teA4WWFV
LvMmmIuJTz1VabnmdD9Fuf03AxT/z9Y9kYk6jB9Go6a6L9qocZVxZTdIFXPyJZx/6qifvDbFV+12
6/7mEXm8SxUPaVtmNZm5wb+LuF6zsHnouLYaY5NPQ5QoAnd6Q2fpBw9zzl4Fze8CN9mwDurgyt69
FUJlQaoh771WZckDzKcEyANN1jm6Ng49f7o9NJCxofDdI/ldTO6s5q2QzJQJX2IINKf6mbiILtYN
sCq1JHdHSNhscEuR9uYI52HnLdfkz2pkcDipo78ovInCerUYH8YrAl4u0LR+sT9SG4o+y3JRgUat
U0Gy8y9oRWo/gDDbMSNLsRvwwWk7ZUDKeWDepG0VwrfzEraHpZ46S4laX213AP0wWQ356wmkyUCq
/pozwQ75oa7Cz8R9DHFL7zRNAU8X8tbXlSA72311zsJl2KhRVS9SYcXiDBiZaaXK9/5LEjQ0ARhe
oqvwUqKR2Co75dSK3Upg7ehRWeEw5F2oFnmPGhn3IKtHX9TQZhOS8e/ZVA3c67Zr6XHzNb73ceeI
XPGh66X2sBfQ8aG3js4fWChvPywoMn+47ElvjQoUptuDuDSdKfW87FX3yYSfVqXtgfKjYFRHF3FI
wwdCJm4UdiyEz3zCFI7sFMaFCkZk364Iq9GX0ZKeDN8qaOE4fRkQokFY2yrhhQ0quJ588Qif/TC4
j9L13tlncEWuuMjvC32wS5vCugfhPo2dzQNDlg3EN3zYa9NeUPkrN4L9riM1HoTvTCl0kdSb2PIO
x5nHQyHHkuMRSj+Yje2w2hhrPlWOO+6LYBwAo+5be8U9o1p/Fb5GgCvbUZsFovE+BWU4IS6kag8m
F7mSIrJa4/9BjqTnNK9h+56Xy5CW/9AdOccQAwN/0RVqMsKTPpivTqJ/KBF/5goUIhfH9TZjcusT
DK5RhJQdNMJLaJKPhSwHF9bSXXQaf4Zx3Nwc0zytOuq4sL37mFSlnBgRWhlrShNtEjti/EMjo/aN
3JjXShMtWvsUmzA7uZODeRrTb8fFVO1Bk8YhAidM+0MOianqWqW04MCcx3OuEuYbO28iyyD641Sr
w3owe5Od6G0BsxTkQOl3IW2ABh1w1rXw/gr6HmNyOw2AftLzFHKH/2+KEh6PiOub30SsR1nV5eKg
fRT9BH2jmyTUbpnqsjSwOlZjHi4kY0vQ8AIL8eaNDAwzL5aRDXezOnryz1GeOyykF7906yyTLpjd
529UfziJFh7P3OEq4KlLH3m95BgpDnsYxQNYRmAVW8a4bFQIMoU9Ns49xUeXn3I1az3hnFr1Uq1U
5dCMsLacj9d7xJbVjUeZXnxQZHsxIXNn1bo+Bpz+1bWjlm9KmPxIYY3E0Ekm0U49XDQxcewDk6rc
0blVDR1PJCPFxF4tVzX0bFik0IKDMNEoJ1EK49nlDZWiKR07f2oCJduY/o1K4izGXyNhTGz9ym2a
iZxmxRIEezTBm078kQ2s20iXR1AqWkX/xNlO8WgxnAHX9o1htIoQ79D6btofcBYJJhsoSiWKT26n
ZqyeyVoeXIrXSYCPIu5tVoPcezj75cp4hUcv2Mef/IPDde8GoDULHR5J5Mvl/oRY6OCTg9fkSuuI
WMFCxOVRw+YnsYzKY3G4VZ+ibUL45RslqgLB6PKXqPNkcl6GlWWH5uqU8RucvjlVg1twE0JL6P5t
KRe8phA+dh+aEIF3m4/2EUliwyVsOKEo5GViwTxp/oh0vNPMJMpXAeU5n8aPxTPrhaqvrEBNb01t
wNim5kuDTqbjaxhi3w7TZ6109jpg1y+GPsIm9pN3bQ5dWKE0bTI8vzLu8Ejmcmo5ge8xRGpzidFJ
VzwG/u9FvBFqrk/h9DKGZomrYjcJ4bns2G6bjJarPW4xanS6YlT3oT8C4S5elrIdew307hB/31Xg
E5CD5MW/81OpoGWDzqhI5rJY85+FPVb3vqKLCrIkzQCHA0TTPfWpLo8p2OLXK2In4BImUoIHWOX/
kGb6oJeC1pIcr9Fpku65RM9E+Mb+XVrBhP3/v2vAf2elPiMenCEdcGQa5DZq3BJ1bHBsVWRLDyCR
mZQlJtC7T5eErKAqT01GP7qw8v7hTiUyPDc+53RPzQQw2htXKIATxd0o6ABDakzfxvfJr6OI+CsD
qKdgz32crg/Oqy1kzN5EHDD3/ZAZgdS7ygxCavgmf/jUCJhiLYLyd0B5Lwd+850tea5NBpl5PaAw
0jIbZ5+oQNlJbEiPnYEljPVXItLQ5H3cWBnUL2DaBlS0qsWpR8Img+M4OQasbvHUgX2SILGdvtvX
ymLK/OsT5M94s9w+hHK8LC05XxxMzynUkWOx+XP28zl97RirBeKFIZsbeixnINZiVBAPB+PAHeWq
Cyu0Buo3PcD5dcuSa2t/ptDH8gaSsyTjEitiso3uTtfUEDi5oZ+9moLxRAwORDkGg6y/LUkhRB/F
hXM3KCKoUgqiRN1kepcNEQkBVDlI4Do6UTeB+Ld5hkDY7sOVEyB+cY2L7DxIs0pZ0fxc8ZW8i4Il
991+IwHIhtVISzRRVUcVZSNOR4ZGGjXDrLayRJ+nT/7+oNf2FvuKZcMh8Khejzx5DeHLlAmGswco
S3/gAtuLx0BA9pvA+WDTwf4DoYuc6gfke6CdcOh5DAG6fgqTFQxIMNASawth9CM3iXgTleff4jsp
cZjXwO32x6DOCxdgqC850FRNsJsEzX07gEVxPOHFHXlfrBiq/UwtXvMhvwWxwW08vkuWKQra1vqE
wEVur6XNLyZQ1ETPTqCRhfGx1fCIYQNEbNzSLhJv0bsvAxzD5Y1DHK3qC79ovnLA/hBR2NIcSLuu
0hrkRxPGYmRT+GuOqgCAkcLbtgfBwqgrEQIuf6RA5i5lEngpPkJ56cY4Tqj0Imt4k/1OLL6M/XM/
QhN8yDlLd4eb8ZwJFYrVmFXHDH7WNpzM5tFOas3h91feRI9BeZ+S1UfCokerMKNZrn00xTS4JST5
0XS5c3MQMb3+xDzN0Iz7RJm1UlfAAQccYleB5lHkHaNB2BetI9sMbG9TU6HJUj/SQ99kr5jEM3rm
seRngGv8umpoV5xUJV26mIio7uusOlM0JFAYPtw4shzvXyNI0BC+Buc3qYrZLaamRILpK+XppuGj
K7JkvsxvBO4OTllLLeH/SZzfWUtDa7DyY89q19NKeEZZxvMFTimN76a2+HD15G+H1K7vLZPOMnLZ
Jfboau8lr9a7ogQZyHs5xWQehWjTkCKNarhNmLC/et3WWXuvsdV4cjy4dqyUsSSWKttyBJ1HHf+1
Z9Ow2HyogX2Cm7bwBKfeTbmktwwnxx5j+t8u8XXzA8KYSJNd+iU/V8u97K98II3gVw2oqngbU0Tu
iK5Od62noATiZfZuYghD+HMwS4HsIm+xMpv00C3lBevJsZjH5IlFI0sVmfoBpKdRxpU1uz6FP/LC
+b+sXHfYaEN7wWUhvUp+qjylf8JcKfWw0MGijIXvzE5wo4uCyl+cbJJun88cCW1jskqqhU0d0MJB
yuAMQpSPFBsfbBdhR9fpsarSyCFd6n0vsPjO62ZXvcESa1IJSgv1KdIVQmMCGk4L7AHyS8MyrVU9
OAr2h0A7twlpL1sOK5LhmezLT7zIwXJKU0064QCQ0DfnEGc4KGQZxYshAoootrhUZTr8BW1k1zlG
rMCsWPDqyPIkppLByFOXWVF1xnzR+m5Ie7YifByT38lpucGu1yFbE0lkJJAknKh4ZloHT3ugBEZv
UNRw0q3SLRkyYUZ2iChTbogGMYoMgNcNP5s4k4oT10wIv/r5OEtppC8GxuQZZFO9wU66GnkQ1pVH
pm5jJzIR4JnFRat9EFvVjhRgXX7/vH+a+PBUSKoQ2hvJD9um51PzquRYLupJtI1h12kHynMw0Uuc
F+16+3GPUOVSPx/j/44opmksC6sYZgXAHvls7oyTFXMn5xRVgsG4ZCXmaLaGis0ZXzKb/M/j3L0U
ZYlg9JbMBAvnZ88leXcfWKovIyOqcAKDMBGiZWHPw3vX1iq0u6qgt8HfgKpe4m1gScRHM8+wfD89
CdhuzTknD3vElBYcpiL5IxkgIShecQUqosS6HqravZH52yRcimn2B80u6G87htq6gfYI6XlnelAH
ZJJX+wTPzPzlceDu/50cxHvynF0wYM5haMJEcrPSILWOozzfsNcL9ldLztkMU/E8J2q/wecDrwfe
r9MePxE3tMWzUB6bjY4i9+LJKcNsuLTMHXKNEV4esjote9fjMZ5Tl9yoLWbl/mtyhTB5kWUiSXN3
gnWk3Ur1iAKjtKUIyyjb2h9kvzTE0hF4n7MQG5+CzhweWW810OytEjm8oebzwOn1I5WZ2tuqvWDp
3LJUEEoYnZfeCksczcQgqa6f16HqJssWUoQcO2BrWOJhd8n6HITruHz9ZFOtHwCYd9h4DtFYy9Es
BGfKt34iIQWyl/TnLLKuRm4rz5gdC2wFrGlJ/3adPo4gF1+aV0RMAWMvFmjviBiogaOuwy04zNzx
83V+3zgVM+SBV0RROXnEw21PKbXT5aNLo/2b6i1vxZAIheHQMbyLrGQODV4XMqIrq3jw9xqSJPra
QiYmPKyVopUnWvz419MqWemAX2rHQrOXH3/bEddhrSjO/T1aGkghsVDDoHhCE0Vm5ojMPmkKO6r8
0e0g6f7DrQkNUlUi6LGrEUorNMsmwHkzduWqcXHHfe9qrV6VwdRxkYpgDkf+m3bTqG7Zai8N5L5M
B9pD8odfqYLmUxm24HjCM3UVXNkh68DlxDpKaOA0YLjnbliBiNOLmw5B8u0OTnsNSuvZFPBRxYDn
fD2LFT/ClbrV4D4MOVyaiU+8FJ6EZG+iripRHEqZdIYfg32e9SfkiORRKscVj50Z0HdFntdIRuBG
6misfVz1iAGFQ7cWGjFiSqCB1jWCdb2D4M4bqGBYnG39ODLrYXO6NGsQwP2L8VqnuDPwZ36AIrAN
bglnoZZN4r241p2xFfhnRnNerte/terVXEzhwze1n2EciQ5vJRaifOgzX6k1FmFirKlqLsx62N3M
mlxw+ldTrkMc20fmIFSGTQCWAN510DFD6VHLQVv4D5nQkWe/GJ+7jHINEvnoPRIPzf1e7UdJX39v
BF3C53zdJ9Biq/BawBh+HpGD9pYrz1PmZs4q+f0cBaB0qlyzcXreZql3683kuu2wHB1TS75m6QMw
2We1dseFoasPAxIpav595riZhaPQg/i2LN+wnjJsKKoy0PWG8NfkmmEx0hgiLZ79uLRbV2V2atB5
J9AZhc6NmyoCcqr3CZbV47qKniNGoDH8QJxlFayix92BT9YIu17qd4pBLATa4QxqpY+Yei5njE9Z
eDyTkC5dE8O4mQLUvEv1bQYow4YkS9+RhIbaHn4DCwZ25aDRUrhK0L14uBY0LfxdzVn7QKfopYMc
9qvR4uKv6wQxHg9ubL3IGtOxjnhuJobpLycTpRht7+Yo/XHnSArIDRidHQQsy29zMtlDFjiKyoOd
CZoSt/DSkYj3FzOdW/64fxF7KGfu+nlA3UJsv/jyPlv3JI6kbNGmU0BmhNojOMbFEHOy8xMeO6lq
3+B/ii5SVTod604+6ywSyapuexR+tZILK3tnV5OZ1uG+bw+E2TaL2HaWDl0VH3q/PY+gjxEYkmzT
D2vz52P9rKWRYPmg5WJAWAWvfrfaoInCmcAwHKpNrPVoCPfZ0/YcnRSY60k4fnuqCPUpRy5IgSWr
wmDc1Yr83WrKmu+hBxnAbOYNWyYazlDmccXi/Q9jlt/vfsKdzIUFCU5tD/r55URtpTVMSVhxNiAn
yeepAegwV2Qzhumj75lDgxs2KOWA8tP3BNX/Wb0v02JZXQREH+nEH03yF5LsvnC5CNuU90WL5ZqQ
BRgjF5SgXlcUTEJYIfGq7KWRhaLZ7aAADkZvywa0hAk2Pp+kg39DBesqcTB+LYwNGkBTkn9kF7+A
kzENbhB2SSWQEFoBXPzunHqFsVC6xUAUArqtrmitF1we6mehqb2AJcdBJUnYSwhNzIZFvQHzPklq
a8twWWgdCtzXf9O0tm6fuQUFdWLUcgo71ACofb2NQPNXwLbPVqZRnrdQsDEJttFZSeIcjSgfdApo
JCt8dxUW45dnGo5x2I7nZwwsVG308zxF99ax+DSIC3tlojI8NghLt67LfjvRam5ZrGbX0CEPnVPX
UudPOshArRtmZeac38O65H0AupOZ4tRvZUMLAwQ2Jg2VcnJKY4Hx4Yy83dlHoVNnjdKYhcs91Qmk
pptXZi1kjbNqZ9FDtO31oQdhVeHUFuE8psq0M+ryG7xI+CRZfA2QbXTdQzHZb2gW1xJGlvZSzR34
MX+XKyVti1S6FdGCHB6ZmJgPmpxWFzKJqnHPUHITJ6RkMooSVyTHD3L9HaD6Pru3gS3w5FP4hhfv
5V5cc5vR/F1n3rjJZMogRoYSHarld8s+u0jswb7qar8aPLQkRGxpUyA5A9ehwVythMHuLAJkgZM8
4nasVKuLwK5KxLdwrY40mDq0L03jqKdY35V/s8GY/3E8QQQRsW6r57BS+aq96DOsKNr51qLBvK+H
OplzFxjdr4Cq8NRgtoYq0cBU884/G9KaLzwv/ldM+l+DNUVtKhgm+fCejk2re6YNqeWEputc97P5
9mwSVQ/2unAhkTlSC0egvr/2E7RDINYQq09CLwTBX8+8v20fXLCfuLFSH2RoU28V3Mua7KBxyfJc
U1LTfpk4h0YwSajCSZvHkKrZHoFqyYxP0cY2dnZYHGHIj8hArD691OKyuheUiI8R49O1CbXyn6a5
BrU+lgYVDiRcudeVFxOmV2lVcx3j9NJAkqrBFWNhuzEc5OqSYdNBzyisnQjY4xdiZsbi6X4yrdxE
XR3EM9KMrcn8bPwEhO/h/zKdJ4HBDoDPU36IAfe3erVvpEesrkUCUc8SaoUTq4X2FaBIzmnSFCzF
urUHsUyRWnp/retmQCIuIxhVwue4LipUYOXPpzX3ticpxoW1ME/H9JTZDD5qUcBXvoCYDjmTu8si
PY0Yt4NYRYIzyoAFHa4T/LtLMKI0MgEGfuWOsjP8bHBddThq8Yr32W761BbQGHW9lu9pVa9mUHnj
nZm2kuwgHF2K4QVgvKL8919UGXlH6VoZRDHFS8k5TZCi5mVqRYEKjiGVG0a8zYjms+10M4YzQyPa
l3UkhuKsMI4LchDQf0Ar2WEPas0a5tb0eiAkfj3I2J56tlUDsc/GnfdmsyNvj7Gfc8KRjLO0BL9T
qQqJFfPI8HnbauKX07UyjsQMSLRNa2Vm/v9L1zL2+y6RLGho3nBycoX402G+OIoCK+zwwllwz7Ha
HxPMjGGftrafUlG2BP9LsGXc/ujOKJutnndR7rl/B+B0osroLMBxM21UyhVbHxQS1Z23m3W4HCCO
/JohTbK9Wsj6JGpJse1zojQsmKKC8H8XSiOGt/EGNKKRd20z8YJYjPfCOQ+2tvs1r1f6JUn7qhiA
tI/JoW/56VQRN0ljn/y6M8a0Y9X8fr+3XEeQavbJnTHrA9qRX9V6mRa7TAUEo5Lu8zInfUJVZOq1
UjAf0+B+iyKuAc7OWkYNb4fEQU1SB1u6oC7eDx3BjKq5ywc0cy/BDcHwd6+FoGoO8O9XM42n5UTV
9W07RY3WkqPONhsQz9Z0hKhp7Cvkgeohwo4DugEDTBZNllV1CrezDXc9r+ovlhUd1/ielp4NHp6c
+0wwvqb6iqvaVQ2Yv0obCkTIMErR9xOqtfUj8dtOSLC68ZSF1vqewdRvYQOC3TsplNuTWg2Ngy3s
br+VA1sSnG+43IRuHHqle4/OBwyDPzJ3fV/Ha7ibo19Ji/17+2cjaHnvW+xsVvFVQKM+O4gFMgDk
OlBVIITIGhcuv9APvqYDZCY6onyApmM/f3H0if+OrEd70unlXtiEvM/IegYJXWZ1ruBn+GJVKF4K
nofB0wWwg0XuAyqHh7wjca2SpJwZXgF8PXk2+l5cwqDEoAdgPOl/GxLNkMRCgYw0A4SSjOeJjQYD
MCt5wbwLH3zhiaZ13JtE8m3LxBVEwSywl3OMnwhypr2jw5eO4bByQ35Q+tjfhP1c4fSMr5sN/d0E
UGpxP5dMlIBu9zBb6TtGpVD/WcBPzX4aTbahuHfUePgZgvict4LJEzNFuwPsxzp1KvJCicC+Slon
SxJx3vpX5q7i1+cLO9MK3xhdiJDoAr6YZF43VGiwahnJfJInMSjArGrYpj3cKHnj+dvXgwiKMNTU
LLuwKuYqfYD2fHbofacO+qVWQsGUX0x/FvuAA2QREe/0i85ixoDeuDJGLC+VhoGaYEFrB6X2nVhv
KqoaSxt4yxt7GX8H9MfPQ5ngCJzLq9CGD1E2Z91OYfGPzNeAZMtDnASZu/2wokmaJNeFhGX2YUlB
gGbVOunr+TwLetECNftByw4hjubRyfsj2MSt/raRGWV+jDiDSKZgz2zvrID0ySARraAKGgB8hNnx
VRPaxFj52UiX37HPeuU9/kEjmeiEj4Jc0E/kt1LQMEPv9Y48MZuPaSjk0LY34Ub+3fvMQ6XfuN3l
wTwzYBXmDilSKfh6oGOmuH0iXVx8ZLIKT6hFhfN0ujxRA5T3rswNM1EVXuPt4HwEe61d3QPeaUku
/FbZptPlEpKJiDETH4RKfpOVrbR/+9vADPtyrdTHR/3ewx3v14eKFavbOXAm14t4CW1E1hG5ictc
+zpCHn5py1lM86MTF36gCG/RTgp5JMlOVABt5Djr2W/B6oZcb1W83NfKqLk1XB/jbd1P2RsmjVRY
vYhU35/b+gwbjdqe2rMIpff7xMTOhQiUYg7Yd7HEunfUg1Qa3OM9udQc2qIQRqMrCnnE/rsC66d/
54C0XI0NCxS6D3HsL+NLgcHYTCEGi8Nq9WgT1IQ7BZKFZ/08T6/5DonqnLEKpHwwlIx+i40vKXDy
xShQVx6BLMq63+oV/Ys1PBQYJC6fdaRkjOsq+HW7w/6VwLrzMIqrgANnLxhUiKUHdJOYaHcTNxPy
MLz7+pKFqK2fLNXSaD7CeGz3ibGnCaOwNqKxegbNsU6YgH78PdZcmHQRtNTlsqgOTueFgnEouJMr
sVMB275unN6P3AxNC3TJ/3uGVXD/tz2h/iAdIcFChZQYTC6mUHOcYUVLBEgCKsCB+QDJCBKi6sX1
j0n6t+w3ODRuQ9l/l6Qgm+BTiCzX61K1r3SXmTwG30j3iXWVM+7L1GjCIgIsdj2xyTp0UEHFmY32
udtACrA7jAwx2aNeMgBw/eXXqJ82qdkMQSEfu8ccTOfcmobwg6lQhzY6rLI5x84dcEJCibqf7FWn
m6TPUBwdvpVsCUZn9Q8pmYMm0Z29n9Z9S3nKbhokL5KoRtsr8qQ7b4uGY3nb72Kpy8DBWMdEPsNT
EYEAb9CX4FzvRO96wLScVC0UT9KXw/BwC6fpW54S/VahwpaszkNfvrlqn2DxF7kBvxZFNOBUz67Q
FRZSr5ftNLvvTbXPfA0fk91o6UGUU6t96y4hzfF0QjvMmUvrcBZyrTfPRoMY1i1WJtNWfxV3oNGi
7DWUWmRHxSQfkEz+aHUrg5CxjccVRj1ed88y5T3Jk+6cvG+mb5xpwrZT9Gdk9FxpiqCjfvQiYd8T
ktcJMHzAhEcglW+QEacIJ1MMuICfReR6Xq8QrixCuRR8AOli7zs86+XhkiTMHM3u3LQ8k8xSdjuw
7sVQt0CeRMcmvpm9rFjCQAnY90776m2+NQTZs8VTmqyJbghBsygcTI/vEVRk5XK4gSMxJRNnbzYv
YLqIZNrx5fuIuOt078/P20IMDF7CtjyT1ROTlfK9BeHiQQzxP569FsJCcZRuD69xfXAQQ4WpZ2MG
WHrohYXtlS2IGoQJ4TnMF3xeoJn2enjASzZe5J/9PODJaeEx6CYAZGzL2z0Bdck9LXv1aXZBSojq
dOqjqDopWs6Es/bMOxF2ztk2fBXAQqGiQ5zifmqHFMUMUC77WVdQ/7MmC8taQqhC+7IFe3o65Nqn
TfSPJw/JNOsoDr0xpV5hi0GmX5/dkl5Przs8i02QHhtKyoY0hQtZ/Bk+mmBYfS7hUuK/5T3c6YfD
rbL0F7HoI5BEpWA6v15y1Jl+PbNOCew3Awz0+Cuq4FjtwYWuYhYUySEveiCGRafcJc15+IyXKHb5
t0FCJKatSPLm9XZCmEu/MxOffpdGs2q2xx+Uwc1RVZhcBOKPWb0xYPHHauDo333ljQs+qdmkxaA7
cq452puePTWCfme4oDvu0ezMJu19lP+X+u92+RcO6SIqUDwzMWGjV0/DY7aMlPhA1CDZctaHFGKA
v2yu4KY1yrmTBhK75V5LIRmIE10Bub+XoRkp5X+jLOCQpmO0UrlpCJETAku/WejVjdYoUQUAG/JW
K6jo6HzuaprTEWBCo5kSJl/UlXmIzL2hMbb2FKPJJAki+hdOmZwQsNDQq2uB4vBddJY1FwII7v+C
6O3cIXb410wpd6QpZ7Eq03gJu4OoAfdt0kS1LHUHsTaq0fpqIBjfCIuzQNioOCQ9dPKc7FRtDDx/
qcN5G6ipr8n0F3YoXCuhvOqqizktP6ib5bN1jUr+G2/58Xihi5i1BV01YYcf8kKH4VRacu87xEIB
h2eP1UC7I7z5fmCv8sZdbFSb3TKE2h2hXLIlEMlvClmAb5ZPv6FY0YNDorqwRvTqoqW37DCd5LWJ
9Ggoj9M7OdDUbO/gmv2I9f8oNBqmuqhcBBOB5BK3S+kqOb4tEoygu3AeVbxrCqY3oWlAB8QFJ/nY
0grqUVxyxp058Q8MJ7LPgsk3xPSxNnVMJ+FTt/YgZ7hlmVarrZyZ1+z9bOAWASqXsdWuX9kNgitR
CMJ7XtI0UihUEu5z3YcwSQQZr7rAWZSbrchBYK04t/eZAKqsw/I5Qnr+mPtMTmtR4SFSebo2gTvD
JpxYHLfu53qzlf4GmkM9vSxzC225pJUFX++GDXAmhbcGug596cy7D+huZGu5JbNTujDHwc+JUIXv
uCOpCXW/Euzcv5DjsGqDx/BwsOrZczaVCyuzvu/U+3L/uekxEBx9y5KX8WkYgV1nQU7YGjPDjcdj
iBiiGhheGgEtIaus38GGLskC7XyoCqXSDb7l35BtjXbSvi5xkOMYGgQUxsHoHdV+29C1/nxVA/45
srJPuWEtWuaG4hHVNTl0FlJTBIVLOt+nYZ6JPJ7NHknMsiqFiVWT9LjFFZQQHME1cw5Kd+zoALwo
jnk2/pcPuWu+MgsdEZhdP3Tdmdid1C3J8/84fB8YEccEkLY5v9HHwa23Yz+Ntns+u64Na7bwcXxE
f/obhy0yCjqU9zD8HDqJxkOI+HeT16SFHyTz3Nkz6CWp4Wm52PJy4r5Z32g2ywX4Dqg9a1FEAhZU
hyefubmZrS1N167+VjLCn06cJOho77L7krIULAfSNwlYhTSeUv9kPZFqLPlv6eV2LGN+Wvi2K/d9
nGc3sLwe9jtMvN7j1giQh9SCFqXgIK8WWhd4w7GECJKDef9q2tdDZ8SYoMDIHKyQGm844tiwT3oY
jTUNlEOmld0s+N1i+AeHMV45lHMVn2oYx2b5tbwr9ltbh6nyvPWCXpXm59ZB7b9cyLyKJgggf0a1
VLRVQo/lMjFdf0rgTXOPQO2urLf1Qz3oUh5XKCT6m/ZnMK8UELUHOcIj79K/GnWbsoKWWUimGMIA
adTlxBt6pGk45ailf2LY5/dokUOy8VsCiksz9PkRpCEAVKWhkEO/8xafv26PQhu4KaxC0HdkVT7I
ufnNe/vXOUT8Hce0mNd1POkE3gAJhPTU/CCsy4RgWSkbnVjRHCIK23wbsmommzl5FoG4iCykGuN6
654VltT8W/NshjNEKlaQOAxHCAIOKdijkbP3wauvafT28RgSMvkx5ep5m0TME8OvL35f5bE4DdxW
OAe6MBBjWUxBahJHO3eZ0l1zX82mEHoStyk/1R4WKvZmTQlTRcsEi9kKSX5VjGLHQuZef9aQLeT3
YEfE4pTt/81mRMejA2v2HJr+7ShuFjW+RJYmHLFJc3HajNPeYCwrxsQeFXwTXTE9+8s11V79Nl0H
ZmnUYea/+adX37lAuZIFqJMmSsPT7v7W9A40dc/2QRFj0sR0oCffzP9RDOVoQqDiCXCzgD8/XOg+
nzYZ7mlDyaQW4T63Kn3bL40ZWIcXoUC516VFrsGzqBlDvBt6LjwmgnnK23BsEMjDjUJnuZZKj56r
jUa7Z2sE5sIAYq3lJXf2SnUNrCAC2EFwblTF1OwzbHHfoHRWeBoYbZZ6IkFjG9rq6U9N/4mufDE5
O1SI/9bk8uJRaJnW1J0/dC4jyrWC+z3piBL759rDmwA+nU6kMGMUqDZ93dahy2X7udIpTVNggZgm
92JBlqx+5JEQwVJDt4ohntoNRKVM4GLM2Uztk4LsKZTGJvrlhmJowDBzCI004wWMLpD2RFl05tx0
eeabwx79tLPiJzP4kBWzttJWPfpgSfsEBOv4eAzF9RTecsdlwxZxZJoFPJCpK7+lNb1Ctkh6F/gK
9fgJM/fjwg4Wb3XSwEH2oRbm1bFjmkadje/pF3PxeIyARAOSXGGhp20AWSPMXr/C9z4uP47GQYte
kf9Qm66gxMaDntzfsObPJFVuBWYWIQoMVxbpaioTflNEGHzu0WNb0rWhOaLzlheQ45C4fkyQPsXR
Nn6jeqMJGqjTahvpCngRYWGkqmAa0iiDs3ES2Aic60mnT3RE10qJ1TwcfPXZheV3u2UV8EvB+ju7
hljz6c5hdYizvnLSiYKxcW1nfKDgD3w3Ne8BDEweGHp6APSXcd0X9cEsvxd2hK19/dnFs1bCRtP9
aKAFtxHqljXkxXssHSwjaqNfFQK+RYDh5D8k61TlyIBYIzKalJBvadvkv0cyNu5qWnph9c7NZU9r
E4pVHk3uwbkyBuiU3wxAsOJw/Ey9E+XMzl6YJ1sLzUKpDnz2zERvKjuhO69h1EuTkioKTBqO8aMQ
bHJXELivurerxvb8baQq63tpx8OkJxluIMsVk3FDt51iKhbjayNkl5DlBHxs3ddtOX6fK+h6vyga
UO2f2VW+5oJnkh8uCuS+MZpEUhlsuwDob7vukzs7wCH4WSdFC4o+xHH6R7SD4yLWYKW+7ZilhBKw
pCARAdFG5U55yizzGmQ3TR90xmohUH5TwqvqvZfnxSKtngtVBBS72lBlDFY9ttz7/JEIextaZOVl
6Rn4XI4jo+JgRExod2PWzJbkKs8S50UCs1Mw+VOtVTFLju2naezB3vySxSdU9FpuVraUbsW7FmFW
iIY/d8U6BtOJcXh/X2J9KCzqPikTFi6qBdFPPs1Zicp3j9H1m6yjuKRqoHLVnrf/fyIFMFeuk2tQ
fpcHXLThZ7Oa08yO17beFz1P/fl99ZdcoohN8fOs5zFawFOjRGt24Bx70TB3AlF6ZOTUlbmVfD/o
1HAjPAfh1FmyrkDU78+nyYVVM3G6COUwhDhui4AXtTJj0z1swrES2hhu4D3zln5oKmxQqpN8lQxv
xKBvkBhpLboFjdBWP4VHIh1zP5j2Ay4sgUYgjiXidSQNRoGeD/NwVzCDhcl4iDoFX4ceHG1dWG0U
9wD5E3ZT0KEtUuHpWY70I9Noq0a4Aa2wn4me2WGp23TwvqIdcBYpkeZYqIi7aFBvqlh+9iuUAqjS
eesXI3+mD0vur/ipIC58NPe0GPcAmnWyU8LugsBjEvRQx7ZBLzHK31pCUUX/3wQ4BEFiw2Kp3iZk
NaNCUVmxEnCJXAnFQDrrRtANBkHicCkgF50xDtetchQ/7oLi180asNyS0w/P8HcA+wjTFvIE5GDA
7azn5JNm1Z4oHHHtRTkmDbioa1Idb/C93h8hQ3IHgVVv884WvMQxFOhhlrZXcvfnIB+RpZJOcOvW
pAYgh+VpK5mWS2KbxGamxOA77ZdPmPq0JzbWHP77YKNuD1eh1grKygsIFYC6nWEek2CkfjXar2DL
eCcKuF/62+gj5nFwDW2vmkOOxwekSEoW8IdvB15RwRwxw4biCZOxzkvT/JeoIqA8ZoWdQRCS/HaQ
+uIuzySIdShXbV3sNBbOuYxDTm6Z6ZrWREDRFlwmhwjB0237mOtJsVUidW9dw3pHxFnJpX+3SDNF
VFYSZ0cLNqg8J4sL6I4a8RJN8cxokH0eL8SdYnLPkXBXbYdTWe2mnsLZWMLScgegYCZhLaDBJ7nO
zPLmH+6+E6ti25YIiDMCAI3K2RZOUlowNiK4329819vuHM4aAYBdiCSr7n3O+RTeQKVHwmjHpOP1
oMRrv+0j6nzEULnT7MgdyvT8o2sN8cfKbR4Ik5NuIrDT24ihOmXr3Fn/6BBU2FaGjxONM5cQes/S
G2sFmGOeFBYi0w2VKL/f8aClHZUYm/MOC1J87ebJQUEAeO5jpUhU436ROubQ0rIQFMukVDc3zbTr
Zi6xLNwKvkYKS0kfY/7MKaBtH0zmihvDsyBrUzhuSWOukXLPMeII0a8drybOVENyfmJjouriFIT/
O6PrpR88mFv3rut/euUHAf3TyFjchZwELD1u1mR7Yw6JHBemHzGkP/MqowjdQ9nGAVgMCOy/6AJT
rf6Yr+SJmyJaLXucNujqLYgF4O8iREZxei49CKv54NrSI3Sag1RKVFa/voDn49BPNnG0XjkKMdJd
MTQBWFfINoHmStksrQ6OgBK0c99ny7XgXe1TuLCZMV5b8PKJ0Dh3NQpGXBqT2euwIo5mbxtK/vs3
EBPVx6qow/PDMOVB+U/7WIeS4edkc0avkGEVzfiVZdtsuk8C0nR1NreP0SAzBTS7vHd+IoUdYwnk
lr7hZUuluMJTYZfStCWgQezH0ozAddYqbQBQ+xS50NdcrJ9ElmeazKmktQQHvfkSUhQd7hJaGKrG
WNyIPXZRttEOuaDCkAt6P6TEGPII1T5Z+TrF+A132H0ifslaxBM7XsRrCHTgcVww0stGVIgyPUx9
bcpCiAfo+Jp/d8zxNIALpbHgHZBEJFTXjBhgWCcBg13tqf2MZ6fzD50+HWBJIhI5O5vfk8XaxooW
VEKDusNshYJwajWPvITAygDaFHqcRX5KUwUowwUpINZ+bxB6+KoiamZ/UFn7fFo2clrftb1ubB3+
fFWZRs3gzQNYs9uXpDPZuqiAYSF2bKwVVLkDmazzjo92LRvPV+Nm9dUaWNeXRV9IjQu3R1afxuA3
CDDvBrFWfvd2HHzJuhY6WiROu8juxEXI8eRFu9hOMhRjpT3Bw3xPj0RS4YvG0eP/6g7pgzzz78w8
hKZOdprhcaIt9/CV0/w1LCm8hZnFbm2biuKTQ8ggRxDcvx02w1rZl/AyJgoOfWzWd5gG/n2kfcYh
lgAHAVSmWS083MnCBweph+in9/0qr5WnV242k6LFP10xHgoJ/U1XK+pX7tH87Yz/bm1Hywhof2fS
gruYIhsUJofAhO6AFZQF74SPt32TXQ02zBZAfUNSbRCnrdrdp8acKkLI+I7cMMlEZFjpIjvblo6a
jwzViSFw22KEmX6yurTXBCLXxhuQUe+K/9n8aWl/t5lYShps3Yj7y+I3Iq3JPCyD/aZb0VY7EHbD
/intjWUktVK6JKycYJZeVYwyxJQ7fh11wqZsGnHoVtDSd3e9qN/XGwRuy9bcutJPdSjvielbQsDQ
lpBpnONq8AEoD4v/wcOojRLfp49W1+VZtuuwkCQUXd0ZZ32FO7Kgk2D3g5yEXWucqj2OpRG96omL
yc2IKdeK3d3+oc46wit9Nc+ONqvLqo/gJUNMAcWn3SjJzVl9fBWMaryLjPp/bQvO7PaQFByiiSKh
zd3SW4FRtRg6lFzwg8hhrTC/zt+7S6Ow56SGeGD1VAwCo1xDiDdN+Tka5dtEYZmzC2D8M697/TIF
xIP1yH6DYzANdef2XR44AHlYceD12ZKS3xUkJB6mvkDvij1CvGI2AqLf4DSID+vR7Xnz5y+qzOjP
IhSxLiZ7iyMT6yLwFk8s2hSvH0iprC15SrlvyyI39Nms55iPPOXPK/2k4gCRAv3l/XFtCDpP8BQc
tu78HpYx1ty0ISkw6fGIfWvRvYMx2Wv4C80cHBO8+Og0knRCA9GPdEwQMi6LQkV8pjLzbZM0EceE
Km46fCNasS6NFQmQITJhhlMZ1HQHLff63Sa/LLv23PjzplhffnXpI7nkLjOsyN3bZdYNc2o8t4Sa
31fBS/NDnwhN6Q3Q84L4EoT2kOhqBxJEeVQ0vMvU/1xp8/b/8Fx2xnSDB1gPJ9KlndNo7AAr+7od
hZjna2/DcCyxk1lcPHmol/Hzki6v5A5LrhN0tdfvn5ONiM+ck3pTPPrco63ElNae/JViZ4uSqFAu
NakxJoxDadULL0yYTUlF93QUusglUqDLRy6WUraQGn7pzKYo7YdpK3Popfzj3hPUbjrOgoOy/O9Q
8DhDyD69wTuhUhUdfiUutiVQEQT13aXQqxc8+SfQWGhUC+VEP9/Yv8XcjWjl4ixexUiD91DQBR8W
FJSNc3hQ66mk1dI71TTgD1mortg14XID6mKCLMNdAacDuEt1Psjt2SIIkkgqXgkj8m8Q6D/OYb21
6VUS0OFt892kIpzE0AEXsjZ/FaOvr74/jEaaY252z8DHqsHPA3Wy/Vu9QdrkrYEUv11FlSUM2PGO
QUtbUKGoQfY4dKI4d+YO93yqyrBFdgvaFgVQ45N1u3HbliLZzabGqdsXVmermh7WcMV48jcc/mwa
jxXlim+mgEV+DpJT7olSXtSk0cylextGfoTUQhmOSvQwaXUyqgopvcuVBScsM3yxRMLsAVpUTavd
CAXwPIqURymvA968N/SSKO5Yx1/FZgO/Y8NxLmoUdDNJEIiDAfIFY9pf5sqZpJrLSy6IUIO1qpVZ
1maut8RIdQQwTaTqTFcPXs5SxwwWcEouESWEoWSY+i9RUwoRupBCTbYQvfSb9yj+sshz9FnT+nxd
uEtHooCN5jbOojPXXTRsVe3a31xIUcHi1MSNbIYXRRnEkfV2Jqso9zUq1G4ITpCMi+vIMTj00F06
4BooW2kd5b49aQhXnavvzJwcEBn3LxRs+eMt+guUaEO3Gxd2+V0DhRKBbYNaJx7lIQwu1vMkHF5z
ZTJpSLBAr0TfsJxV8H53xjSJyvdbLTsHXeCRCo9cGLOoGFJeA2+X6zNmN82RC78/aBl8HxCXO8sJ
9Jg3vyf4WPHhPvOi+6hxBwwW+sBXZjc022HSdcr0e+k+gnBOVgRQNkMufFQLiB7ZyhG4N1QIQR0G
4I17O99TxahR2Z5QkQYnArR4ZQFEkpD487zLwHRBfNwv32ZUV1Ff87SuiwGaqdfQA4N6IJP/iVqJ
SfKNPz0prSJWLCg2N3uIujxBl4yBG8DMdSeqYT1SA5TcQ6+YaWRNTohYkCONnoS3PzxvkGLGvHpA
a5cBb3oWuSZP24iTwkUgzw5Xf4VDcYE145vjAv6Hn7BUEmU7HE9j8HuWZ4qRM2E281s/aZ2uXfgF
Xa5rESKQlMuE2S/LfsKj1UPcdWkzktPBfIJGnT/uq3JsW/8V4tZgtnphcbOpoDfIwsXebvS/zPsL
fNUM5ZgHHcEli+KjtilhjYb/uUTnFIB8tYT/sqsTaA6qMx+EwotxNP3bUcq5jsoGy0rFDhHeoIKW
24PhNVbKYxPazpYVogibXfIdHKL/I23ODzKMiQhlc17fKw+eOIiexz32LhOWtBaAU10UIxP1nL2e
qewR7dlQbN3Yr0PsgtpNWnAuypKNqHNBGSic09f/ZZ6/K52krs4ukdfkxLGANQbGRtlVOK3lD+ri
2/vMWuWX9DlftB6YJwwgzutNsPDvT7IIokI5HLV6n0hEfIe9CJd3piZvn8WhoX+UHMz2SKw7+fxV
wyejABd/eTsrTHMdru3yMEV/p75OcaPrzueNjOeYV8xf9I3pdEVFppQWPZPZJX9oZuPTQRmdTFPT
tWFET4UwkxX+0IARthBg2MPJFv06GTwjPLt9KA8hJUPZUrYcu8iB+R2tqlPVmi2VLrXZdwlmUb1G
U3kzNm4TuhZntdg3i/yoJImfd70tFVRLkHqh2z3MG3a1W62RdhW6q4goRAFfZdt02QiHWYgZX/NX
az2O3gc22ebXJS6pp4RE/I7ELnzESQCpRvU3p2J6IyYBHSfEbEUg3iE9YwTMDqMu6arEIhRPlcYP
l1dArnJWtuhW3fHVUp5Ra2ftzawfzIq1RCMSrOsMQBxGClel36MBjN8hXCEaNtxJ/UAoMR6+JVxq
dCO+a5tilQpWP5bwzOfRiu3vsDkO6xRsRWIYGI62cWjsZMczIQ2BDKGZ56Fu8D28Tl+pPRncruWh
eLjIYVqT7p00iV5XUznbxuaFSVRzKofDgmuWQCy89jfZYqoWh57rbOssbJ0SAi8QFQ+FEe+3GOTf
UqLNiGUhlapwCpZejNtPzTSaPsTupojyT9TZr7K1H5CiR2fjmtl0KUP3nnNyxQFGp3mV/WtfWsHj
yWw5h2y9pTvOM493gDNpL4TiebFmrax6DLMW792xo5HumLRyuO7lslE1qlGlTdSJRqkHWndZnfZ3
IH/s/qCGDf6FR8sIv3lol5X8vQj6VI4Kfe8KYbLxoKlMRKfWjTwworNneqYwORXAJxRIJS1WiJUA
Zk0TZ0JHmDiaK/M/Jeh2inuvIFImAAm0NYkTMVzIXCGtvQtORi9xb110bdMRlhGV3lCLNfQ3EWgH
eyn9TrsAF9llU6JXAlAtXh4rC//DMxCuDS5TFHjCqs8AUJgoNFgDrFazsH+fsuZpTV0tlucyX04n
CQ0sylsWNincusAsdSJanotRX5KlmOhq6KVV0fKkbOWAfBUDcMPCFH3UCEz3lh2L/67fU3wkIE1Y
9tH4vKrwokRkN8GbTLdnWd0FyfEgW59P3Msh+mWAk8gYkFC5apTCYMoMixK+P2hqvhHDT8T1ZmmR
cNOtpodnjPWtCNimjzM6JMWr3TKXFfQX8v07dHbtStpCnONKHIfIHf6GWgAuuaLA0pOt2ZQ2f9L7
payIQ7Q12/F8kJGmOylR7GYqO27V2GRVa6KuOmG1dxHbPv+BTaoMZaREmr+BpofmK3/GKwIGY/md
Ed8vtLw9TmCpN6T6OuS2cptmdwkYL6qpIzHVUbHw42ne5p46P74uQhL6sOoSD7pGJFx43SKgtPX/
hEvXA6p2fui32A9SdXUzdcVQ2KH+NT5Jy0TyGYh26wB1Mui4SfPjZaFXXu7H9gEQO948PywIJcjl
cJjEdvHryFKA6PqBIYQUV39uIQYL715d3dRr60nC9NNlrCqBQgzzOhJHE/ApVbrtJv46pPjaKjt3
XHxSBQcZQ2FLG8GCpkbSkXZizmV519jBwywtfZcrIhtbj3CcE4KO1wE+A9pxzV3n0vCdW/2mdHW2
ZIdZ7Vo+/ioIJzx3bM8Rz4/g5ER7ux/F4KGomePs4lWd/4H2OU1sBrqhb6hLMF2Ljq5Fcxc6Wdhx
dqKYboBk+MK64bN5ZjE5YfUgzjYU6Dnh3fXvM3Vyw3IxV0mOp49nN8CecfPDqmqc4epUtV9XKH7Q
093k05TKw3gtVcNmAqtzbvaCb+ROr9bFmvA8ZXb3IdEZ8z3eBMf+5oo566ax2YQAmtKjsVP2Da1K
EcdhyJQouYdKUgMrQNhRfG1zGJc+wHe4PLby/oSyCF04zJksP+u4ETK3bBCyjdGU4wPKoN6c7uiu
nPR2UGWTQg+zP61d+e/Z8OuFXDb0rcNhiCzutlN/FtlC+taWslghFD6gN1AmAhk5Y7iMt0ANNT2J
twtWEptDK98VUXmj4FEQsm6ejeJi6+XvneofIDf2T9hG6cjHju8ukRB9c7lA2alkNUa/fK8+SZNA
90qdXH48d0WwM9fZe7e3Q88MsrSrtB13mzJntL6WPaVDCOUHzxIYi9R5Pm/aI96QrsHbaTSVx5NV
FbF8vEtsFDf6YvJJLD/fReF7ZSXfXtgCU6fKNSfyBGq9lDuvvCiqT/boWS8/yTBLyNDcIff3jhQB
gzYLD0HJ9DfyifYKka3iu+Bje+slyWX04LiNadfi4xf9rGT3e8RieV2vi+bd89FoazqOlwA9wxl5
CYDwTMOiV6meLHSVq4W6mqBqZ44DWAEm6uL+IXe/5ZtS6vGzlsg0wG4Qgs9RVSZSibYgV4TKRzym
v0OupjI8Z19Wk3L1IA8cL1gd23n7FwNZJt/t2b0LBpn1anWDB7wHM3RJfizS9xmtwbo1K3X+38/s
wRW9pHbEAji1XktX81Qs28kB1bPT0jQf+tReNwZrgzfNZtK+os10cFj3Go8nmlpCmw5dafvhsC5s
09n2UmeZVbRqWaK1RIQxvd6HtNcOng5OJNm9h5o1mIAAuWvFSwuaHA2sa8aw5/Qilhud2a5v6Clg
nMd5nweB7vsgOFSZ5UQxG9Cl16NHnNCM37K7Qlk4bhVyjTD/jVliP7Arwfab6yEkgEh1I2d89phR
Mip6X4f6fbRrL1dQml3Ojh4rjEn8ltFakJVH4TPHvnzIML2SfNgdk/uo/CJb4UVckyMzXGAXGCrv
hR6XjTu51uTIBHbLYtfPRLlgbvXduI1aGtIreUoKH8aHz5CS0SI2KS7JCebvBPtJZbokrqV5AgnZ
lcF5mIpTqRZPsyHoznKYsOZ4AjgmLeuhEBUn7mKoupBwFwH1VchaCbFRqVdOrCh0o582daPgKKRu
wxOQigCB80I5dMtEFuVXXywZf4QIvaXz8krP+QeIOYbzgD5HjizyTlDSeYDjZAYsWAkUJRT7uEPc
d5be9P1BErPsQF3oGL4s5ReigCZjuRGatFKw3QGb+6awbuzfEfjlFn+KAT+pj8cpAkUIhU/EuhUx
c/j1gtTVs2NsmDpWotGr6hLtOgvXTnRTQOn6R4WpENCL09j0f17uDKiOgN8A+gPiisnAsE0vSitj
bOUGGHwCvLcnOPAvn4Z4KV/f7hkldfBlDsP4bOfZHIppgY6CADGKmYS1OKxWfwEFjZc0fj378t39
7AVppr7P/29PV76m2ah416swy/7auprNOfu88Bx/O4vcNQFbBQHPEdCgIpBxzKNssZvsy8iu+EPP
KeO9emmBLOXXfMh5eDzy1kYDoCtGHvHO1g7N71FkG7/pnGJqKFZq/h3y3l06yH8WCFrHx3RIgaRS
4St/r6t5Aa9J2eNYo2kqlMiQgBTX4zrRNMy8v9ZpmlOr/WutsAePdVAV5ebw7nTn/Dpns12juNx2
DNYr88xVXWvY3LjbCfPLJUpl5O0y6dj2Zz3+FxGxTmp8F5oM4wy3WMJIFVb5fvHR8g534rtCgziS
IB0UkFKsLK9RaBayfkHHX5KZ9P3Pwm6dvFo5vYrkoKGmS6HzhG8rYbm0PpDc/NH8AkfiCC+5swKP
QcmQdn9dctJa8KRVJfIUpdOP1Ha5UeFyrD186LBN3mA674zfP6skrs9lMXbeEQnXzLrNLQhGjkEf
fScPzvU/6bXXOY3QCHnYwHj0UMImxe3Xse6dGCILImk+XHo6bYQ+JMNKdXdueIXkq8wyahzcXSO2
uLCT44vLQo4CjUjTL88gOmfdTtEuboP3FDPXc+18vhso1CqUHWCI7i78N5PngCIb5cxv+eOK3GBy
T1aYCBVLuYo2TElU/97ZVCMDyMJu7EOmYD+UzUw6Qas6+fUR3aWGSiifAgwXxNK0qHPVCFTFgcc9
3zQU1fpC4SPKkWhMTYB4lF7lj8FsUClbXwDTTiVgD8AD1YOMLtEZD34MKEpAqVd7RDqpdkSx6dU5
fOhMI8FnAYyFCfbi4j0rYM+zvnh8uu+w+b+UtHJlnwAx4g4ad8UPvJXxmvYGybXlsbGdSMQKPiUU
iDACBEiFU7skSZV0dRCLGOJnYH5l6AvvSANKW4DZro95R4bK0N/oZ3NyG1RWg0WIs9jcBo7+ijIe
Oz+RHNsuk+6FvrxTsGMBBQdLDNu7Oa3DFLvUnkn+P6EAI57u4FvUDbkxxR53I9cOt3kSRVnVICdZ
PLBwItdwA4l4LHvAyki27EQMswwI/MoRJ6/PhTNICzn1n5Q0trEwN37rtgjKxbE61WK36e5HYXLK
GwEIyH7HZxF36l9GCr9V5JOV1ms7gcnP5j5FNBkkw1Ua3bgi6Lc2e8PQmisBX0+kz+WQhzqc2AnI
3vXaya2h9bMjSs5LjF5xVqjvz37fHOMEZPpsI1jW5JsIFqbhR3VnyPj90OWeTV0vZ6cW04Sqx+p+
4L3CEHbUJ8O9ct1rKvaB1QMig8wCBS3aQ04yaB3SsxhkKVRT2LHDKIcL7WD9oO1nim3pqUZEbTRv
1RlZ9+M1YMuM6XANics0LyNUG7jRhlgfMYRYS2cmbajzC/QK9OTgFyratUr/vAMjCQPcjU4hujBE
sAglEc5e2bZeOhrLrYEbnaRaFBHCuO1TAir4Lxil6ZBcIX0OeKHI1P/p8R87rcKzrxYL7Vw1v293
9DsZKbIJK0Kl/I6KaJxBiSX6I+/l8vuOv7abfgRDT03Lsifjsft6REc2j2ulmXps6rKcAPuAff4B
dpaIIigS49P2zmQ0dNEsEenZ+C59rDeXGe5dQmS7C+4UQqTrhi7MZeRdAjFhUokN8GZ9N/t3yL/m
0SZUiH4vZRS0HwGXzQEdGa151FqFk7+/+Z6tXBMDaBpJoP9KUvRxdideXosyiMUg6fUNLXtxy6Hn
dv9BLUmFYuPlDnBENrFp1xuUAH4BBxdtFY/SGa4Z1I81QVi+NKJpeAiJX3FVwf96DUu+WEItUF8w
HI6nToQLe7MXwz48REy7OHnqV2GWZIfueWoKNhvTZ3OV03FOTGH+JmzMIh+XQDovXJ9Qh3bdwQ/W
kCIvZiH+4m5f+j7oyTXQ/WDkL+CyGPad5OFX1Qe17spc2agakSPTavXYHtyIiU/op5UoV02e5eRj
9fGfaHAjk3nDff2qIzcCrcJT+XLKkpa0X49mLcJbP/mGnkgYoBKZ9uULlVD0pR7dgINXDfB3lPuH
AJ+i3sKe78yf7HZHfbHI7CFTjG+VvI4EbsofiZrecjh/MzOiQacjESSTcY3LGBR5IYXKB/xDkebY
0GMofbYQ6oS75JPNo0DQSUpwz4gIV+VGW8xNkPyO7WkrO36oOcbxyFQs9Dg8nCTx+XAkxXkKJpkN
kYj4X04tLB9GC+iA7qVGRphJ5a8xAELJgmGRgY4F5jmtzSiJ2iwY+rMyYONMtIbXTBZen43ih/Bu
p0jzrdI6L9Z30mX7m97aB2g6K+SrTwhriU7GTmfzGmP9hiip5cspomndWPdUfMS530q+7BbSVqiF
QHPU4EGAoSoq4whL7V+VfnAOdrj/T/UoD8e+cM3V4QN0lFrKqGY/+Ftr1syBZcU3hOm4v8iTExy1
H3N/ucMmnD9nouR13iPHkjfA+NXZJGQd5OQZyxkU8F1GBVHZyd03El+P6WvXli6c+8c+d7148nHN
R2s31YpT77dUPt9DJUym7pf2eKDAmm1dGb1LXGQR2geI299su4CPIeBoToOZCBfIR2yBl4AD4w8Y
RUq6o1CDLBbr1ebvsMprS2H/uRC/wQ8AESrVdMEjb/Y5oBxJKwiYFjXuZJEvOyWSKwQ92kUPf/1/
zIPuk3mBDs8mdIF5Y1G5TQZBSUM1Kjm6BRDzqedG38nvozCxEIN/sdaUwNGVDLj/HY0hu2pYKZF8
OOHlayjqS9y30W4WBGUbpBKiiyzMlRa48UB8ZERenqQlDqQN8m5nWku3B6qkSWsuVrrj4ZKMJtJR
iehB0ufSae2w61+EY06ta7aAoq+iGap5tgy+t0r468kKGqmc5Rkx7lgn1HaZ46MXMQcbRkUjowOi
fLPObFV261WvtkEsE7Ro/BOcvjwmiOZoswOKM1uinQ3MKosY5dIbuxx7q6maNaQUzOLaMPuZ9hrj
s+PPRROa/y4gbzu4z1bRDRp7SQl5W33H30jzqlGj8es/00zZJGKP18vJf4CHBZbRTHToX4xIMkPS
wEx9T37e5nd5iZy90NUvgrhlFVDFpvXY7FobQEFOZIE7sNY3yNw3YwSHHqToyQiaKlrLCKWCBg1M
MnYbdghaBP6BbVB54+g0mWY7ZdUtln0dXxfK0+DYQWLe1TY18Xt5V3IsXJiUg65/hkeYaMHU2KKz
jmJ5pHkSiwUUb/dDQDvK4CZwMA/isuWD/OFo6FFnnX6qJeVP2pULqu8m7m8YN98Qz/dqvYdpLiYJ
X3x1JbwXJpiumSxclscg6szZNjVUD5RK/8x0msh8HyiuAtJnKgUOzZbYiRL+nxwfEPja3nHzqYBk
6l5TzIL0FUs50drycG/njE3dB1nXSuK9P4dNgiCxTFTfgeRrs7CxkYrbD+HW1bPLSH8HZ93cv9Qw
c9NOfG624a2nwDzVy6GI0PQgPdN2cwKL8DuPrA4bKIO8rZKpq0haN9E7EOh3PPMsfPBRaduvrTJK
dq927KuJVRmLJiBKycKXSoY5QWrZmZL3k6ftXeahQguvv56ORXvWtogvk911UYDmVYUQc4auOXyy
eBkWnBA6BlmumLg1KI9KV9bv7xlX/ehMPvuWFVUGuBCUQ8Ee1oYHOjKeUOgMNTnyfKgrfUxbDu44
/sgOYj8X1EB1ZiYjBQgLusTWXgiIPrvPXmQqMOn35FfeURzkUZL54x12f1dzRflnXiAY3f4dZGAO
uhW3yGTz9QAFPyqHcOcsz+FQu34izM/RX73/BIHGd9eXVquLuL49O2RaM8Y44V4OOEl8Lg3wonZV
cttTl8RyC7RbfgwWX6UoVhqA/i/PziaXnoYkd0J7CvSuxUAn379f3xoVjKrmPtNb77sLsOKwHTOi
K0R/lGmFGeCxJBXglLvw4kteOaMXe05aoc/hCgRJz/XOVgLSC7E1aMYq17VdBqV/Iqzm0OR5cqgJ
2NVo/DFyv3nsdZCAT1NEP3+5yGhdSfHbp2pSZO4rT8NHiPBDs4TpT7B966KgSe3/D5Krw0s92MAp
Usyu3WaKd8i7XjCZZGDDztLR/b7Us97ervJqqunb0igfPYAbtpV8cevo7PQHYnzjaPxQmwJjVHFA
rrJQI6QrUAVpvAVanaXaOMUxTcJoELWHRzJ7H69VP15R3iljc4LqLF/dve2HObzdSSr+itN2Jifo
OcDHMJtl8Y7M7NO2yyoiG9iTXBiSL7GV0mBwBipQnMqY1RgU3DBc2LeC5c2hTA7VLgtMZUcSAxJm
0ZTMRsz24xSYN1NDNKQOCHyY5jEkClkDBPAsEvCAHFHWZ4OT5842dgb0vLTgwYPafH9nvNR+xInI
+VeR6CNfjsdEVjn2pDKobuIBq9Gqct0EdBDF+D1NulkP2rN+ayoZO8EB+18sFIu2t3kD8/sfbsJH
+vplXPqVfe9BW5XuO+iLfogHsLdwbh3b4nqUe7fPrshmcJWDf2y+yjsp7M9Kn4TIDYiqtyjtV5zx
VA9Mb5FwdbqxJOc0VRbAwfPTjzmwr7gP7z9NiKERg1R6Wt2kZ7qTbSeVOtkFOpAK2nkJp7TFZwzA
IQvntyaS+njvIIKC3myUN+VhvOejIawDwNvzC3dFhS6M09oZ/ihz+mlOyokSJMNs7OD2hl2eGcAR
at3Bs+08TqBX0wFAzH6miPhLefLZvuoa01T80pNjSwsxkta5nusUVpGsnTcX5zqCluhBdwg2bhaD
3IoqREMEHEJqov8ZcJFaTOoO6oqnA0zpnxzWLIBpR8C1fDS+ig41k7ndlGv5EMbfAp0xwciv5es8
bGWdm1/rUFsloxfosneIzAXDEV0ifV7bzDaj9wCr2WkQ7F1189XokakgB2LJTlOtujw2RTpunN9q
riS9zYZv4siPOFNDF9rdboohbCinsMwkeuLYvgpzB0kMTu8W+6Pe9EvgXJvzuQCrkVpw5w74a5zz
xW/AFsdMKNodXhEIb77Ewh3oaB64fNTZ/DMDrV4SZW66J10JwsWBnIhSwgNAVFSqjBSdpmYlwuzR
v+iGoLl7Yx+ywrQ7Jox3TzJr0vokepYIk/u2r/tAz6PNQw7VI57XYuucLSAjPJJiEzH/ky8qPyIU
D2gBUGPHUfkUuFbudyPAifiODDPfYNQuGXtX7iI7Udp0mZzjoNPJeSFYg8s5yCdsaWAI+myooA5P
xD0zy1UzBbQ2v0UhFWZuNPuYNY1gHAHppgQAITvbM9tSruew6foikKkU3PHjxYdIP3i5ZH5kGZzC
mQR0JoXg1wsbYHZm3zwJqm+MFp8f3rjLYnebiPI6M9vb1NDAKSpbFsT32fgoX6GVHcYYsCl40KoC
xeuDP1BaF7uWkHgpRJ3Xe9prX16KlXXhwJ+sX1CwifzNz1XCrsuSpA9CAB/tdC0BCyhC5tFkLT4m
oLovw3LGAa54ZeBHV0TvoS+r4er8nBEFUN6lP7qnvfc2VI+DUk51GRZgRZ5eJknTOPTspULRVBsu
yN7855G5s0EqbHodiKjh6SGJAq24ea3C4oF6OygQhtKsCk3gd9FyYtvOlvVZmkreJWKM97y2zLT+
uT95s05LrSR8qdBQAJT158VxPrgPEkAbdzrJ/m/NZJXzqh/kNPJjs6OlF2/Qqpmwrbon6/GU0Zyo
wPu7/0JQql0ZBnhHJnp1bHLFoaizw2dhzyxdHur3GVVW/EwOSrOVqrhPOc+2IdGzY62x+66kuITL
dH+OAuxjxiI4LgNQeveFNbw7OCy9SPrbMHR4T+wXEXSL17cVxNGs4fGa707/MmzrXQlemc8XOMuT
5AQ25rKk/I0MFFoTS4Q8q/TVF0D7HAm3jrC/mjGH/BnaKd1VpyH3ydhKjIOlMlqEn4X8OmTvsEf4
G7ptTpu/MkDFGR6UMYa1yNTAOjGDME/vq8jkaO4fe3ZVj0DkvyNrksCiQ40dZmbS/k69Ox6xb61v
eGfX0DLxDvQRbM4hW27ZGEJNaDaC5ic9arPGO2alnC5gXlgxrR6B2SisnwroTiaMaSs+sBjV+uCm
y+7l/R3FWoFyFEWRfEiP2uxtRDI+PJklpDvGBzWP1PyV5calEcLgYoR8azvxvfnMYKmFVhLz0eak
ax7zsgQ1P9SAgwXKiDvKVhBDW2XLHeSLdhrQBpMOai6Zl14wjZvTqdFXhdbTk3LNtQOJv4sLZJti
f2IyJhwA6XoC/rhYE18EXW5ZXifEsfBn4xvCuqqkyuQjyFQSs0M8CdWEd8CIJm1ois/mEOr3LyxJ
wtIyplgfVhlW0Qsu/K4GAwztNulTCaH+qTBBDVII4ch/ou7jdQE67h2O/JUW9T8fy2Fe7oGwd29t
su8u0jFWfqeDUt9Zm90TN/e+Jahfl0UEsPsZ9xa26LgxEOgekqBGS1jyTCWFn8NvT1WR4YOhLI2Z
/JEApCRVrF2BuiPP9zFbFk1IHexKpruRTUPTX+JGblLWpSLDTMoCccwYgHCZvzrlOVhtk6iUOrym
VWHtRMkpvahu3YdYRX4i+Pglscil8FIGnqO0gghWALULZDwUNokdgxaXnjBndOEt0WPY5s2IIUap
KAegrOXMqvBWmZTWxPgoXR99XD7RGErTbUt7Z64gsHR+WgTRySZv6gGaMQD/54p1qoN4r+FQ/k6G
ta0I5Lan4H8s1L91shOiPzDIiATCoGV629/3zmBrnLyy23uNKNdutYrus9QyxQMXP/zHfjO/LWVn
NMRXVEEE+pOzN9lCPrvaDbsFDVTUX+0NwRg6vhD5GO96gHl6gKQCbTjY+yM0lZg8eQ/qE4EamaRk
hPIWAyXEvexrkcjVeK3JJh4Uievmvvm4fZYxNfViB73gHoGMH5D4PEUyhkfq+Ap9uk8DTca16koH
p8ALGdsWn5XzI0hWsfhtvgt/XwtdlYvCWq3dPbm2eJYbAInr2lKhq/q23O3OcJ/xq2BTMRkSkq5x
mwwrThHAxyqeSj9ZWIuHw5kyxRF7b61IC8xROD0/clFpWDeFEcNr8wjjMvrXbKpWjydueslEKMzt
YLwbBgACvvjMaZXfhlBPbsfY2cr2AgSsgVQmwzjQGtfGAXAM8TKcalaKORtv40MsV8JEivh1SiQk
x4E/papXHxlNGT+bTWf/48aFMA59rDCiSXxCME0F5v6H+kCJWzbg+gvZncJpeImUh6QzyPc7tk+L
CmZt7G03NKEmZx3ijuM8b/IVSFNB8pKv6qQ0P5GATMg5FTsEV5rNd7/Jl3xHhDUV3YdolO69L9Sp
tugadmN/DE33hwKO81ahTUObdgGfYxTI1QS/U2mQYVoWyw3Aej6fPXG8KIpFeURqpqO527zuiHZg
c+mhJPNpihCZUdow6sopnIYARZAlii+0m54y9peeUZrVgveXmFYc8Zky+7z0++2sN4RzjpRAdkBt
oulgbGncuy5gHhc+U316Si4GpqAKDjL/tKSMmRWq5sEo6da+Srua+0nhcyeixZUEaV+JeE9PIXGW
hqvA8RSszlw9eLv6ZZcX6wExfX6GtEniqKKXGXv7mTRQrM7aWSr634AOhiF8AIWS76L2wpXlg0/7
QZG5+9MEiwbDfB0jeFo6qhQhi4CX36kiAhxFXcXZShSzoGP+cVAF6ryvn/dBDotZC4y0Yw5nkaA9
iwRqGDsi9YtFukyvygtJSKoM33MmtGYdbRDHZJn3q1/o6QpcEfTZbDqvKrRoii5WESy0QReB/Xbh
w0goDoNumG+pkkxo/evtdfuFJmfIs1DYeyEqQkeGcsdMOKiE6NWIqPRS3n8LP+pquy4Wne9wmitG
UkElvswjG6ybbjPUBPU8blfdYEQ2+9RX51cMih9k93KwSPfRoAby+Zo4M6nPkpok4Qnbq/BzH8aG
KPcveJszk0J54zEIDfMoKSQ0rKgdKjux6UUZdPWuGV/40k2HZLxxap9gt1/0hdMJIZXB6Fq3CJY8
J8rSpCcDLoNzoGUu5u9zp1FshL9TKDsunJwiWv7UoNmiNDZZJfztC7MruQ0pHVlmmp9uFU2ec3zR
WzU09PBR+oWwAOTzBioike8UOIK3iXcWOXXrOnVCli8kWQ2FSyq3rjb7+rm8x9IlfIuvvzRU96XP
pMDs/YhRHkugwaIeO9gRiPrmQPGhvh5cvoc6i2mS+sUNI9OvbY3A26ImbUPCCGt/E+jBer5E3HNk
dDRsG2KZd1JYEUAYfH+F4+833G1dtXY6OmOlqKTs2c4cHwfPnymifzV6yZqQCSCaI9PkesHzksGg
B1Dh5Oik2LYALOVGWQnXnZ0W/l+cNrb2JOGxsFRqveMOn6Y7Hn1nU51JoGwm8JSsME8XL5cJpeZG
b1lT1M0z7bW14Kd03clZeo5XIUQW7WtN3rUfvKPUVlyXPULZEncegkPJvvQPMSSgJn+fMcL2MGtN
tS+kUO8dgITFD54WqD/gyKmlcPwPRvX+GhrkH7eR+/IsTiqgSWSlhEPoE8xrAzaEjZs1sZKtl6fB
J/gS9iAkG75SXhQ5A260Vh9TUux/3dKHPsHUxtW8db9Ld1p7IrazC5USt5TChxIfgp9siHV2syc8
HIb/HZ1qI5r7gCUXqeG4ggfB7/W2RIUPmrE/TKiU3f8UWawj4F660+brnxiEqK4fUyuI3CZ18cKm
TxOxcE4NqGfzwMDzf6EKNLVxOYBkntC1vWQ2+iDFPihmC/HDBi/0hKyd3kr1AEpQACKNkVSD2bai
XrcCXljI5vGkGbeaJCA8NJXfXGVaIqZA5tyG74NL/kFt77g1L0Fg7HOTrxZuP2j+9XXBQVofrqBS
j436oRUNAPAZj+N0VpY70prhzHM1LB3pZXY2yOGnWMOJCFIq98bHZVsGVf+OdZMO9akjPKXpt7I4
haRpuXiW4pxKgP1b27tnh2qupMsAk20JvdSgClLt+rZM6OM56hn6LyoJ7EQudO/fESwBufIDgHBm
EaHLMSLNQpRzvpgPajY/cD/TjNLsqV7W3wPLQ5buLV+pLNvkLD6X8AJILyzb3a0pEi4UE8oQfRjs
vAfySUsC/WKY33IhKMQVe2bXOSpXVLCmMYAJoqKbl6OCOqlQSGLHvR4X8tKk2pufZYLZXkQuQtsJ
MD9LnUd2x0mQ3qO+Fs3cDop8hJMD0UtgwiQ5wXuX2dti+V8VGES1MlRN5aLLajEM1LVUFAew/cVj
lQwGkp0pViVORiY4ICVVLf1RepYcRd+IGOkDDIUaroE/gugDVJLVykO8IzHWwegncPwopAnOH0pQ
K++AgCkP3uFsbNZaZzk0q/4rtKDIX3H7bp7FDs/E5Fhu0jciKW4hyqjWNkx5Q4UtmDbzLiTIYpsL
LDbfxjZFbX1Zgm2XdEmk9QVu+4sMlGOBRwtNMMC7ReeYW/SA2f2aOt/wbYfmzs/6gJhYQvdzk6GG
K7pJnrvbpB3ze9PhQMlrI5qdNEjvIbHdcUAjiOX0JssOAR+VwFvBCjMLekh3eWBmyJnOKEOxDNL1
LDO+2RgMzx1ECAQqLjcWXimoGTlqScL9mGfBB/aDyJCQNFhpKebaEpPtJVJr6u3OtVHGa9MKjIcn
DX08XvUi8VNPkh3Ht+M7f8LP/nDr1iFvr/OQgIA5pN8DzO7EAlE8CMQWLi+rxr6P6Z169M1zEJFf
RcMsVw35ukoDOn812Goku+o3T+I+jx8P9/YJbI+LGtGDsyl4V03fSpZPO6u98mgNeupmy5aLD9PL
vyZgvJWvrA9z3Wwnal4xqyEbIMwzQAvcWbvVdMfNYqkvDFBnLuRoKH9l4rDJyZEWKIJ/GaiueMBn
xyZ5JcDlWdRF627IYogm7nXnPoGh2IPHLZwWip4zcvW+xsZpovkS5upku5W+YWJRqRbkUD6gUZGS
HoYbZWVCgMCLSu0ur+/yvnmvTBvymBUZuX6lbfJ1A0O3yZ+XqU3la7SO/lr/a4BZuGGyoDxOLMB/
CBVhfXDtaLgvieULxiEDQFKGtjIWmIY2NDrOWqvScw8FuzN2/HOfftLdqzasY3hRqnHOIz+928lA
cTp8lPaCv/z355lXU0oDQFETxgFreSLluiiVtxseBTKwE/uBLCo9QOgHalrdY/cdGqYo2TDzrKok
NUyf9fzim3HLrWsixtMIkO9kJgrMt09sasWGhqulZ8xGbFvAUnAEzaO2rYcd3iy4BjxXexXgpE2i
oiC6pc0McU0rqUW2FjMTVtd1Rwx8f1onysQv2ULkFaJ5YO3bbAMMtMf6ZSad45jPR2iCxqHe0DKp
JL+fFI5IN1JwpZ7lLx8HELAUpi11zwgOF9VDeHKVd5syNOnZaNZz65WoacLrYA1/GB8t2FG7y+dg
NcJprH1cwxQv2njsk5WiRHTjpDm7IhysnDxvRkOrPRRI0OraqwoQkvGp7mp05Km6sx0DhrT3Dqn0
v/tnhq/spZlElF6UCL35uLJOztrCGYsfU1cAYkeFsJfLfReUt1zmUo7tdYVHa3xqXaD3CMQoaYQ9
+Y2G+qXHFk7SE5NZThsTkNTlqjvzkUzrvSF+tfuFCts36HZIkTY+Hd6e0zWdattVf07us4s1JlL0
GApxQwyGDZ3TMUxGJ7SnbLgRs01iRmAhHvrDDz2GRuP/vDIT5+5jppmY+w2l5p8CN/5SVnY6etHE
oVAdCNenYfaftNVRLjLen1iAAmjqIBxuEpxjD05e2dkrJSnZU7anecdMi6pJ8+LGINUsLJZ8wypF
62zx//e4Mna6Qfoqq1s8ecxqC5Xb5wXntjS8OHWxRVvwurzuZMg8kTb4gaa1cAt76d1RH672pTSd
hz6g+HEF+bVBk5pVFxVFERJukYQFYf1twpHzlwLSpR0shPR6tc4PNt9stxTmhvI6eBrLdTEH8IVv
DZ9xdn3B8XTS7LJ8hsu2/WnSFN7zvUd7Vmqiu36hDuBhlceLC/re2lB43A+fwiAeFjKiZDxAM/D4
43VlED6QgGq6LXuvD6fCalJuvgI3fhVMEJlMJk/XdLW7hW8u7K7/Sol3nwjpGY1OXCS/81Y0olrS
5rDHgQiD0vIl7ldLBgyjSPfryGNQVxbPQiBVI5vdvIsRLrWd/Eaz8yh8n03emTJc5r9J3IP/wl/Q
iy2V/kTRKNIp2n+bwEN/DaDoW+ty9rNYWEHe9BqQYUUpTyRBhVTERd4lanrKuJEblrS0/xghSF+E
zSvPI3kl49GycFxywgkQopGx2jiFLMdGr+mDfMJAE8Siz017YNlHkC7qqSYaAqzqP6nNXH5zbnpW
x6Emt/6azHL643dK/7ksDjKRF0XgjD7ETKhsC8Xb2Gwc8cP8yWBdBTcM/ZAxUq4WxgvYWMqffPFC
GGLRrNRLpGIyGKlp9jPdCAKYCp93AB56jVVt3qDww2vB4jA5FgJDH90ZsxTc1aL/A9gO5Qri/yBl
E+xeyrmcpk4Klr6VDJDtRtcTjWhG65E1v4bPlQ632BbFjjCCUD/Z5mZcd99gXJ4nROx/Pt6DX76f
KHq2aDTJMrX8gHVWxiA4KODh9A7NF2RMJLuOio09fMvXPdDrrphfLeRFnU3Ra1SFJh06Z2/01UGD
TkLqotpTLK6ihIlrR4Qeyw68FZfXje5QDMzYz2dci8LhtvdPyGOIkiZnqJDri3KV8FsEZSX7WlEj
KyR1iOCDVpAfRr2eVv4nWaTW1dFke8n9C0PjWJchmUS9xTBh/Z7idqH8r4oGOvAKBmnfinHjEcj/
Y2eLwQP07UyZasGPsHRA6mN1mAyMeMFn3j4gMulC7WLr0UBrA6jlbHwjjzUZqwJvfz4X9c1GcKV1
oS+Fkt+St9p7Yx6icpQzlLUG3DzuBsUY+tWyMkz4k9JndPpSS9Vo24VCK8o9dKiwnp2aAKInh87t
VTGJTksdqUr5xSA/YWAzV4nbWH+TSfWB9jHmoImtKxI0cZARrP4IoRRnMi8QvNF0nz9S7QSDZZrO
ofXU0LJiw2nSvvZc5WrhZweGiil6g07GAuV2hFzeU0jBEPRXDOf8U86be/g0erOAFCzQgyjlzR81
1kLSxj7BgzOgZGKnob/QJKRBEFPbcnAms055YXXwV5oJ9ZToZMdSNsG0BkOf3syKutBAm0oFhOvo
VD/EQHGvi1RHhjlp93W7PkGap2TSYVKcAwlN+lcIjK2AyeK0QRZxCjJFJtk2/EGoUJeMAc3eI8rH
+hKAdCpPaWWBxYoy03rSNQEkVl0p08tHuWGuHEV+UZ2rs4sCl137DfWQeex3XxiAf9rkLB66JcNT
txQjdAMF7+Gki11IEbM09S2lmckK6stWUQFGfIsSWFyHCeje0Sy8jYKG1/ah6n8rVZyM1DjBd5b5
mmhsWsDbrxu3oQI+fceUJ6K3iZhl/XZDqXnvoMGQiMoBrWZRDvQVhsAEbL6Y5xvgkCABldrocp8q
nbcr7xla5hN99UXUOzThJS8NvPxLQwzJH97IylAtr9wIIKptfIhBKzUEh2RO6tD8WXhzlsrk3pA0
4V8izO7MXikaL3N/eSbcUETI5dKMTk7B9sv9KjiNC0quoYIfnQLzdwHaFfGsqxQGAGdH3JaFxKuB
8xkkhx/NgKl9YVLZA6zsUBEgev68uRugNCzTWTA47qBtJuowpD7NSOkhFS2YwRwKhxmXC+Uaha1i
w7tv7OQmdjKKNckLNPxrogtIOkk6vSTuftiq8U147Jii0/qIDN9pjQbGTIaCb5VrLpLuOZChHl+3
w5LsxyTg8CqmrwnaWyL2J/+oNBVSShkgxydKR19jo5qcV3ub3r/FuqjVkrak97prIzZzF7KNd+g/
tqcMe9Vo8hAHHabUdj2C6oz14InVRx1zjYQ9DubTf80V6WwciP3pRHlVXoWk5VhdiMRVAU8M7HJ8
YHXYlPxLICt+87O2sE5WoUL5uH5+pGvvcB/CcDx8zpE41V9ybacBNE5O+0sG+CzevZnWXuj6bjWg
0mkzpz34YmV8rojDILjmb0tUPBkz8L1QU1Hy3Ugz151YdLKoUukPnZqH9mBX1BGJkJ+5m2TlZuF6
E8XXG1vQh+7wOu33/48FFP64vZNK03oFOXDo96aMpEvjGX31IBQIxFdBW/U1yKywzE898Ieasi1H
0kjjF+6Ma2OwKAo9xN8/7kRSAsnVQ/JEoN9/8uvKi+zHWPI0HXSjNk4aE+U92wDJaiDXMPBwYm0E
NH0DGovLFxL8fpP90/hAo9RfA7Q8NRE/Qy9x6RDWJBuU3AhQcsTOEGQmhAg/Q9jTv5oeimQIipYl
P1xu4/DIPRvimmJ6FugMRoDMYEMDHXaWUDzmI+XIcs554z4RtvV67n9pj1iyXJOqPk03EA3wCBwJ
lUfUo1U7FLfm7xKmJW3YsdvR0MvmTuh1ZG6j9jmEJ3kpPKh6yCgmvY5RL9t6WZ0GYMssh6asN1/I
H3M1L/rBvkPX2NQcHBqkksDwDlpHdqhg9D7Dxu4wosXeM4vaFSuP35HzfONf4xW2r/bG2eZwiAeS
1EgZY4/vUFx/CDhUc3/9w3Mj+Qcd1Ea/r2PDO3WXGuFhJqW5hUkd3hVcy4mTuXoTHezEGP/8CBfx
ZDVjFS4IuPT0+pI5yMC3HMlEi+6IKTDttX5oVe+LWtR/za1TYBghSfSRgCJ2KYE6BntxbpTjRekQ
8hv3EIU5OUIQM88zAIDsnti63zoq84NXBqmn9wmv+QEH1ZcQls7IuAUSXuQTUwB5yIqpo+BAQEDG
bvYKh8bxOYTNsELUFYVk467Cl7LWGRFW/V7OP7CJ36tbDBuGksjALvtBpUIhj6uVyqm/QdKXCgs+
xrqiUB14wq4UK2tWsMAu5HHMnBpRW8Vv/wAd69SnFm13ERTIihJ/jD/+j13sV2RV6nit1S2V+b1o
64Kh+qRD7SHa4LF6160IDhg5BfUclvbHtT6Iz7PXi8wxc14e0Azi4YHTA9T1OZfqXl11zcOLOp1j
KKzh6L/yw9H/muB9FBrbMQElF3aqD2UmjWk9L086izC2v2oT/3KSvQo4V1ZPqLNTQS4TNy6egj/h
O5xKrame0Eo8tXCms6s9wZch7XWr47h3U9I513J68aO34gh8Cubtx1Qd5kRJP7BmQlDzaEPaCChE
n+YbohLOjCeSQhfK5+/DkaeT7cHaV7FThPiTcx6Yz2SyUhrx335oeAwZ8EVHU0kvz3ftm3/Dv1M7
imQ0xPG9zFEw0jGLw0DO/UAL9JFU4jTsDMOyExGIVgDYomqRBD7Aapg5UT/pvL3JS2oqLbyUh/Wi
6Ns9HuvSCf3iO4Wp1c53YR0YPxUd9XwTqeb/wzbt9g3UsoOatfC/sY8vHWwjdxzgxZwNfvqRLuU/
fCqPq4EtMbxJznS1fwtkfmyej83xJeG46IF6q5qC4wjOIfaObbRgWZtHib+YxYQutUseu9HkVotx
6+YeL8OPMScgnlkSXebGejzRjwC6L61PRnOzWq0UXbwjF9hE1cIGP2URIWvCa6X+K2bdENe28wco
bsYe7EMLoDL3WVdeFqPovmAXI+bYzaRXOZp6pA8hc5vsy9/H2WuwmA1zVoSwGNY7w1U6t3Gkz3V+
gOAv20OCFuxdyMla2UutBPxZNagfIetrXYrQdmVo1a3h84UjVDwwKv83V2RwFNeeTthuTq3BBFvL
yOFaSIa7sBK/EgFeoF05U6I/vQqAACO3K+QXyKUlz0WmXYDagy7gzzfbde7+CsIlGAPM5x3zY2Sh
cN9OjKZj+ojz9LW+7Fou2FFjqNFA5KWXye4ur4tr+YX3iNYl8zAGvEokBH2/ljYo+rWi3ME8GMjW
jF2PPDjv5jYv9/g5yl9vBzKphRUgPtdNWqs+cXvz5V0SalTImQ6SE2Jr6+MVQ/e5wuM4fB71cO0L
XHD1221Ugf/+tjlENJzSSUA22toMATPpS5faGPZoIbbydmOLBlBZnF0vc5SnkK5Ow++/5tNqkVK2
8LODZ2OyvTKDKZg8dp0qm4GVfjTKVMTwjX74si8QhokTaL9SXipZRX0epGHR2op+fdJDOEEKT7Vx
GGtYOe7c69zwI05P03p0hq1EnwWwCu7Wm5l+F7uH+x5hzRboOwSVnmUNt4YL+oadiyOQt/hRr/j7
i9G7WzskIETueSgwAzebULBKZMkqSdzNPEY2End6MlzsLRDuShg/0BjRqhwQSm8mCapb62h7jU7m
kFr8YIe1aWRTOWuPoJUhz2bixaBzD4+c25Ma2zt3TdZQPCGatxU27m2mgoW2wDZzZtZ8QBajrvDv
lNcwfDW4rBUwVtedeq5fSoUNhwA12HewrB0LOAvMP7H6k7gOrE4EBqO1sEaOJM0FI3y6RQRFnrgu
Ya/xLjKK0wuPHU/FOR7CgtBiFDjK/nODVJkdvRB2PqwJtu3bZ3563cQKfVZxOKYrCuztP+J1O5gT
Kd15enZdvL9Re89iAbBAY5lYZkC3lMk6M1baT38vf0MDMUSfFWeYay0XpbefNCQyCM/gfDsfwRXt
4TLGNN6Q+Ug1voZVQKxNk523lV/ugMZeTfOR5GYnP41YeZmEEcppMWOWPkPIvaDpH41V07pzR6yf
ZSfCp2aitSwdEF1kDr87Fb6DODBJL0pZw3u3k8scPxHnL/ubPVNKpMKCV+Uc+C4A2XYJtCc09S5b
L/OxJEEvviGlNUWJEOFOwzgm8Ra7IIByWkTdsc4YEKArV16Nnvb513j2zrsEPMwMiDIpGwfeAH6c
32Ci4ZWCcH+Totz3n84WnP3xpZwGGaW4cIjvKAnKp1cORprLgqEe8Y2r8bw7/LT1gBs1robq1b7B
ClEmEX88lp4gJRTtCd+aj22xyuFT0H3bQ8E3+HCT9ndH5VKBpWiskK0+Cjk2HP61ySuNFTjIlcY7
RJiKV7U4EmJpqofl+hgPZdth4KyzhEP/9dkuSplC66AypacAd6diAjBWiHi2f1L9YZi06Z0dQiPj
hRZEZHTmylp+EJ8YB8X0kMQsv2V2DNF8Yjj6Vdy6zg+t7PTAJXki9EkJrRVHvtK9mt+5z3UcB/n8
2Zc4w4/PCFFfmmyJLmr31QRLrabdXWqXAJvw7PDAITQ1qB3yShYyJ5F0EtES1hPLTxvvhViYwvNQ
aQXKYwcyaCL/IgLEO+otM6x3uMZHEHBtXafNp5ChoLQPWVmpU5WD87AIK3m5ETu1jh7NlMIxHBfP
4iHSYdsPs1yezMA52wGZ0pOfy0i9RCPghlS3pxvjJYmN1mCJ16ZQ633AU/8t4n+XAi7nSw5+0hZS
5Hva1wyL4gQkQDQLwI/DuUKrpce8PHRV4azlUPmP8WGdEASap6alqF586Rw/Sj5hw+oz1u8a9dtT
kvQ6QC9eY5H45rbq2V00gmpkVFiuRqCozwWu64XTgi7Cz0ATzIZQAqLHQDxonCI+Z5gUuBLeG7Az
M9kq+bKtAzg1vQ1HAUjcDFeqdV1F9VfBSYXDSsd+Q5fHSQfsu22l7ufjMrLbMyqJ0nsYrbfw8qmV
FX7zaw8FMjc1b+7B3n/OYnqhnddx5JxA/hmYLb93BriKfGBGmgJeVNCVdBXl13kHMANzwOX+ymrt
mbMerRLvHdVLcYXpvUOpTb5kQm/31eabiFLfzP4GgOjKReYHFeep+1S/uUucU8Io9QTLJwmTKQla
myqEgh4bwrpTnauLzzfhetTBgpBh7yZ2T03DoRLT2a94F2dtdc8qB+OcmOr6KhPA00yTSSCNl7AD
sjGdrFdB8FOPth3yDVk5dHXGzV3xnSPX1Ei7GVv8nAUGaHVvDAZMMjsomjDfHjdGEm1bDAuOdoXW
r/pGBhbaG4gp4RwY5MO06Z4ofZpiiZ/PvrjY5SMpslWE43l1djP2sNL+gwQi5G8BFRxBvzc2ObF0
4LhpSnUQmznPr/h4iQli9LHjSy5sieO0uiiAskz5eAF+o4dOazVnSA7jIV+T0G7OJp1W+PxeWZUS
T08SHa5+6jAMEHqlvE7i2oRC+UsvFEBjQ5Rp1AQQzG2hrH/y81N2SbB9oSluEXShFZxsvzL55L5Q
HyRs2mdmiPhhjgSBqPhMtK2sUxAoHiPf+NFBJzqEdOITKaXZzYCfgwTct7bhgVC7ZzO8ZCngkuyA
3SIOGwYkRzfjE5cQfIFLFnNHC2RcROyXk7disnmDW4EIAT46bla+mucyjVvNVM9OkCqCMcQHdHo0
iHfXuo8YH+INj6/Q5Hu5QKotsIzJuBLayDcGXS4MBcMH6rqM0TdEnzawEdc/3lpP3pM/cr+txQfD
j1G50ZJIVJmoLLESpsFzv2vz+caaLeXbqYZI/e0GAWUuktWbVHjZg5dSmrMS9xBillZ07GlpHx82
M3GMV0F7MM2YHZ0nqbDa2u5I1xmhT8OKZ+8o4Aom8c9tdii+66dYsK0nLAykM5nZdYlRgtaCQavh
PRMKNc43crbCLC7SjB8D2xs3kMiNIW5UrH4oUfCBxTsBKHdxA7K5tyefDLzoJ+rZKi0LT8gEuAWz
WvR64WH6qNVeMMRzuc6YbB2V2Pt8sdf21GLOWzt8ZJdxsN60nBPkQkkHQswiHv/xtJZANt1D9p+o
RWjiIRmTCo9PnB1xUodUM9fChsRhxIKVjr1gra7cbaFO1YlqCtwxhlpfb0wrVKP+ebx2zvkhqYDD
IwBu3kLzHOj/M3HeB1OZ/FmNO3Aa4NzHr/FQl3Dc05bADyuJL5gOo4jxZrF/mmHcDxlOzLgAO5k6
d+mlRmKQf2NpKz4T/LiUM53MqW3dRbFKLDTIlapjbPqMXJGhFRSAa4vY8wrmATZ+QVGMO+TxQ88Q
qU6Fpl5ELa7jMofLtkF2+5vIu1YUI5buf9ZYdNNWOxTXH0omB7fKqdLQTd3LYOppjZGpvDr2UJWm
r5F+f880QxP3maArQXYs21nlTJAZ/8u8ZQ8OWYK5E4ULq0F7h7wJWFN/Apl9IscBz54XSyEKNXgY
U1/u7nKbnpxep6gkav6Dl5uRCRQA2ej5bISnokexiMUSwGhMFoD7pbZtpFWqg76dVKSJPqp8qBEY
WK8EgzE8xlWefJ/xdyKTvSslpydezxz+BO1IhDqrwLihSt742QZzds8AwrDQz5k4OxOC5t5RXpSW
maqW0PrR76h8IrMHpwGA+Tg7oCYigI9O+Bn+PGfaH2yiNrLdGpHyeIy4Grotaw142j4qDif3x9YL
t7/mUCAM5mwlLqYKd0i2ij1Yvpni+ksfGsLD87L1nyj6bEjlrtFN3aO3VHmvk0XKF82roMc4Riek
Grd/nBHLwDJaCMrWumPysCV3TKTg27nWYjHWhoj2g0r1e0NyCYia1bliKhhvaJ4a2dlrJYBfx/B5
J53z/3Pmtfbyw70qS3+KcE4c0M0TaQtUeYN33Olhq810IrHWudA2cC83VHaTTAFKOe97iQDgct23
jN0iobgm3xanIZSyfQAz5LrDPh6WyPkfw8HojtjajfufQ0mnoeNf6Zu55twWS5CobzV3oAE/YWcp
OrpEYJj/IR+um4+XhX3kUoKcQT2PPQ8Sy8QadPfZSsvtYAuEHJyGQFS5IjQfBPKoWAymqTvgKwDV
kMrQhQNkessZqzbbZ73l5y0mFKfT1XlmJ8Z84veZgzTyzRVZllJmrWDnYPEIYnL+mrM7cpEAoTq8
cxis4ho4iTteM5MLWRQF4w5ib3iPI/jgPmyVAFs5In5FozpegwEttGJffD/kI/O5SwpBXf75/kqa
O/OfwNMqbKkAM333NkmyiX0il+ErYIu5/G1E3O8GB3u6FGsIlD4tpMbqfTSit8viYKOsTKoMevQT
Zu7Y4WUkJiQxbjI/uRTkrp3hLACCS3TGw1aBFNKQDhfZmwJRoZr1zTmzCSPPopzjdyHbHedHj4CL
Iv/YKVWQNbVOZErqE5nkB7hF++bub5majyOUE+wNEouzKk6fOvTvD/zq2Igc/9MsUjzNLtU5ZttY
n6eJNAmxPK+5I1K/tpq6to7DSWrhkUl46wBYoKdGePxGMCc8znQml3+5aF2r/EZiuv8UAzlFWch/
whNFL3rmG5j6jf/llQJWq2lyU8z0CEO5pF/9x+T8QV8M4SlUsF63yFm0gwXJewoZmvmHF/sixYA+
0nfN04Nr3zu9MPs7Ty4phFzHkJtWdnVarKovHypyHPpbAFRfGPz2qqH8p/YXklcv0xy+YklIau5z
tvY7ElZbFOFJk5VaOTwomvr6jJk3SsQPXb27xaV+J70t4FZcdaKOHxx0csAsMx7MWZbndnrF7VKV
9ZUXeYFA3NYRymUFVx5hzrQaVvIVo3ptnFf/fekTkdWtPdo0WajuJIR18LN5/UddNwxalvPeUbsg
EGzw/BiDHadPyK8ux3olbTxCAiC8A4Dzb/uyROu97G/CObBiE3NDbreBWb9SyLhgo1rpHJM7UQuQ
9n9dER9KmnfYADLw5/+zluYcAW1W3xG6oQMEBBHIUVTCYmD8ZWFzJOj+nOZR0Y/IkP3uyiORDNiQ
PdGPhdLiBTfYvW96nyda7yI1NAb7KOhnqGgtAU8KnctjMTN95ICXK29fCWGXwQfw3ljL2R7CYhYr
jDUwhl8rUu0OEIy/bPjhmQtuxJ0SDB7jt0tf25ehqmeDc4rSJSIqm1x+FhtFPqf00uaSbfXT3kcj
b/WQ2S13OrlSQsRTsWZI0k06silmEimFX1bL2qbhBBCrTa+JxYNAbkM5Vy60TeMScsx5BR3JpXfQ
xA0UkBaP8n0+xYpxhatqVBNQfYqLr53eyV8a5J6vbVM8rY59nZh0bDGquqhKKOL21RFH9Zgc/BEl
PejQTrcybSTmEoLLTYPvUa+ZzNLH4hRVkZn8DjhMbPxIVEgcW5R/zLAbxwYqeELrOYnQ4UUQ3RKi
Z109FqtRZ4NUi5hPQJdyT1pclVt+TiqcyztI2lifXzWohCLpyGzAhVXa8vsVMUzZ/uBkIWcfKE/8
ZuTRaFyHCyZNsWekq3MXQGQlzxt25TnznBpuFJ+wvTyKkhfAV1toY5XmiuWhagJ0Ri0mk5hz42OB
YkHbtrSTPpJznk8HoG6Qsk0juav7k4qwdgbgLgOQira3HT3lSxx8DX6bq88TYxNDSar1KbD8M3q1
1XDBW0la1uY+PpRYFiQtT36auT4+GNPAoCNYbQDeYLiQPqKRjrMOUNNv3Ow7VjGhckz8NjNbZCK3
muOFgRbtVdLkGGAkyynIF1/KCh+YZmew4y37S1IH9RQsriyAXWEg4wuxrJAIzRVYfRCtG0E6hi4t
0eLQoi4KBdieFVqSWXBUWSRL4rVf7NH0ZRN8zaYnfgaOooj2+UnVDDoq3EG9OabENeS5mv7Vqfmb
OwLYriK96xa3w6b+BUJb0YVh7D8UA3Q+VFP1+L8zZDkyu3c3GKXrLlXbJPCjFrk7sL6kg2Vvd7+G
ouTauZm/bRDv+bm3m0+XifgNZSZ1E0z+p6IS1oGmwf5qjcPUZF1M2kxoJA2cLPdFLbJY10GjEAQP
CiNT74AtLyw2Cc8CJYV+/yzszbUR+L5yYLLf2XIqqM+ec5d6TRDSxRyQQAb/EsUIPPk+AC2V7ROg
S+GDajHmnOtlxC9oD+/Sbj79zWtZBLCW9KgS4xhOLglypV8M9fydyrZJGQ/gmq/8B2UKjzKO+wEz
qJyvMobEu3MyRv9x85qzDw+qymym5JPDxy9ODSr4kOZup4RXoNcIJYYzEUR2By1BsgLQdKghgJJj
HsJd2AkBgpKnpud7qH7RQxBTLWpvRro2pXP1BvqPlfSBYOANUtsvHNv1362hUQc3s9jnOzVQ5EoY
1fsnDoFihtW7SuUGTCrusCYRWr2e8nLuGMPR3OhGUXmUF8B5RrzwGYICmVB9mmSe9XODaVp5j3Bl
VzEs0GVyezMgmhSBLqqqnKbynvNvd+Xx+TRo7k184+bTgozxiKOGWBfYwM8z9DOjXRyOacXqhH3m
Pi1Aiu04KAsdZpH/WxLeHApmMjtwhau2FbCv4zY3TGXHa2Pm/NxCxaVluuhyYyYfoWualHqagk0G
JTINCJyvQNDmH4KTxTKTW56CCEADjdLbH2Az/r1ig20hmyi9yIql5HJozMHOpPvOaWK6a0v2QgpE
NbIVaaxFK92JMnqJGua66vjHASYD1qrSFvTcMOvij5Z8nFeaG3gR80O1Frtn6cGqIkd/AFTRs6H1
FkgvmrkFOaOYtwwt8wekg30gUXjDsJWVEg3rSFblwTATHBnZ7bW5nLZO4KKxeLGYgYiLRrQ6iETI
GlBp7Ka9tFxHSyqlePVDGTPPw8TK5xxhqkI0oIYJgGb+rsnZpd70KHr8H2znZ98e62ffFyCK/BTI
519kK7paSs8arT7cAcx6NL+c5IlZXBeRFnwLrCwMHymt5pPoYJuVWKqDdEfOGJ9MUN199jA380Fp
oTmdZh6loCBRIvXYlNQof8i9Fuh90mGLAhVAYwXriYmZIf5huoZ9zuWTFOzHN1z3m0UVm2Sj9/gM
6r28JhIgRB+90Jw3NC9aKfx5EL7oZylrBqql6uDgjbEfpZtNmFVWIAXU8wxnOLz4lYCrNEfj2YsJ
epQe5nfh8gWRPYI2549u1H62k12dyagc01kcmtvNdTUiNyCWfsSlpPGmrqL0iGv2iibRC5HMZNrI
s6WMjMHl4IfQougzTTKSu68a0gWOgEb2s7UqX9be81jIogDc3+yMCI0nGTQEDlRlKlasNJtVnZtm
KTsNEUPRNdZr0I5KNv3RMNcqB9LflsY3BFYnjf7H4iKHg6HJwxocl3mXVw/vePQBoTIkK2OkXGkg
b/Yj2miwwJVCIeS7uvfMaXB4duAEfdT+irfzXG2mue0hvp2lM+1U5AYujZRgL/xSelG9TGDHKuOc
Fa2hwlvUrlS+mxvaQqyRAhTCxCjmYUyoSl9qVTcgGMLzEHnQaHoDrSuaId8b4QbIDOl+xlOYv8UK
L5TjvJlyW8OT/YXOANRutjXKf4UnO7aTKfPE/DX8/ZUJzhkKgy49nYQeUrrqtJ1oHBeMOWzK4xJl
8bnoLVQyNS4ql5HDsS0i6YNmxSTBgK/HiokO0RTjKACIEqTdz3IYePM1g4x7uMy5hFPe9xXMbalc
ekN8ka+iwLsGhQ3ForBbOIgEsniV4/N57rViLftgVFIuHBJjMSyqON13xRgazh1fapY7RBg+SUFJ
UWfbOakIONQFmAw5/uv+xgwsfspcWlUFfhl+YEnEf00xOa3qbwRBUTu9y4Shsj24rY8sXjWOExUG
MrGYnY+nvyGAzHronQgwz4BlXHleDUyLUpGywQOuMQyhKWzUpuVVnYH8Kl/9Z2gSgF282l2sTAwc
Xil8+387OsRyy015W+UrSJZfQqGfHSlUqf5BUWmVdb7f/jZayfXsVVrzzZWillZcUYYqIxAU6nc0
f1/DKJzfcAXyg/SlcMOthOM9FGf0BdzrimbVw/wv5Jhr44elYwU8PJa+adc1uZifWZCaNnX1FT81
sn3pxi/5XWlXcmN5snY6m08iP6QAc+rUV2WUiUW5adNgvdYfIVtBrdzBMXSwqzmpTh1I+t51Ex7Q
Jef5bknZRWGhemXaGH9emR8oq5lyJWFc9WwyxctrT6mafxkdQeL/sVTJDqnWXS6x1rCJpeeAwuIo
QKBqRT7oUFB+GMYBMiRsqolWZzEzIual0qo/z3CnOxwbh7JvpaNMJQ04qgJkcm4JDqST32JPYmMW
gtV5t67FV7Gl8S+129ndVKiucSeXRquU8Mn8s5yH51KWwkpaVlH90eUhYnv8X9rwJCW9OnCQsrds
W8IT8AjSHdEK8wuVYhJSChVti+jwXLqwuF523+I4D61eMps8rTBxQ+oRshi/0PVaJPpwNIe/aSwt
31zmThzyW17XHZcv2yBe5DZu7i0QODrP3MY/tI1xweg0fKAFyAsbTd3RXVU4iPNG6EZ7YZQTwBIU
fYFG2ZGtZPcn7e72upakmRwF+BR6/wDSgxWyBbzV3Kym+WUF0xhldD9VE6bzArLIXIJsvDNq5R8c
PC9OtyCcYOU5rNvxlVHNM+XPbVnQQoO6fBNpvHYHYPIHB4xl3UVnWbbwQzu5Q9M5mW/1Smc3siVn
KCui+HtYVLM2760swciLzZRcAMCFkFydT4SUV786pz0AB9E4oDPKpikG82ukoH7WzRaqzF9eJntq
VW1VA15lsdMR2oU8wsg/wsK+9cYWusvCyyyANPxzrKWQ7gntL5jrcWlUAj6pTJhLpccNDYPi2TkX
P1mO31O+ejMoTkBzKp0rmxfQuP4i1kMoubEIU3lLZQOBvKPrACCUjB8ABV2EKBnAr+GlMC2HZKnV
08SJ9nUd9+qqOlgA6EXdzE+6CQVq1ZC/o2AfrOegyMrIpsZUeqz7rfAltMptN5U+lmchO+4mMrj6
GMEWMIVwqVScFRyVTQNpO+e2PSBHhTyWY2IAjtKjnun8jxULcjHa2xfwsiaT1S+3xUYxakn86Sjt
oBQM33tQWqi6QEM8MY2e5hnoy39Y4mmi/zSgw9GKGgBS3EUzb9Lqek9ZH3I4/8lCqIKnVviSPwWX
2wIPxXazS+1nRJTOuZUsewn3HXDcTsCqsC11Ywr0l7TgHqKMjVbloT/lSkfu2S2hgX8JqVB2+Ms+
Uj0g+6TipXP/BbO8UW6ivLpuU+3sECbnZnz9PTjTZlnNk9J4DflFXCac8w3MEF11Z+kn1/5i7Q51
95Lvy+tNkQRZzI2Z5+14TPgAavJi+XgNvOs/lns5WhLBDVRvgWWwDJXjg2aYsZm7ZwdfArrXOmUP
AQ7s+Su3EGWxFH0ejgZ6YTESCkWvkHSjG4Fk1Q5iCRYrjrZkqqE4ZQXQz0XG9aOEe+ADtY0sLe2L
k8i3donMZWWH6Lui7h6WbOFzGjU2vDqubE0ak7x4n2QJpTVOtTmykzI453+TJRzdykv4fGs4jIyj
/N8UQIh+IQdA8o1TyueR8ZhFfbfgGsCe3CmBOQwiC43xtzvYtVNNNpB1KN2Ag7IfqD3wXgIy7YZu
nsVt67K/bEie+yjxW2bNIzdHQqXXYtVYCyM2qaEUFoqQBZHbwtzi/sUwL7jkLppHApPXFmZmMkSl
9M86avTJGiXr2z7LETQWH/oY+7K9+KU2BHypm4pwLYRjPufg913lzKuZwidpVGmW4ydn8mVR8Ope
C3X2JEjDnKT0ShgzUUHZXfWQheknOyO6Sdf5ggwIjsSKUzPtSLsdy78WS3EZgtmVAxSUli20vmR1
skImNndJB0JqIBnMAfngE9UxhNazm6AnL742+ED7RH3aGQGNvkvCx9K2uvoV/MB7ccejxOey2QSk
lEh5plRfbbSg/qgRNqB8WwbK8ToyQtwNbzXvF/iDyfm6jQnKIsfAZaWXrvilAENqUZG5yzd5qAKa
WiyBg/mgTSLxlYCdPx92ob3x7yqzU+VVbFXOtsJyKBdLW80PVLIS8O0O99oVQZcir+uPI2csN04p
/zXMAJGz3kYdFqZ49US8dkrHrjIrv9Z2eHlAYh4C7znup5SHgFK427TI/PMVc6jVuFcU1TUrZQWs
J4b0UjT4ttmswcMifT9oDEyCyi9Rh1bMGzq6gDHvRV1BTKSh7VphR53xuupppgafeTId86AIfWuG
k0NtuwxLAeMeWm1ZxJfpCvXf5dL1lv273s80DmBw5KfKNHUfhlMcYj85e7zuE+xC9lVe9RrVTQb6
UCfqQ5up1X5vGnLjFxPajpG4dJ+oXCW0hIN+hGi7/SPYBJ5JSb77Fg4sdVFPgQDQenskNBU6TG0y
Sy+Zo2PnSCg0EXF3llIjH7XAua8sS+V8nRcDOAVfNN/XQayMJ8An4vPs/Hyx6aZcieKUjIFmZBqS
Pcq+d+HIZbpMGVOPzQsPNo+8fkIN9SffE6eVZl0JjxFj1Y7jcMtFxabMU0Y/s4uyXB0rePYEaIQU
6wfnzHpKNJtUi7sMVfgx8LOX3PHZFG7hpiiYg614WBW4xrb2CneGBo1yh+ABVa3sNh/p7q+EVoRW
0csikdfJ72eHDj7zoZi7kBF5zhBw69D3VFvOm6rRfUgOrnhIteHpilLohXy/PeNmSVrmLr0oEuVe
MAN8HDITzigUPpVVHZ8VuJeoPT3v+44o6osH7VZTSC6ieC8NWmAQ70hrA5NajZyph/mvo3IGN86/
EbQlUpIKrpoHD6QUyZ0cGPbb270oPiYvsdR+bGMkPLCv7VcOav/K6C21nd0Txn80/nwW5f6Zljyg
fpuG+E5pCuCvgA9ZM9tgXn2S6ktT+wfNFiwrX/JV29nAyryitOLTNhj3VsDPuTzRD20QuqbUieBt
7nhkr14TSXDr4Q28DRu5gwqhcnBkZ1XTq+xdSWH4BcMCkmyVhhLfb7f9Hm5DlSC7psUydqX7VyX+
1IzlGnYveduCUbdb6kKurNKpiZlztV8RmqcRgXtGBMTsbVw9r/R/1zhjCgbURO6aZny6uIl3IIFn
s/gUH4PBJaf9iP09U/QQ67vcJhgjK0e+nJqc7ZM2ZD/s7WLrH4Y7ksyYYFBdrMWwNF6cVrduBPPR
wazIo5C2j6Zhww2r6VVHRl39qO43fom3xXTeCtk/gXc98RPUkjX44Ua4OEG0NbToJVV0OL6L28pH
f+A7t3U020OhE9+Pmaq9fhY7F4DQp5GsmanEyqDOL0bTLJsfzH5zSFxd9SjduUcP2Xg6cOzACQhm
mGGYj4Bx1TNc6U+OLbO8XSSBQFxGzYZP/lGNEPePLB4NogcIA0FqzHkrvlBmhLVvi+YQIVO4/KMy
BD0bFUttV90YTvEVDvTku/+6TxA4vvFtZGstBaTbGdhK5DLtsLF6A6MY+4JxLsOCEHqLGEzdJ52G
/j5ZeI48lw2N/jJ/sdGZ40SsDi+bogwoJPjjMBpDmVfw+30x3lelGpsyrKqLuYlll/Hfu5gwwBE4
l+0VxKlT9s3lYtkt2CzAOcSeekmWTlA4VP5Nwu+69fFUCQjXMaF4PspSvV4fZsqUg9HPmCV4ANZe
srkMqZLuIdyWaGdqL6GKAPNaNULc34hP+AppFdQOGBzrCO71rkOEGjZp87J84RCSmVN6XU+mabfJ
xsZmqFLkT0YhZzNl08m1gIN8cK5mw6SHxeffQR8qXwFVDOUb52AKmyUeKu2vUz6iUwGCe5S7ydMi
7T/3eBvnfn/VXrRkEAp4thKt5VtvA02VVPcC+D6vbaN2eJwWNWb9V/kWPqDP44GfE199eWAxSygM
a4ZRu6fgpXaKaOWKXhIFqdP4YOarhJXfQ41xF29JamSmOh4K2eiuLX0IB7m8K5mfwr/BfkxsaWU7
o7uf0uiOz6vaucdZd5gZOxXg8C9Id2mzt9jNQuz6lhdR5CnCrdaa+lxRou3zXN+OiCfcX+1SDEsZ
FSVLqu7ErxVxxAEDgk+Hu8XoiwP/pnsAph5FyRfEBrsguvmiApwmwss04JonLxHJCRCz8HUcs2A6
DWW6CfPsZGeXknAgRNx+7FidxM8NTcpBHFCwsiY9UwhEgIDW2a9sFEAWA09Eat03Yd9MY6NcgKPC
+PuN3IVo+gV6fuPdB22Bf/keuibTuMCHFnpfGVIoRDL/0TTBScsrBG2fgHtZb1PkvUhKO2mzk5AU
4BBPU3W4oGIJqHvyTedBKNtA4monyNb/CgzUA0WtLAtY2wfzyT8TtND6TPQig5+il3S36sU55tmp
go/7xo3HWMAA8kua4q7FDyiahXxF3eJx/MYnHYUqQJBJmv8hwZoSCQFLuzD1R8Nie4jso1vbgD2C
Wj4M6PhqijmTW6MDw2yk4M2UgRkAXY8EbtAU5VFmOZJ9qtysAQQ9T/gHkULzaQUNayduNJ/9UMjL
JqdzRkjsPeKIjQT1NvcId66cJ5fY/NhZ1/vPDaqIHCW73bZA02w3K0Jn2gIMnAEJtrcGfugGLLU/
vCQI6lQo4uAUy5sBvsD7I1qzyX3fT4wOSTCpYJDINdo7Az2RFpckc44VxA8mYJPUQmEQv2asbkY7
kac+JZfo+93k0Mw3eWSFedLx4JsaNmwE/aI0H9mmQQI64jora5utewnvm8qqmZVQnhTETljO9pzi
H58d1ILgJDo7JarpsUZ7ij2O74cPwRUJwfRsP2GIQDHq007n6f5Ev/aRPqNoFVDWweAFW8R4P1sS
K28sZvUM6HNnsehuNPLN+YQE8EMOP6At/BvI87A8tL2kk6Hy+CbhOmFPkEUij2sXNON5WnVmxbBc
x5jpQrJKixu3wfR2OxKphtSkT7iKMApqukrJase55dAF8NcIKnpcYwNuG8h2l2ScGc4m7SX5jAJR
oDZFp5aBbzxU9CAW/AZbbqzicaHNEuM6dabEkVOUzjexFTMMhDfl2cAJhoN/MUZfYe/tcMA3WMYZ
WLtk+XzBh1ERCY1garW9SpkpwBreTiYkaNU6cqvCkX5TVJWPi0ru/tBRwvwK5SN6f4SFkrEL0LT3
x+taRxJC1g83veNdgk1NK5oTKnbsmvL7snaHtPQ6QaZIhSwDyubnDTjn+oLdFMNXSpFsOtSqZ6qC
9x+BRnOJHhk5QRvrfaCJsx4RxOrklm7vMybs96P6WT35Ajwjr37q26Gp2jnzlHmjmQ7JcKx0uush
5tM5ElopFaedxTVDS/eJwpEQAzTVRedJ3XHuef+7PclwY6XLkmoO3y/i4d/DUbKZfoW913ECr0Pj
/puqDPn8Qr311c/SIi3Wb7m1DCCZw9M+iNhLxx3ObssI7pL1QkfMCreI1wOzIj6UIC9WgjmdMzBX
rNPrku5R+IAYF/TmAmVNqxEmiIpM6CqlJxtTyU7Aec0GbTS+o19u45ZGPIGlwI08KcuS8tiqrk/S
zCFKj/hmR73pVAo50nGhTNEAQ9IPa7bXssLgbEImHNgVmxN3rgikQcRjwgocEgubuEFYM6W2wziG
wH3M5jEFbF7pDMMq9MYa00AW/HL+CNXTnSpgV31ZcRn2R4qqclSVWu5wYb8r2vAQSL7QtUnBcgi0
6n+qReWEAGZXeJshfQ6kIrGjvizHxYWl/AbDnwmafXx9kyHGblSfK2/yJW8x8uTKUksS9by04nKI
w8Pzz5JImPC7eVC+0lmHEWG2+PKaelbTApjPPa5OW+rdjZAXyy/TxQ7Q6QAvlo3ehrDgEoO5M/dG
h9Q+8t/LewqymIYuavJOf6bcimuwza6AWc0MxPs0Hpu6YPOTYpXKph3jULNInoyRod0+C43sD1Y8
Gwi6p79NqgWgFL3qGPEte8sq//9BeCq5m1sSog37+Y9goCnjROCzk12MT7mSbMiJiT+uPmnMw38a
RElp366gQfPUH3NXmt2irXT0ECccsW/INg1ZHGcnLTy3p/VKast8YwlVUtFIMaeesCAbgTzobAKW
F/lxuVgZJb4R9k4qXNGa/gLdnCFtPp/wB60L2Nov36JadBFVot3dyjR1ng2h4dsLRhoYRo2frh+p
lOy9kq5Zyw++fc2maFn2kCYXOi6y9ie50L66A/gMF+fR5f23nPGbqV7n2pbQGdCSEFGYq82jjKgv
gYGUWyZULYCDzr4YvdBIuo6XswUCPqQIQlN6p8G7Ykp9eVaAIRjCUjGJ2dZ1JMqxi9SGn0zPLat0
ixJlYKZVcDlXwR3P0pQX3AIJuLZM1nCiG62YJuaYLmKxiY0+G5dFz/UXaNyaNOs8NcPdEYEu8PhI
RunsQhzQHl+VS0DS4a8LoE2ptI7A6GBRCWTfSakvT/BG22xP2i3WRBzl/4TPoRgZ8XEGdikQ2lIF
dO1ZiBhHb9wSmZafqkbLGqNn4CsDYZ9uAgo1bOdfkSoKZnS6xXN+HJ68/TfmM9mt72oYRzrr0wdG
nF4wiR+J7CLXGHGKnV2+q08n8nYA/ioDgqoo1culQqr4oSxSOfvsra+9pNlA3OyNqh4e0PoT5DwR
3ozCVpzopeFzoUuLN2guaYm+lOKg5Tvtlus9TjvTF0bkOps69C/9i3wLf1g+CU+1fLAM9MMrpYVL
HRwtYyzDrA/MSFXPuQziB8Ucf7fSYJAO+XalcQUPPoCaKlWCG93Z0Hi9fUk9S6IiHLZecBXAtTt8
HEjx/kZPexpgvOcFRim/aw0kLl0hM2F0IT7UlTdVqicCcC/oPUdz9+OVHNv/EutA2oEd9c4WeiWN
MVMuCsvq0GWaPDesyyqg6zR2kANCZrOCH5nybfkU2UJEaDwz9IPX3Sw8t1xTh0QiXMrgSf3Q4/mb
B9KCD0dmFl1pWK0aemESDZFvyo6h1IqrgaoilyJzQlCS6S57wb1b0jG1uSpQDVnX8qPD9nmWhLMe
AWzXev1+LY9fZ8ZdoEnXIolhIDv1JtabUgdGnTaJOHCZ4eHFfz8r5Jvoru6Z/Cles4TUJq0y7F/u
4d1N1BEDdVMlJZ8J+zKOQMlGYysoHqQRynzBZDP9atfE3x28EIdAgboPE6oGPt/U3AUlDwBwtKsk
5SGaMS2gQKdFKyXe7oC3wLkJ3kpyzbpQ2+3sPkNDW7vH04FWO0PUX3yeSszC45FuIzWoqnh25oFO
lgVqMG7IbclIXxLMcfik9dTeNFNUsfu6kooqRlxR4D8zdd96RVhA+L4zp4i1T5YOoMwQqKSTkWWY
qoO9r/zvY/QnEcUshWzz+ayjMsTk3zll10o2Hj856sq8xo3qImsDiSsM2MsTs4exkZETpFoTWuAb
qBM2ZZ19022b3EAOEatwt3PSfcOQGhCNCdciNjNak5yPSlE2Vu80AEFJ6K/8IXWSWy0uusjhC9Rl
LHG57aCTGIP6KynjY5BX5v+ESSlbKLeEbl4O347dTNvvIyy9c5svfcHl+tWMbyfoAir49pwVpdHV
l30tGq6rEp8sy42uijjNnJmNsKeaCxNWxd+WrZwHSfGcYQgiX4M+K9T10kmagaDY5U7O6StuBGV1
oKHH5V9GhDup/YoDfjc6xjhbY1J8/Ji0WyMOu4f0b6EsSYBuDOtp3NAPSsKwhN/VU+/rff/VB0nv
NaFRp+yyMQgXyEPvGLj/mGgTYSs+ElbOK16oV7MA1xg36O2VmFQl/0Z2lJiKonA8zn1c1EGON7MW
gIo7LRaKk++MBvj5mQvbvR2oaThmH2pM5k4lWZnfNV07wMjFQ6aXx6VCq5oJa0FiudzemitT/8ea
d5oQS3MVzvI/3LF32PQaeztqzJtrrgEMKB+j0otCsRGts1/rHjB88vNOAGKyF0wRzzcrGt/s9bwY
Zn3MQZBBsmBVGJieTI+JXf7wpGXvGtVYZWVLQkjG7QzwyNp2nrmkFPL3ckV8myCTU3VNLIotgmVX
Vz0VlxahoXjJW3N85c63WObayqLk8V/9atHGRcr49Krk1jZtF+IlFg5+igN+nSq2QZGNEz+PYjdh
v+8Bu76f6tWAoSAv9x/rgGn0I03xOJU9k2dAgvww4q1Own7wfTwv1e9BDQsZcB4g8hssXSA7EASF
soZrb2QCzutU92QjaAZJD+CAs+rmABtWmt7Dm21dHw2gLaBrtSh6jaFVzodkDLs9KXdZySGN8M2v
Vy55OBHawLcWZ2yKGWnbXc8CpDu8WKwjPGvHL3TtiFdodIQIJA2i/Y5CT5kP/g+YWF2R8qOqT4vp
UvaRDI6iaF1KJiIDBifY4oxvw5j3k0kFgIXClSA47p1LXVutKTxVDuR7D62oTTmmpTvwxo7NiraV
C2+VWG7n4OLO2ouc/5o/fWDy6UG3TDPjOK+J/sEEeSijWQp63PVboghMIZoN1TiIlwhOclEFAVLa
sjaBLg0DJTwHAgNtwFUo7GK8z+Vzgg5/p27m12L+gNfY/eIIaQ0OK1mSWvVxYgX45ro/7H7nVyzq
7HLWGjnPNlxaijvNEL+uEYWpb4bEqdEuew5K9/41uLv2Y0xrfgmW1wzHvF7fzDA0wpR5gbd3e2jb
mf7dY+u/hsOwhk+JdIZxqhBJtdKx8v53UoRKBbAugy9YvvIbJx9+EbRzvcA+hjiXqSmKvELuJkep
xS7xURsF/myy19QPpQsFewX+fYFXRnYNEKN/hcVyNAF6YsHTbodsK84kP8A6NFXE3HGFMDa9R4q1
P0irGeSbieB3tjmLLguOndpjFRXc67aBlvDfB9BaH4m6jMAFYI9tIcb8MEKxXXgSps56Du8mviyC
9tu2TNhHx/RqBE/VKhiWzX+/woHP7SgLV0lNx5cSNSqrSA+OvvSPCSsgPRZjf6uLaUuJZvw0NfLt
VU9n3dlpKeVPLS85PmGNMMDVRkGTU8RgPCxDyYY89RJ2wXEWrMt2vt7HACR9RByLkrvvrnMA401m
aJRc6r4np8vznwRmw6lOWbFUI8KLRsTNnbxiFJo8wM3kL6s1QOkJ1WiCpoJAJ/FM1gh+yXOCR4OI
+GqNFrDxP9SW+B94prtESzwVIRCSx1DPusaQOZjdXGovnoaFOGvS1pDiAxUdD1oVybV352IzcHet
Gcfm1DdAPkKY96xbDJ4SMuhM/D0hrQBTwfUQtyjehpf6Pe2BLjOHOBaejzysI9y1fEnKqlmaI3jk
9rA1sbNJt3NazcqcRiUBBxLIv1R+yNLjncVKug+HX5oT5cfAO9HE5Ku3b0ty2HjA78pwpa7/8/Mc
vlRmLPoMp5g9g0q2ax8WQtZ/n8Tkza0KNKRh58+ylcj5gACTGl9KNwheRcwyu3An1HNeX7QirdPp
1g6T+NBlokUX/5d8v7cJhvCzKNu0es8t9T6Yu9Xq+q0qhLWl4g/g1/FWdnP1OVXWrv9qfX5dnYR5
lNaYOX/QPtHX95bC81j4V4+49oJpdusMzW/91bKmCnVV8K+MIIV/C1Wanu8qY+HVHOmrASe3uxNz
E5h/+NN0cvH5xk/8J/+jPQ0Pr6/6HQaXagjH4RaVTjNOFrE3yCy2CWbrAK0uYvH1HfpTRlpaPiU4
rXWJGzW1R8Rg0fVQcFPQM9Vh/+i8EpKedi29zQEni9YZ7OlwtZaRRhONwn9SDnGUTbjyn+c6iJmL
JcsxPrfeDoFICaLIwjnm8zSn5gMm0nPvjCyN2lt6CmJ7GNVY5MfBXSpzuwXnsLqCMrb71C9AKVA/
lM+s8oHKlwLHimTTb4wTtrYnof+0pi85aGhzKfijYWVNW8P2bx9kLX1jvr2wv00u/jOCXHOnKqS/
gedCA5GnOd3RPEIcDeGAC8PkHxcJ6z+KZhNyDlfzMogCJnLeG7yFYDwv7rIAqQqSv8TLK1zCO3AJ
SGz/+ikmilhuakXsTiqTUJlsVVki3Jo13UFYtmvrjXL98CcscSD6cBJZgxvv0Kq8mOc0kNbVn9qz
mDG9lINSTydZ8VtZSsImeQS5hyO3h4eHQb4W9nTBWBiJrIArDdiewrcvr9pOysweH9xw8Wn427x7
k+GrS3KHarSlHGfYjHLtCyx7cAEYXGnMJXZh1W1gvTDTCmKreyzpCu4MHBZVoZvYqKzWUAUTdrYq
Yv47IVpq5Ugf4/Wdyq6KQay8XaUeda+6VI/HFtTgV2KaGdIDKPw5I882PAnZbK8n3tu6PrGugKWM
cWzQyU5GNzG+P+n/2GOcTvd2jGkFpl+CAPL3+ffR2fTKhz8a/O0VJRydSy9s2R+KHHhjbeDOCtGz
OzP2jYCcxUKYAh1wCru4903zXZUfwjPoKcXH7PzWwCG/QXsxPvsRvRa8PyXsYsqBij6KpUdA47ks
zNBsoD0rkBLXTX+z7AEdCq8yjJpzj2Xqa1eKBEQcyMkYUxsHGenP3rO2gW9tuo06eewtWOHGYw/l
d9OvSGbwymvjO5Je9JYEBWe3epDNbxieH6CN67JjFiCkWaqzRXeYohnrVJFDNuBiibBUXz3XiN5o
9Dvw5dNIJCTZBfFUoHUO4NxktCldrFeeka6I6d9ucHS1DZQqIAxhVAycx4MA1Ql1WK2gu+r6GDXk
YrvXwi97rWJXWhg/yfr5BEQAfwcdxrEx2qlp9PhEIRIqB0paGzQQqshlOcHzwtPd6ye8HjwJ/dUB
7vKrTQ+72umWsHlvoUODLy4QLrsXXxkgN0ySnlGjhEc1wufXyFAi8ikQkCdqbU4RxMt/yDVKASIY
cs9prkerxLiZsHEaIY7t2p0xMv6nuDsfaA7ftA9B5h6EKf8v7Ea4ZKgJyljfeZEATpmexbmBr7oN
V2upcD+I/WOMSM3DPwAJqehpvJ8OBz8l/EM8ZRw+StOFRIvC+dIoBxdKTwuhZ7tWAEORMBZtTVoc
AnTS9e81Am9MLRKwceriPAzNGRzA6YeVMD7VZTmZnHPB4zGD3tjOeuuknhQvlCt7hAMlVm1nC3UY
zQcYkMtpWFgrp6tssj9pECiH81iUlEowvu78V+nGv5+kBNue1sc2z5IsLOloM/6uJzTzdAzMcKJQ
Ua8kTav9BTkByNgfPYFh3qAUS1Btz140e2M9ShfwZUgwkUIplxMOaGRMxihs+AxHtlDeQvXiiDqU
H5TBoI8gw51Uv1DUAB/UN0ETzvyiOR65jwQjIU1newkJS+zPIl2XTOXCrJWOU6BXpDDaHSsT8ah+
BgImITcXyqRXulMN/MYEkmxFv6fhEDR0olCIUTSfroi8uSMYmXhLgySUkT/zQNPi+Tm4gmxMRbTz
9oR2w2Q8NbZhZ3aeubQh/1z8h5/C+PRUFXjkEKXLAzLYxBDaIgejKb9OMY7k8xWn/oUEbExFLRzj
F2GfNi6RgOf4au2R4WDl91QUryspgupzN2WYiS+fEZwqNeWFo7Asz6t0f3rlDBDq6LDlwWutsTPa
7CcNnhK1db+za85ZzxBg/vQjScVDh630OP7JEAT74FGEtfPyfrl6whGDCA7UYASQ1TKnnGYx1fd4
EZT/sKxJedlmJYIapZAooOFXyLh1WjURD/yN9SJVvnapGn07GEm/CXVD2BBFifMP6ax0kxuqgfat
EMpMux5wxnU/RVWAzcCm1ceqUMG4T7vpks4xVKrpjWQoQUHO4iI6+//2SB/ynMSUOb4CMXWPOvEb
Ts43+UUgCmpNN44NoUvkxqm3VefWoSVml7viQxr4Ce6eUf78kBYNBUCFUl1rulwZR1qfFSgL5plQ
Wn/cGcbSy3xk2lF7qO1ZE3xHElTTH1+aCtHzd5FWmyaU8SZZhMsUx9pWzGDKiHfBwva2ZRB81Gyt
0ZHEwXTDf3VYNjOEs7ZKPXxQrTiBsg0U56Xsy/y4k+4aXJ+Qtpe6oNI7VvJ83Oh+hnbn9OQVMBAx
LBCZGcCioK3yZ1qsMOn6V6N1WWnOuCeX3Olfvv/QdW299q+5EzRiYhQ8KL1p7dqVIMLcXgV3nIHI
ZpUxTNzn5jxpaX43ujhOmPMyA2TS+SIdrNHXX/kdS0O/uvU1zth8iCXB52nR3bs/C5ZEmb6z2HxP
vH7qx10d/SR3DT3s6a69Za51lkh4IwEsHQF+yZ2uB+c2xYBNcB07sF14M0KVOpenUuPth8ks/lk6
b7fI5YPWCshqTAn5uVGGdZzkvEI1vbZbTXfFuRS3e646TPM6RTkLRG2+oTEdhqtaYdAO+38scBoX
AKuRzfhRaKCZU49E0mHr4jLoP63YHB8yfoTkiAKDnWWg8q59dkkrzwW5LYpvHK4GD86NJnG9pppg
2jvHoGLAlJnIsCU/WfvFgtXk+bcgnk60bIFnMi9czLPbXzSFvPItQqT5p2Ca9BpndPdXLL+FIcqP
Qguat080/4kT9Z6ZqIzaU6WFywW6KgL/If9Pl3KAGy2pccOeeBh+aPaVom8rmCbKS8ciVE0E3K7C
tnH/ZSaCoUCXSW7Vg3zQGbEUK5HG7LDxmFZ9tN8yaM4ZnF++8/OeJBzpchG0Sg/q8ZUxNM1VcofF
/OuYFgHBuzgWtsad7DF3Z4e/MECO8YZtI5/l2d1h8O9o90faNDvIAEocRmJF42BIExBRB0mK/Z2o
ewLdmB8ueCO7SAz9wQ+7Vz7Jih+PgW8bodTWmjpm9vaGcFWuaz7KDesXaG0W/C/4nP69VoQAJVsm
hy4P5RKHC0mv7qkzH/KTzHmNf92pPQYgtqjS+YMTo7jH8e+6dk3Ozq/EBzXE1kkO2yRmS3ssPLBK
yZuLFT91/Jyx36TLXlpamGbfBOvS93/0CxFctTxHH6rPHiYzTw7Nr0zelgyl0CoaiRDavziMRyjE
bVftdcd/cOw+gLotRX8hRmE5EuJkn6XY8ZcoU9AiRGfrC45OyIWmHIQvInyAsypapKwINMomCV7e
ZGRVQuK/gYu7q3gECuJBe4gq3ikqQgMcgZiFChvEdDUT1VVPEZNMOjUvTDKl0VuyhBVM21PfrLYD
9xXwY2y6ZmM7d8i2tGTvfvy8v8tyejBbkWWNAG3vOD9t466BNjB/7Okil7ZFKm3UKtIiSywnCgTg
XoXrKwBAsVYpcr5bQFrvfb4yuW+IBdRcwD1xndQF62NEgxEMr6GYre2KVHce9Jt98Sw1OeMog0BC
SuJoQB365AklHswHwdO4Ef/e+Cg7GzVNpC79p8dOTn0DdMEXcVgQzYdJvFPyFnevbwj+Zin46A9z
a9SFU7iKE4QqcBnBBxqWpGOXD3z+nubqhXKu0I1xBc5VvQMK6dUYj6F/T2Xx4udWPRG4bZzArB7A
IFmJeQxqRViWD3LiGYGqi0TfuoDE7vH8pb1gRGeQlScPqZsnp+ep0FX9Zb1hwdjSXGJo1OmyKYI7
Na3pmg0H2XwFXrSGrKwEV7KAMDEilLJxURfk8KV4qMfFuBhUiEIYnP3FsR4C2PURixHpBW/tSsTA
bf1ohgk7J/TbQgaMvMATNcqkkPxYlf8jVi2YWjdPVsb7rwHFZr157i0JdjN/I+Of7z88o61AHQ9h
SXBb7m433AOvqPYTpjzLN0RwWugZSFanUj56ngtrx3eoWZUkzqb5zh8lD+zy0/g89J2Ac7OSpgy3
FTsZaz4W8y627JMKoErz4t0DHIkAQ3RufWmSdukb4lDaOhvHUoOi8KC9VYw+elwsUcXoB5zP7fOA
3gOFCrOT4LFQexwKqrS2HneibEmBoVTzCushWxmJuLWYXTeW8m1Ki25jAr+50eR57CyDbsS1XoIN
00qljiPqhQJE9LEklglquBhX0H08jDE5vHfuUfbREOJIBVTgBey5FNR/dPTHd76g0oRK/471e/A/
Xouwkq8AyHwVpZRqCZOWdkgKn1z+PBw4Rcm0Osg+ClKnQzkQ55iMndD9k2Vv5KU9Rj5zFDrUJjqi
3KW61MrMogebynXMGokYktd2nT7vUtirbi6lEF3oOGAcqSw63Pdw9T+iTp6J/Bb0FHa5Nw4gPNWe
/ICri7QxUb96vqxyg+uNg/Ha154milVJAqDDQ+NbMBZIlGf14sbr7za8PSCEjjx0urFjXmQduGov
V/OSvgsEIAVS7lIQSlsgRhlrsqN0iRYjinr/fkn+X4dSW6BxDsB1Wb3j6kFHTa/U1qNMZmwtJ9Mh
XKYzDLl/UNzwdQm/undY6UjmCdxP8dgClaW5QZyUXidYzNxb9+g/CfA1G9l8RHHLkU8/K+oelwRu
V8qu9RiipGiEWm4HCv9A7E8D9vknXpSyRyS2+U09nkHuHAojVZ3tLU4S6FndNwhYC9SBQ3LiOZb3
8qBCVjry8Hh9zhzcf4+Vt8z2s3iYdTsvqxehib+oaRjIeSkfzNTEgVPbpdlhq27TzmacHIYwSnCz
yE1V6Umvv8G+skIKB2k+I5Fm5s+TAKXsayZzuAA6r8Ua6v3kS9ktZIk1HZviXXjEf29KzDjP44l/
wSh8LKLgM9CdmzI/56qZi0lXR+vblk/UXqwGZLyqs6OSplFQF+qAgSYXIScox+cg1A2J3i6mYiLU
MbIybYfeflwiNXawGCYkHJk/SpxmupsxS4YDyMP0n0JCojR0U9R1bkGoVF54A/oGnF5//auXs75P
wPCX9HpqWDquUzglnD+TD1uuhi3YzXrpmtTWLXhn80ELxRIXPwPGSRIUtID7zpOTvNKnWNQFT/de
Pcc5oTmr2J0RpBRbs80rqYolbbwj6p8iig9jGTDTJEBXM3qZVwoOzgmUiZIu4DmfT316CK1ELfjX
oEtaAVHx60v+g/YVWgw1xS9iwQAg6zwgN7uuLWrlRnbDCtYhLPIEgv6P+3slEsJsv6KFmgCRKusO
AHG/B1UZXBIszFmnF3SG+9I8IJRlqgvE107ryUeHSCeV0wckqFvFNEe/2yCr1tyc+btcU323Bbqa
/TdSFowD5Cz7KnPkLg5JfVdXgM3t4LlL3EVGIWLpVPIpP+puaUnY6EkQ0QIWQzCfG9w6Nt/BlZZa
9tp58alYHlMy38jxtZf5q2BymE0QZss1f5DYJppu9tzGEjBdCtCcs/Jn8BqNjq5kzCSqOqCRWLtm
4HrPbI9J0ZLjdVDivCGzULmltL4ZVMBETjAzK+9tKOUee+S1M1WXo88vEdcjd123TBzrvdaYccvH
QPMmhRiyEFZXZnyQVKW/xRlQjfDDm/46mDu1/av7OaGnMq9QHES6r/TG1AoCfTkkZIuJb8atbGg2
T83prKWwEvrycorxlEd208+M5RCdOShh2Bj5onX7oY64lv+23ri+v0JysVsXU205IP385Rb1JC/o
BC3Ci45xWzOoQ/M2YopNtqlnQFKrMtuIld2Ow4NcBdmJOPt+gl20yfCPtcTRzaL7mUNSNKYcBtEN
7iP/aj9ttbZh29zxqbrr5c/T+iO+7e+dTiE99827Sut4EVXOeB8THuZRTJoIpAh6OuhFwCqS332q
6ZY2ldug+dd8DUkyw7sCK4jZkA6qApsn0R86KZf4fkrCSt0kzTljh1HKk+C57AFaw/z6aBTpRuub
rXJKl1SfLRJ3KDJISBkR+cc5KTTJ3kyzks1rQJqqVzbRF7eDIRPLFaNEwU8XSVrQJ3Ga7eaCkLmV
2VV/aKeHh9agO0CRAFAqBd4MZTWfs7paWZNhyJb66RpUm6O0yJcxz0rpaJOMi+jj6m0CJws8HqMQ
9MQeLLIwX1+KnfVpPq/2//ihD3CQyNCRxs6Ue+xmCyZimzeujgKhqeVIWF82FBeSNo1HijTxqHyi
GwNwJiOqjDjcDrFSQ4VdN84gUj8P2xL6WrCpaGxbcFNZ/qE/9ZDva5jRW2t+7LwiPAm07h6Ws/n9
gLAzGqUSaq4fKoMobdlja883JXd3/YKVbQ18S14mPsQq2XLdx75DvlXX9AF+3rVOSIzScHnGGaOo
D/E5OV9C2fYojp/G+BXlBicfV31IHtz0+l9rpdkq1S4nIBd4mQFDHjUIqAbZGttx1RHCJnPYOWUI
jHGwpg1uriWIOauWP1bQclgzv+1CjJl2Cyb75lu4Omu9/EEm+nCHmDf4ovcX6rav+U9BrMXpPTjX
ciMAtaBMdVUfb7hCei7z0+YvKq9BLYMqoFXocjyweU5rSGfynr4obS2XnJhkDKcI+Cr/T/B9roSF
jvdBxln8mZ8m6senCDDrnXIMDQoQRv46N8guPVMSj0qekHs95R2oy4o3YtkOPo3tHl1HEINvJPeR
PVSco2Wf+X8kpW6SyL65XSFa+3lGCE8hmwB4qmj7SJWzmY7k6qNlRtFkMYGd2uPaRuq1cZTKtRXo
VykGeNbekA1HrPgga+Ri2O3ETyPGR6G6Pfw4xsS4IdAQ4+yVd5XRS7oPGoFD2faqUdEmufZiUX/+
RL08ufdnxZLkyxHFeagSm5RpjZ7YWtuVc3sceVYSqd54vDif6ttI55UgOAf3Tr8QUdmU64lbVtLA
0Tjps14N4zyiOIIJDOOGIsy+uXMnCMTViuuUuyHSmOZ3eMfZODhMuar8/eQi2lTglVFA25pPbXZJ
TfR8QMrv6a1yXJzNIjyRHpLyFK8Dh33nDrOZfVcE4jvW1HJUmApIdi4LVFKPY1wsa0hPs2Y2CrQA
28u6woJ8/drDbk3Q9aEsX8sH97lnbVPwafjiB2sakzKeyqMVLaFjLYMQAZBPTe9vi8sBJfAnVNko
T3NnyytYu8iPVnlN0YOstr1Xwdis9wS5TxzMlllqtvqjmgXQbOwgdRsIzW2nvHGrF+kr+1fWnCGV
eZc4fbPiy5SV3ayLTRStpuW4stHNPv00tBU/FM3q/B2LlgB0sFq7cOUp96saNr3UxRJthsuh9a5H
0tKNKtrV1pvgjBHXECvq77176i+uVveKk7JM0ol7PPVcMnXhip2XEKQeZU/wbHDdNLkuoKGxB6az
Su7ZmcZDTyyNWI6pWwRQHI5awhxm3l7fBmBzHL5QxDpYmpPGL9wTSvlNa2tblEp6zY+GAkhsCYQV
n3cL690k0JyF+jBXO0FypZCMha+SOW6kF0Z+Jw2jZdVftdHit9tzn3O5v7/8nHZKFQ2hTqAftwgP
8lVqbFPCrydQPmoLibDGDuvsAhM10bR8E0ElWtTcI+htpSQmMzP+E4cgg7mVwxFtlv5+2fJQVMFo
Xj5B472oPIZ1q2hXNkWMU4KvJJjuA545Lk/DZNy6PWC4KxozZkoaK9x815im/Xdf1FYpbajyCHq3
0MYPRgCus6ToXFkGZXlrPK/3xUy56OC5w6qzPk7zAXb6U3bKYf4sZUe/AyZhBa4zfoMWMUAcYWs8
np6nxVCp3Uh8BuWS6+mrpvgQdkM7VA2Z0bLxG8l+EHQPpfyB//BJrMJGklvdiUVkLKWM28CqAN0B
sqdaSdTqcfFGqGIgPcshXkmVBqLEb/4ES+o0TRZi4bkOZLGH49MiR4+u0uaQTmA8wKCoWbPQCzu2
T6yhaEasaCMsW1GVMpMyFoC4huUE8WTolKqge+lYOqAlqzNRAG3/xvSzgaOIUdCn1NZn1RPrczTc
jDU4kxLxRWvb3vBspif6tqVDck4YR/8nKwEzyqNJT1D2hYYO09J4NOCVQXgoPKCJs16okD3/0pXz
VYABX9UoK2VE9sR1VSH5X2oPjQVJS7bTWCR15hjJITWy1qPLidmju0eZK8XOMhYyVO846uES7Wdq
nW187/CXGjFO4istSo24NqZ4YTvieyqYCf10ptENRsGk1t+lx8HTL9dIII+4qepCQuQxoUCLdpqL
konA8TDZFz2lqFLumA1rawHk/U0U78iKL5l5wAZUo6FBwx6nEWixzxH3fwFSk9fuFkNZ9zKK+a8j
9/ccLIcCM5RoRKePvV/jVxxIewNZCQbEvztKTmaLAsYhMBwamG7ZZqUVUEqQcIcV1206IRWgaplW
jDdwvVzUxWXTWYMN7S1bUmQcD3i2wTMJ2t74Owtxmu7/EiGWtfkDoB7bj7FrbMRjRZsr9Yemc7Cf
xb+jLYWhaObKYr+5CO5HPR4um/hoB0ZtpiJrU0oampjWEC7nt9V6ECpZrxUtLnVO2Gr1eE14TsCw
LJyTfVIT0rWvhHj1qsmrLcfSdygjPKj7mOeHqyAMXpr2hRE3XtVQJS1OPLJtPdqgivMcMG0soHED
siz2a2v+A4+IdGnlTa4x/sjOfZTCsiN9UcP6eCQwEQh/MXgPZWnn4zdG7rFFJMEFRsAhCJeOY0BD
bZlL21ptQdcld+U5cmOhZNk+BpLp0w6AfzHy25CsFh6KhPlnWSXXNk4zG48WcZG0kJcxPtzS74qD
SBCQdNJLFd3FEN2OM9EsCDLMZwrNrmVM89NuL5nVbq3qbaW+Q4QKSszUonoF70MD6tPbN7jVjn7p
mFgNvcwZSTCYthxPekvCvLTWLMdD9NLSmgfHP65omEQ+O9iaAA99K2KM6j5eBIrzx9ohEkSkk761
I78mfZiFbWerpRQIPJkNxW/HJD77p957/M+WWbJL+xHzGZQ7qfqpbnheGWQj2W+ur9WwEQCW8Qoo
EbFyaPSoaTuwTvX9xAKR/ZKV+dLRkUsCK3AOCVpOQwS0z0PxfM/ymrrRKcHnlyo+0xDzilYVqmVN
Cu9ZuMcgINwmzVh9M92xanmpPK1PmG5TCtABldInlQqVp7rEBL3lP5fUHBkPh8J//q0FD++0Dp0A
3XSUcC93p4Fg0A3Yx6yUQ0QE+Tx7c2jTwGUDze4B1FZDtnWyYuuoslwW7b/mklZHhEd4YooiEi8a
gIyfIov4Zzm4z4CVmjC0h3YMkFB1TqHefm6QnTHSHCfD8SSpUM2Tl3mZlNrcqfYauMzO117BhfOO
aVsNzUQyr3RbZKJXwoJqgU4w927vTaEPwfjHdD6ZqPsYzqyaY18CZGkSKHzxDmcTG+Mr6B0Ps6m9
SDkBdawjeX4kKYp4GflFobYERkFRlwMS2Cm4Z5yan5a0D4hwjAiZxTLrNYFki/nAKff5OR16kSBj
vt9LWCAs+TNa9SUAr5Jvt9895aKxi811+fhouzRhEIoWx+M/7GWoJOxuNS0WIfJBpJtr9EDUcTUF
7R9hBvxbGaJMXtbVsN+aNGCBsyo90TF2YW+SXMB8kmRYhsDDUGWeBd2C5ymZMFgxEszT+GbW8dxE
dVld1nMc4VhQ6gUouYhtvTtnD7mjb0RXGxZcjY5f2yrj38PNV5nyI235mv+Su0wL0/C4s52UQRIz
Oy8fE1X/yRMcbWtq3NVjcZZo3mONIkkdmdVFsyfhLv8bQdAuuCpD6ZI1plZFpXYz0NHfJnBipbv6
nXXxk5Czp9T9uBX5enpBEXFIziNaDOV8JtWRzZ9V+VSJVB1khImu1FhOtHXo08imW9ODXAN1HNmn
m/b6/KLaT4jy2u0cDRwZEXIXLOLSZz2KeixQbIeoUXuJk2TLvo9VYo3mUC1Qi0Go2a7o5qhxYf5r
HF0DcgdartKFInepanYUfzmsUpF1PKPGmOdIxBaxUWxw6XmaJDCiZpYg3uA1aoEXUW1149uB1jS2
LTEM87PA1CG/tqcrVf2h1p+xkDbiKmIpAx3sFfJeFrATe5Pabog5sHjis7fwh37odFJ5tE5g9l/i
lPS2pCmOlV2HHpNO2wOv3BPS6NqAgMLMZKyUt9ajkWPqxI3SNl+vlC96QqAtMeKLBSFxLgOuM6Y3
kNOvwhMtdubUrfB1Vqd4M0bVrPhVgiavb4Qo3kbwslXze5bIRaV76bXjx9l89VF/ENhYiNKAvwny
FTSFAKFQ5t6DDhIxHe0azQsCGG9mSC4SFK1LzTstWSW+3+mP6eZRs3fDKe8U5BqlJLAdOiEze2tW
Ec6XfdCrcgbmcGKa/mbJiwSBK+y2OA9/GUbqWbBY5FwWWnpDvybAgVq9Rb026c2L/PpRQlgvKtf6
fohmvKzBdZblxS2XKQj7P7RKHiyyNkl5d3KAfkKdnLtH0WnJnmUoaZvBADzvzUTYrOTUQJLob9K0
smEAEN/xRx2kt9NQy+GYLfGE75PO9YkgB/B3pBryLs1FbojjnUJxVxZ2W1sPx6fVpCdptgp0ZfJF
UjYjZbv8cs6NfSxaOMBBvAW9DCcA+ssup5jdXgUxKA7y7dePqhS/8RlAuNIgUP/lZg03JGStCZkm
3LUkq8zGFddGd+h9y7qcI94AvT8hV3FncVGX/XpedZOLydvLD1bFhlqMyoNflikQWTbzEcZXFv0G
Y2bTx1E7eWM95g8/irscWxLsj0cbMm/omPShfbVtKd7ib/yMPnwFiZYoUb6FjbXCjQJRg6hMtHGY
omhey608NJY6ArwisIYNdi+saI+3ZH8q/uDnuxG2XUjq/0ggoQcYke2rvqjVE4yc3/d8VzEfJE1p
0nOxB7GX96sVMaiUBlM3bNePBnZvnOKF4oQrVlXuund9Fz/oyIoe5rAgEGqO/P+j785C+/vXcqHh
wfDkqVQK56+8gA6UNXrFb1g3F4HysG4nhHYd157Vt/Pdy66WqhDCqJ+F+TpdwnXstI+U+AX24Uoq
SLYoHSA7Lcyno2g56Ir75B/K0g1Q9rlt0WTGElACYOPDTXAfb0UL8r+jwIO3qZmcKInsk2AP59Ci
wfEo56hCiS+9kl4s5UqVvxjitqJ6R46rIISjg8Z0UVzo+QIJqUkCaCCiR55iiSF5ThF2mdJ+6DgA
x8ufoKyz7g4ffagdShFk6H+qFOiJ53AoT5bb6iBpDrobiMuydx4PhNv1ClxD4OH8TSvAwGOUOJeB
fzrFbVXlpVVNgCjKNp+v+dW6hV1reyqqQuMlV08Z70myvperLrbx4sgKpkeLlGucGtT7idkVxWXj
YHBxxEmxFRhFNGaWX25oOwybjgij7ryXnnftOrAzK4yjTpTKdhsjL4iJoTxPhLxGS9tuYP1quhpv
6iByTk8ZuFenXvCIj0RqTJV+Slqp+qFvwVOnmHvytc0lnIjnZ5xjHEqt4rbMxUfM0EowYCsEZa5G
dd6+1C5bWiMiXFvJ6qgEkLK5fqlRx+WQcEkJWuFjLLcdUImXKdvsEcOLZ9q/k8WAivIcIu+44Fef
7nZSel4tWxr54bbUtL4q6IGm40YgMlYvsf2Z1JT3ByXWm0njWWMvJLpkZc329dpjpWwaR9BvtKUT
A/9vbWseTIUAEkZrT7qiMTq0G1QXjdv4vfO50+/rW6yqFjWH72URA4R68sgOV2Ld6s6PscVTe8nX
whfF7ZOnxSQv+X4+HL11HhKMssavzmmBdOl6LptDMIcaeqZzdZHPSU83bGH+ss4E7SvUOhpQF0jz
/z4g8RSfZlXRWEiVxKT5Pt+6ebc2fVBjc/HM5cqlPwkDPrKly2KLHUxr2rOJbVtWh6ICdRKawedZ
WJ/3xwP9XhHCLNcrJo9hzZKOtsUwXnazc5gKM70GqD5FCWw9hu8TsDZm9ZXBzqgQchfLrqzcUukB
KY2xYMCmgPmWVVdDgXCygTRm3fsmyalpBh3MaD0OfuUhMjgzIbpAu5LRJFnn7T3rVknuX+N6jzV4
H8XKHx39US67+xg83XMkCEfO3YxrVtsySOsMr+XSETnF1ZdiuPZvs0pqVRSri2wpRTGZFNbBlV2U
oBFjnxHRUVHTEp7yCDKVHDidrkA23MDHMLCE0o24IjMcaeyiwQkOPsmu0ZGqO33SS3fPKBA7vbhu
sxOiKxeRQWx5CwIoj8HfQggtC5H+A6/2/Gg7FJY6kh+KC3TY2amMYBwYZPA/2PAx4QcOm8etQH+e
/jTqOJEbxNRGVVYuYSM01Nt2olSfytS5DA6YwoknPflohs/bfIkWlMRC+t7SAJQwBQc+XoNCUvDs
EvINET8msr0qRIWVUBHWpg0nPwlJR0ogkOXQZ8jahUkkrEoJk7D+mntzrz6HQnO1BHr06U2n8wjd
LL+Ap7qGtKIm3RLaXH0ihFq0Qw21Xuphviw9AnK8DWDaMqjoR0I8Fp+hA9/AW6g2NDmJlclBJymI
qkoWM9BSu3VAnb4WW/f1Ua97sBjP8JipeiBXMXPvzdZL7jkWToYI7q7EnlC+tlCjK/Xxy/9O1Mr5
cN7GXUnBnVl083tP2LSi6n3i3VBjPmo07iLCGwG1PzFlLd7nyV+GZjLTpHomKUAMF6OxCaYYiYNO
jaKlmIRWMauIjTRJY/pmOybNfCmQ2ag16SCc6Vnt+LRzMHboU85/ijvLQ5s4POgXClKRDEepmgwi
fiy5PO9skMJwPm8MuuaW13pIb/QQ57UuBIuQCGfFh6hWSWKt/OuhSHlaAIB07LEbYdBGouFHONuw
4GyIB+ekx5g1zaG3bfWrLjDp0spCLpyJBAuEuIBnG76FGF2m/6jU3gHmf/C2TXrIi0yPdnFjyZRh
KqwOHdwN6ZTMZmHo5nWUYbQSqSimquCqadwwgDPk9RIs7TEsxwwMGIPJDe8+vA2eXIsfXd/T6fM5
iDlNz/D225T4Q1AZ5M4tEleNXYt4B6dvzOxxTCEZmax40wHF7Jghyl3QhS7ES5RqT0gOtzQIpcaI
6rFB5IVDo+uJGhP8dx7zybROEj7Ny6g3i32GOLsl51lLQz/LoMTES5o7kz/BtpFgi7AUTN5ioH0N
TeudmNTkqSRe3C7SYf2ptdssKmHfmSDlnj4vYbg01Gt/kWyx6vqRasN9Tu9147jfqEtDXY9Wkfog
Eb/8hnNnw8UY7hIbHXVNc/LmPklzBvfmNBm35iQ+kWumtO7ab9PgcTTLPC55Y8YBGVpLXF1+YZt9
PcgtGqQCLtNVB8QXaDVOQCLULry3rO78WeTtS/ZpBV4hgWV7u1UOFOSbsja4FkIM3haS3abB3CBc
SzzZTGQ1dEBytlQyfZuDf2yeL2nJAjEKHKz2R4xnPpEAMoX53XDONT0VfwlRll9tz0ftJSFRzhET
ojjsvP5DNFeG1Alvubp4NXjUQ2F4RezdeuL6duHbok7Ok2Pzeg5kTHiJNC7u87PTR8rvHIs1QVmk
FMXQHKGoU7Y+6ddWu1i8MqZRXMEzUp+/BL+mnMtzLzekwYOo2Y5EJcat/cRUyOlxzjy21u91C3af
GQN4PbZ+AZkhmz/+6tKUPbc0zC+Bl9iD3N8gAS907kOcHgJyealOel/e10nts2SYPcYgsFntPcUH
YwA0Nxcp0EkRSiG7M88V3ufdOaxhvNf0hrPzlZlN4WfuhYd9dokIdAhLPB3TIlWL91V4sRpKGaXa
ST0S3mnJ/vYDT3SdtvTJYceI4/wENW+pepNQzKWeyr3R9Z7AZuGqU065ZtwqEPxBLiP+EEIYltKP
KVw9XxDqXhXw3adxG5emQAKd/deqG0ZMR6eLhSbFM3aMXLpW83sFgYcbQYaVsjUatede0T5AolJx
2wAgjvBIORK/U0NlVqCyMBWVQqJldtCCXygzyapAnEnJn6B4HJDcoXvPG7CMfkfCOwFaZZRP6j9E
H+DDfWvZtvlSqOkFPTBvZUO7UdbfLzhFgcj0OKqAQglCtz1fp7JJqtNQ3dI9kHT6artMFalv0N1d
uaodruIJp29FgOy4aw+BDRxwOLA/9r1EGUeE718QX9Rkh1+RxKx9v1nWD/OPBpwCt6A1+a0Vz1fU
oaxlDUVuMNiVDorngoIqsS9Uzr701tcVXEwq7qt/A/16CWfb3Fkhq8zvsggf81WkR87KvthW2tqn
QCBRiR1aa8P0evsq4ykA/5HHoxclf9oI2g6nfmvovKMI+r1ZkdAryu6iYHSVUnLGyjhai/eWEy9j
/A5M+OVhAWhkGzXCV1svOizWAX6F/WpUqPjUEpsGo05IL3H4zf6n6iWdyfj+Zazcz0RfAIMiqXSV
XCPDuAzw4D+7U7kh2UKOzQQeYJP5/eLNtInLS3jw/IZ4SMara3AOkQ+Z4FtbWC50lBccw5sdajf1
CZPT5obCTBT1yTeoVElOM7cGr1nbWwLl2XDEhr+wodacEhJARQfKhc878lQM69lsZSNnELpHdvVI
veQamI+pv22fTwB1LJkfAvOBn+9DtFyYij94isT09imAIQOHFoFIVSXhnHV31+OPRnltOd9VBFS3
wg98FKX+tkhX87e7/fwg66nEqhMcmG6kxW5fg/wRmu5gx9Mr8YL27m0maXB4iTvVqS5nFRF9vhdg
E4OoCCEUjFvamW8ISlWC7aGRWTDPqwz41QYPdjx1zDKVl5OoM05WEkHpI8qfdQpb3pbwqX3s+Vsa
ni3uZ8JULmddtxfF40xW793pZ3gXjWZThvJ7zWU4jBNTTqApf5afnzna0kEO5eEeDe5W7OJZay/x
H9odsDxkmA40mSo6GFEdJhUm19jFpu4TqvJRCpJRPfbqPft6NqJaRytYeNyRgfthueI5AdcN7Mbx
XnQ/W/nq5EFqQSj6VMXkW1ifoAXP1DKDk/Qnk61bUWpRMB013TFTRnozUiRRkwMI5aftIVI009Xp
WjD0AYan5z7iqQJd+qA44FUjf4c8wbsitVODcSROLkUhFDOycnY6nqrmGYL9+aomhDCMbmk7gmoZ
TcINkIthtLQi1D+60Fey3LQC6lZLXV0zYAsPSRjlyfu779FEUuzfVQMMN/0A7jxQRu5NWy09QG2U
kA37uR7EtmU5oI3PBhGcirB64RuwGpyYEl27IdysYYj1LwFG3VrQ8qxGv/xbDYgHXNIYxOduMcat
BbGG9xtbMX5XPVgEDn4pAXCk6ogWK9i7xKV45cKXtRtGI0TyvGiuhS9hv20gESVch40h8LMR8tqt
CYIusgl3d6hgNOM+6VilclOv16NU+AXsNie9dd2ml7SMQkbcReLuSkKa71RS4OnWlTi3PgEwbE75
/3mmlGbES8AynX69m+D809hJHkDAqL+cymd74e2rr92cUL2c3L0iXLrvo/IIMX0HVJDnXaBEW9/f
lK0V9rP1lECqquBp6GY1fmNmj6PlgGkfLyTUeDsgXoi3RHsV4GRdhqYGPBJolk6pa4Yx/RxgQaZC
TukjjOJe09i3QbY3fAgTeg3pWMGfPV4YkjGAzUB+TTG5lhD0U3eFCBOmVcjRzCYby1fYJMqOVO8x
f5+nf9TBndjqFwPq7jXuEWUlSCDLvSUJt0bJT2cbG69lV3VqkjDR5ssOOmUXig8TUS7MrphChvgS
sE4IWw497IAZefn7eHmlvKzcX7c5sOzBV6yjOgRfFoA/SpbeqLV7040kIoXbS4s/LJCqE08+N/pT
Ci12UA+BaQqq7DDSrA+cku9nDwiR2Mr755T/+pEz26QFBTBfV7m66xEei3t251eJksyoCnOIdIs8
caW4dxCjWEJODOXs3eviCHdWmk/wlFHIl5AGWF2SgYPBm2a0q0FPMzVfiKliPvKuVoByp4oDX1/N
Rys4GaZOpRCfODovqqJ17kfyWEbIPkZdBJePjZp7FzRM/Vo3sLNV1IKwScOhcesSyNNTUUToNhT4
IyHUQeOHuyUO1Gbe2wix10CEt+Xlb40FBuka81VhlVGpB8/xwHxAHq4ob/iWiokzTe5wUiSliKC9
Rbdyr5MnQWtbvdhYFz23QaZaUBHmHcKfjRmq0lzBHf6UQ+olq/r7NN6e2EdSUyZDSWh0NYPlwOC5
1RKa0wNic6CSlOdyWrVDm//Z3UQZA4/FyqtoVffUIFBaOMRqpgP1d1gPbB55pI9GxKu4YOdX7go4
WcDBchfjLMSTjdf7tuOtKyDi++KsD0LzqMtj8CUZWAewaO53It5uZsqT6PEMKuVn/xwLGMk40RPd
SzE6rga+9gWPWm2NAb/lfW5h4P1zPDb6tFsz9MHwWxeS3PcIVA2MgOQsSPVZaWS2pvXSBp82ucJD
rDDlk0Ayr/ucBgaEMyM0XiQUJQw676phR7EPR7nNE7MDJd3/QJQMZ25OWEw9Ah4aOivbBOTMGAw7
f0K9aM0yGDHdh2joEB266mF9NNUIDEipXqdX2huUnGMoPl0yJ5D2G8X0gN1y4k2FWH3JhAx4feD+
CXREl43ngXQCIWh2eF1axqkJyAsAs22Hu48rWI0htFkdRFxr5wSEodJ8Y9GqHq5kTO0z0ELhLBkC
AomcdaT9ilznsI0yRFNGqVAgwn8oY1c7A1+4scdakHKa1efKy0nIQItB9rFgKMUSX/qYDQzyR1uv
5JpnGRJmV6HBhePC44mIIZbOe09R1uVrkWA8mLRr3l+BrPC757K7/z54OFem/agJVfNDHgRgQNau
PkV040IrjL11XFLDhIGsioawIbwrcttaj94+sxDw+RqUu5yUgwp0di9evdNJdicPbD4pSyhLOxiz
e/cwVICMu3ui7Srj9SWzW1BxO899F5mkLv4s0sthyG4tyswxSvvTnG7EVb1JHYVcGSNxFF3LoCiY
v60zZXTi3F9qVI+yAJ/NNitkVAW3qfE2GiDETN62eTWWDpaOHZdDcFkP2xly4+C93pCIT7xWfcha
76pwflevwkDiuqWYZxqTR+lgLbWQTOdTALZ+Bk+RzCzRmbD9Zt9xHDdNnB2MsUoo0EuBDlVb3FlA
rNbC/FbGxQQ1quN81YFldYeJo/hg3+eGHGio2om6IZcoGtg0VVDwjWB8v9TvLtrPxMhvsl8Qw10j
v7gqTMtgGpaqoQmwy6u/QdWNe84upZjK36o1LzDtvv6pxLiww5h2xjKiEMXYNAsSMIjhiYHSDdJf
VpZqrYKMMwjccqkBV9ffrhVmFj1lNwvLYxKWZ4veJnVYpGb7phkYTvKkkdlVW/rq35IiH/7j1fox
zH8W9LGM/a3sv90jQgyECJTNjj9ij+nOvJcFuM+Vi1YdINGcK6DXBRFKT4w0JkfiNu8qGjdugoju
kWMfaSl7WZpnMlD8SimoUEWLGsNoMTFteb30+cH2tFQKDYyBSrGl38ykwHowNpkRHSAUmPkG7uiW
A227t4qgdeheDt6QSknsw9o+k9Qts/CYSBzpEQ18EcmuFBlxpcsAXISayh6dQ8Ta7mnPoNedqvoI
IWQ1327TRUdz5ehpShgA8/gXZKFoJjW17aYOGGMZIZmlM6snNvmOU3BeYb5HTNOGFMS8F2TG0Lt8
HPmgVPfrTCdwHW3wnMrg5Xwa5LhNvxH5kwNKArKpN3PCg8JzrDniITvPI9TWGZyU6wMU9pomwtu3
B4z4h6c+kB7QpL+Mm3n8SLora0IDVBoAxV5IcP42yQ8vkUTcC0k0Wkk9O0lUSLZ9COUvjVOWHtMB
6trocvF3/mm5/chQGqlHAwLw02cCB7YFbygXVbujdtbc9pzK4apFlxtEUeLt9dJ3i6R+s6a3alyu
gajW7CrOtVNFdLuWx/eiOBWN3pRoYzMf3JDMKd84a95Gd9I3TJ3yxuQVc5EUexFLgW80xmU9Skea
7grhzlZahFSRR6o4jx89g39WKRvDqaXwvOLIumYYBGBw05O1m2KOAB1bVZx50o5idcU83ry4ePVm
lPuO/CnukIbVYFydnvMybfl6r57tbb15IU2SaPVmq2PqkPb9W9QckYJ79en++Y1js5WwhMxMDk0C
2S5+WiNOB3vjBh2yOt0lGOPwTRbmeJgt5VSdE32SbuOo2YxAbO3jpzjz89dNbO5Sc0qLDYcwEZHW
Qsqj8qLDOy04JncreTK8GOUUh22zk+HrvimrGngij2iaWMSiySG7dH/E5lV4MNr1LPthlLwsshrb
ls7dTeEX5QsxiQf2GvaDQMWpYX2vY/AZ/2cOT11wzRDcNwDOJx5YRJxfN+aXzUZE4kzUVA6tGVR5
9evwncWI0w4NNI/aJs1lIoeSMwLqCu6tyItK3E5iVbvCEuIQQo+tLjX5OMnIMYPrHTFSExn5rdLU
jxveXTtlbgsL2Yq1Q16rYxZ1klw1mvMGWdTOzd7E2CZ9bQWT8uTQmqlBLDaazLrL16WTfoQRixo9
bRuHt/0sPbaM1GSsB5Fa/SfD6R+/l3IjN8mBgyN14JAI0n3NZ4DgjBCW3ZiyekD8hK/klxd8KlpG
IqWY1TtT9DXOTm14cQZfRm3HwIvmrr6op7NVigCzIKuchQ7HzXYpAIcriEcJi1y8m60sNcpTa7XV
XYrqIaJExvOcTb6JFb7kBwawQb7CMENwVluM5dRbTow+nsRdt7xBrhOJ3hGatGGU7TAFmapMWYh3
VYuMPDo1PDZEjiuxUT8YSoHkRSF6qNWilWo5JpUulV9mM38OpszE92MuouIbMzncK08O2gqLVoR3
Twjgk2CuwItys73qL95R2aSZbvwbvUU/et5GI4QGiinCDnJSTlixEt9llscCdhvwFIgWKWMsJKN+
uOBwwSYVFdcDHnc95g4nwWQtufjraas2A9e0dYLBrISYddmllwzP4w6hT/kszbXNpoAio/jA/FhR
0wBqHtbBWWz0HS04HOmaCQklHAfxJUNHLFcK4DasgXpop2mSYurq7OM0N2dGE5Nx5aQ6uo1qHtMe
Jk2H9rJnuz5TfBjNUJp4aNlIWV3CyrpLw6gmPWKl+CqgssMG5wx9e++jD5aH9MqddF1/17ubK5Pf
m1TdPcvcNusXgfpdvL6WseuBeSqgbDRMrPql6pnJo+f9AK+koM+mohNFDsvmH9TMRDqPbIGUOSRA
PJQNkkcBwP/6/15gU+66LR4zOOFHAz3VLQlxNwKIcYc4ymBXQYxcYhAtWZeVXYgoT7Plu2KA/irI
nk+T8jr4rEegFlbmEmjuml2bWccodyGvU3u5QeIgBpqIxENCsAWyJHRcQ3IIqTDz6LqrAtIzTH+5
vgnTgXZk3T0HTjD30dkoeFsnPxgOI3beCf8msIscjeDlhs+mrqLVPNEnUtCWD3rE/Q7li8XlJzjf
gI2XVOGlxzwx6ELdU0/vkmW0ZNzui6RCG6xZLE/LJfjFQuaymxrkOu3pH3KHHuQhqmaOJYFrh9Ng
qtGVqJC8C8jqTa1r6e3RwUfzkkkR29GS19WGC2bQo98u2+hoofAHNXJ/DeEh1XofsIywpaa9HFW7
J2xxMVRfr1GKIbXF6HfUJNMEvUtKM/ne1/ArDqh+2cuI+hCPMbCK/3+Qrzohr/OlCCi+1Rwmp5ND
gTxYtywl6CVD/CM9KNQnE7NmWX2am1UzkubC7gNZMMQpKyyNRjL3RYu/bzLDD8QakmW/fMppBpI7
17I3DvqxqQo73jGbcdhfhIyszloXy1Fd5H96LpWB0+oRea2dMaNop2fQZcwE9TgMBScUyx3Yz8tj
TwDCQiSF1Uv9yumhjjCYDaRU+p4eeszrcXWCS44umQ04KcKq9MtVu/AA4mLA7VqNJvkGvYehHr5k
jc13NvFpIjOyjpzmTF/c1PnquNJNduUuRxk/nt4m0KcctBkP116HlDaQ6pAXdWiGrI7V86GEHReO
l5vHd4b8pq1MxWQINZQjSYIEzqQ9hHmE+S+FLHLdySYr4kqoBS+zDNXdOFRgmgOUMlwHXqMf/+yS
gZsKT26f5kZuYse0R0rhZKYI62n86K1auhkeAgFqwp1axPbubbOrocyJ7eLjQ6XGhzBDElQcXZau
95xhs8bWONybRHb8wHfdbyikjBLIstFlsU+zmqoO8xt6sI5v74/UePnsqjADl5R9NpZJNNRN4pNt
GQHemmCSyZx9PHc4LgceNh3t/+1TrTdCvn7+09asWii1ohDaMAZf9KPGdAgyZcUYI0NlQjoSlYpU
Y54bj2VVnhQEQXa3hoyYfbzu6Srvpxk2xKzb3JyGOILbkLTtg+RTmcNBHE1YLKrAkEQqTfdcXjw7
HTBeRSp+sdUUbCtDl+SB+ckq5nxraFMP9Y4Qf4qfY8O3YBrIyvs0i0qDnUD+Fq20/yoym1VtbQ+2
O1A8wYOkYrJNRCnJ9u/2TeF4O/VFWMBelqDQH+YMeUSAwL0Pv6A3z4k1OOtu+fJR4Gf3L4ihaX3d
UPDmOSYkCtU6TPpvBINh+qbe5zafc/PWUldx6cWzP5wuqrMjkxPH/GzNoXz1e6hBgbrDylgZVn7v
J7joEfwxtC/plegLBj7Ft5yLysOtKyjwqtF56u8kCfb8JGllH7qvQlk08FLe05N0S3+lAnjRndON
dLnz3O8HuIsiH7ZTe7Y1jtqAqVSTjbWKXNaVSTuXsb6iaOii2VV85oysDHc8Dui7v+94QNLRvbqr
Y+XJ/2ZNVL4rm+Bh8yjq6D6ArVSF4o9cFiGVSy7ge3slWkrA28GP3CGBUvq1hfhDd9aGGJfv7pw8
AhbVY7r9nvYWkM8KW+fERQVz7+5HI3FCmksIHGASc1D2XgXjV56TtpKjkLno1yg5nsvnr3oqBJOw
Mth9tdlq5AFcFYA6P2167zKN5FqFvnEl8yKzsAKlnLRNSF3RcnGabUGFz4VQ5duJAYtY95dbheMY
lKWVmqp4xSwl5GdEfteV8aD1UnR8scqcIvQYxcvsEOx7vG9AbRLQjdfLz7ufqNmFfXSLXtKAm8ku
E9976UNjlSVci60glU4K7LrZtyN7lMmMRqNVuZzNUY2N2v69n+B72e12L19fo3k3+oOvHnK4uGFc
idNSIj0VimqMPlVrUIX+BN6ZCd6KdKGBmIZ45B30RDXgio7Amb1e/qA5fLqu2pxKQTzKmkSsnUhA
4adQD+Z2WZrWwsFt/PvY3IJIVgUW6yfyKyYbPhDiSt3oxfAzg9EStkqh9mgidk1JJjIEgdPxRxZ7
37JI4vO6KcYUts5VIX6HJzWmGxJ6AH1DSY31c/SZEAvzuCG4hapHV/uV8UKf7cLB6XtLs1TZ4TcF
NBdoUIfYpUgY+6TGNhmsfMaGmyN0Wtn/vYWP9En3s/DUKRobVvEX5kPkjEe4mHo3RI/PD1X7ZYji
E6cxZCPMXOx6ObTUXRER4iKx5NKLjJlXBRYfFV/JUrLASulpG0e0M9gHWmXOLoKFPzEknJ8BarTw
Xu/9gzHnikdZk9uljxz49JUTxRsFZhL6Aos3esXW+67NPNeT2XGLOU62RjNI+hbMuCQ48UUoGqo0
L0VgIFN/UHpT5QPcbXVbYurSA/EgZ3UnvR0iJDYWgYw8/zwXs4HjqzIwPeeWS6NW8qNkQnuWzQqm
oupRvy2nE6UsYlSBoV3yqKGjEbNiqUbXSJ/eJ2TjwI8ukhsrAVi46YSvNv5psPmPMcZFdDZLToe1
x/oEv0dl9ntfTurmb6s6vXyTdws5DmqFMpGMROY/tvxS7HSZeBHCICZMtq63ZW2M8lG4bJwYHcO7
O86qALXT58ixP79DVHYO8gM46JChjzwfiGUahWZphlMJW7E5GUmlaqLUcEYTgNOTvx4mtufAI2j/
hxR2SStEcGP5qOQv+H4sInOygfndMNvJ955xwA6tXiFFBopbsitVsx6Rqva6URn1MVjMwjWdc7n4
ifS79yE83aEv1FFRf897d3pmcfh6VzclugfBZN5E8Q3ThUz7DAsaImZy19vXUXPViKjnYUL2JXYP
Qt3IsJraMSQwSuCicHuvNEtlGpP0W3Uv1vMUPFKUnt1GfG1iT4FvF4owKcTjYGWQaL9bvh6Qfpqg
CAU4pWLw2ML6i3Z6xzCesUHo0jBk401Z6ovZxl1ZNpcMYSYeo1INb0jXQVEWR4VVhJ9EcMaDr8qS
F2Ug+/HZ5jqb8Hce8N0MtJkLllqx+MJWWfVkJeX6fpbM+iobn/8ZZzDzaLgWuMlV+iEgyjG6r8vu
S5OsNDpX8Rn96GNSzhFAO24ZNplkC/6KJrMbswJZ8ggleWJN8IpFc5Mmmax9KuH+8NlqHMvnQRcv
M5WUVU5BULeyhdLqIYvqxC3YvvDJXr6ryNcHLpj0w9RAny2nRVkOFdAf31X6l4RrsVIZKkODAElG
Qfh3tybTbWS6qJXjFV08Jowwum/1yhOxzpJ1fzHGyZEtVM7/L+CtMnycv6a3QukJwk1vPtJQh7fC
KEu+dt3nBDvhkrW3Ruf6siP+2LEPiK1tqa5T/smk7Hn8/IoAm4dCfZ3u3W/ndjTLqARFkf6vfp2U
IufYw/wIDFoCP5S05KVCeTj05HhiewHMXxHdipXQc1gwHGdh/lmrlY+Rhi8bYWLbDLVw44C0k5sN
he/UDJVTpobn4sJ3DHeKMrbirceWueWUP63qRJjCErA3rL+z14deE8051Ynw26GQsbZqymcx67z6
W9r1jTw18ukWT5iPNlE3hmqUT3o3D6kc4zAb+GMTlcsmEEW4QQjwriIF3BxiQ3z4ywwEAiQKH/Xy
SQJJUFXwgHZsE2d4JQSSHaLACkvg9lKZnRukxxPMoqL8UgoIDMrJibjOk/wYjy4GftHHTz4CVtge
u44p9ITq0b6quWkpdNt1HgOPtMApUXwJUm0vSgQMYupMJtODmx0srwo5ypcgYMjEP5/wkW/el3BL
IZeZ2zzqBoWaZvBOY09z0cLrtZToXDxmNG5NxU+iHBB+lNpTSpTHMOR8w+UVCeKEO7WZCN1pJRp5
ItSKexER6wnQd30A9u9DHtq5NC5Ej7joL0TPdXOlMedzWofOlgTjKRuYVxJ2Z7tEPhMmYjHsjhPF
XFo8DGtS8asPaYbxHv3be5l14+57jXlKWqy4DqbaAe9h39uvbllKebTaPaoVHDoPr7cxd0Ogp1/D
cKwO9Lm+wkyDPNtDAX0lJbIBB10wuVG6RwhO/8noOJgv4k/3udMeXzWQHgexiUuxgNp65xb0heWc
r3Vhdf0ArI4fFocVajPHCTAIE41d0TE5Gk5ey0YVJaWsKcTimlCNEWScu6ldgogl7ggtvDRodXb6
cSfnLeLIPELrSzug+tRss/49yWmtA/iK8zEdCBUgYHHwPuVWxSUojWjVQT/0HYyiYJd3pjBx4FdP
p29fEsi0gv2RmTYkQq/NQMnrNaMxkgmT6rK+e3mYEeo8WtrXGUHQhKsMt+/yosxlQgZE4V/oRw5z
FTmy+qhilW/k+pMsOJAPRC46hyqoI/jlRmAXXEgFlv90OqgtXYUFpDfGVXhvNPL2MYkh/zUBXx9l
AMcRIX1B1n55cL646iXVdk8Eo0pYA812ScrVq0JHCHiyGouNkWVXfI6EXu3ke1tGbTj4RWc7bbVg
uqbZD8E03Ef2Kd58hmw8Jy43M+dAFiRfYVdD5NICMscLJsH3F5SU3pKYeZ+3h2HohehTQ274PIK6
V45CVXT9Btj1o6fWTOSUQ93QHe0ilH7thmIWmOrk/neSugOpI5gQOs6O5dTu2WxYu8tiwTpfUBGe
FrqCsjtYzfxUTZy5x/xB7u03B7uCnu2zQ8tQZqyDPzw6eowLUYKORVx/acHhr9N8QQdGZsGt2ZnR
VvVl40/83w9/aIY6tOsjfv4vwGfyHtdXTvwhuxP4WPECg82zK3e5eICZdva5OLIccwsz1sGvEcx1
29G/jJVbVKvmhgGiyt3fAsQXBO/GGLNvyG5HLzvEXmfDqfc9plauwsisfPv168KxIVu2IG1giI4l
EJuRhlA7oT31hZGt64/so/CXg+xTHMxudnKHJKrE6/F9hTzwfZ9kJJqXVBtExf61ieim5uf7+ptn
58Z8+3OG6WWK11NBkcCREPFir3Mqnil7mGDM14ZP6W2t9qTHjL0ai9fNnievOPZmDJYLO44ZAHcs
kH+yvcyt2BWDYhbqBl/rOxp+9G7c3HmpStt/cTt0eGgC7oVtYOerqIRChTeiMJuRLx0uylhaQ7aD
ckJ3ulIUq4Sw8JhLPFchkcoypVrAVcLNwJVIvnmNSfJU2NOs6PdvaQ0Dp8RmXViaATmpufSuE7LQ
cZDNWVPGxtShxuLMZNTtPKka+1Qyh52t9MISBa4KmxJEMh7Fxqhzvn/1QBu+fo7G55yfMb9B1u4N
TJKgD5/PnPigPeU957uJuUUkEJZuJo4z+X1XrCvAMHGkRoTVBZyDOwWYMeLYJnp07fnZjDdlgL2X
d18JLBSAUXCb5flUMDGXz56zQZf09FbZCyDSDiDU6WH83W252XCJWha47T/KxPFi4Kt76dDAQOWx
bbjDAYTUn2vWjUnlBqoU0n+2KrAcBwvS61s8oo2tOIPuBLmL5mTWF+1g+GQK+m/LGWw3ja797lgo
b5luI9lBzwkV8vk9zK+FqrqkgFtQDdmOh37MGnmNbaXfQnY9hb+sHovk/O6oYaNh7SfUBOvSVQ6y
3FCE42LBRjOkAgZn7k9ot+yY4VxNO48D5qfCypd7RxQvNaCyjp/3HPynlsCx1U+T0FWHb0OMrn0S
JKKprTbrVs7qTftIwGNF8SRoET+hsWmfU+Q8Mu9MGAccg8nLCJ8M0CFxIMYABsyTH4cjzu/Pevjg
JZ0bwdtbyXqXsoTUCx9dC9rBoRtaF9QsB/04HMn+G13hzT8yw8B6B48QYhczZNTjubC2BLPX/DzC
0rFpfYnL7IMFASa0Qatep4eqb8CtYeSRUu7LWd2HpnVp3ehvxan1JEKbZ17Anj7GwnT3UjjLokT3
ichuSotgKXKQyoSWoIcfQPCyFAjvtDp0ANEJApmzlNw25ux42HXOwwHjSj5a50kEWU5BzXgaVLN/
ZWwbVS2wB3IVIjXgfENKwKmEnOC7Svu5fnWu3xL9SvzQmSKbBA2lwagsQ0Xd4BLoH17zYbses4sk
HEQVuVLwN1jvvbsCCyv5dWIUh0XRIuvhMwqySKvLXKwUWess/+1h++UN32lQXiB+9KARbgbGuONc
4ls2XwTxIsJeGrqD9rxpbJ1B7OBnS972od8v/Xw63IqD3lFobnmLXHb2ZN1KfDwNFUQuiN3GPXB8
Og9f2+FASamAfvHgpqHbaGqO+i1Ga4Flz1fEefKDrWBRwhTsfIOv093msYIsxfU9aLr8aqd7mYJP
LFN1EuD6bUdnQfwCblC6H/I1quFyO71VRoEqlzewPDw6Q25XYA/siuac3GDywySkBSZ6uw5kiSEV
euqyLZO7/29SdPgsakHzNow6BSMVypj325SSeOfWKL8SzSV/rUI544zSSSNw3wIFjioGfMIkcfr7
YMYt3CW/+2EuzFP8JpblsTzpmputdq2P2cosqv8u1T4ptxqZfGI6cr39jtYTGiz392zp9mcydFxI
MNSG8O9AgR/mq251bMEGVaKSO6cPle5W7ZLRUwVyc6HZtRksJDIxXVEWpchNQ9c8ojvf1PTXDhrg
ObqSO0xWh9MqVl1j9/AWAKZVz5VwNOne7/JlY0/VbBh5YyZ+PQG84F+PpY8APaA6xQ+mWWYuDi6d
euexkVyan8dklTO6vznx6h55uxIdsKCiWoK5DAqc1/kkPK/jNmFUzFAXBhSDXlT5ksdpQ3bkMUxD
waZEJk8OXLbiKaqCRBqRABML13lr4lVd993Kb499HwJBtN/l6z5QTFx8LMRZKqmz7mi+eAJjDYqR
Jc4kgZWzLSlgSfqVRMV+iKGJu1qXiQkTxdznEO0veVAVIWTLK8zlHul0GueOC2B9NLN4FT7JfUwD
jLA5/QwD+OdfHMuLEwPPDxNEhKeCfrnSDX1qJa4qi76uDezPZmKXq0+6jKtMwA9EBiPr7iEm44vG
bx5oWnxn32svUJm8K7KatGm2jreQYSRgDxLlGxuqupZIuzvpG+po4foqlOzxwzTWuIX2w9REMztg
yeA62pif3s7jcyEH1DAUx7binQcofYz+VBW9NnO8T3Dho0P6c2Q3eMfP5ydelB1AZqXubaKXkLwd
xSQe5GEyQ4Q7rE6zff0TviTdCHMdDogDigBB7Lu1T3HFWxLaFfk4luSylOtr37+N494G+5FpyHMx
bhp121awsUlH5/TCQO6WY/pj/7jky0Sm+8SmbVKfxbc2ZvGgMued1gpqXdb74774JZKIMqQhJ++b
5sDKj9G/g8nk4gHGE0+uunekES5n/GVUlydiY88rR8SToriYh9bO4ZH/GtIPL18wDmZl6lTTTJCy
uowi+fptvfCmUtN3pt9a3l8awm2W9IWZXRZLO/gUU+h6ZGFZx3y/+P03WHzGhBxy5mrhRnhS18YE
dVKAd9IJetbRHRvJcLuWi5IM/YRev44lWAI+6HEHx5PkN+G6jF0PyDuRENqXrdmRvv6rBhvMDWCj
/xLC02PjtipTf/8FD3yDvIudFNBZ1hiU9b0a7RTcKXAahny6Yk8EQPdnggfVJ9PhESXTTF6L53U2
uh8MCnNjXzOJJEc9gU9X2FKVFX5hAM8WMUdrobGwzVK8xycDc7Q7p/S0CbXaLVKfdWsIGBmY8mF1
Ed7JgA7nmR3xqVAcC3cNbNZyb528vZGFZEi6dDvd7/zfpxB5YxE2Zr2jjmOjkqglR3VpVvyV7CPE
mmLRHhg4MBi8qDDZN1QpIE7Rm/8GOCDL9K3almQtATnd5yjCEgwlrBC6zHcqcuxEC1yH/nMr4LBi
7gXleAzwyl8i/Kj8pcoLD9yGULepN8AQJqxphm69lVoWoWcFto5JCdQkIMxOGHk4cLsdRaXo5DN/
tppdfoj3Ag1yV3UvhfuQSpfk5YSuspIh9CnQIBJ7rVb+B/qz0OHfaZXUz4eg5og1CaOgfaAuyXdG
poYbvdPawHPxYQLrxQBsRY0Qz+17tTdh/uhtCiJpCMGW+Kww9812YZKzg9GmzLd0/yg8EWvBTenc
zD0mk7zswucVTtNzdQM6NexWAALCX7w1a8OO4T8YJxMJM6a8O51ajV3OBA/yPRkt6Cyt1+jF6/b1
SaIza2cwVqnKfNS497ydzSyn1ZHkWUcBD2bz+OWnzyZhNssAWuM66P+bEOmS6h3RVqZ2+B9i2oD7
GzAkSXIuVKCL6Jo6BiyLzbDfLygCUtakkMmPoClkaqk0iFc7O9o9s3yztGvvlwfDCplrkg/LQcfB
u87tOl7bsc8ODhpEeQ6UdYz1ShT1FdruIn84j1A4BAMdcP3bPQDnETmNGI7HX87K6Dwsu6+mzc1D
irbk7LvFkFjNrW1KgXR/H1QEvC01r4zlN+Q6wOlwtVlVmc+fmzm/ZeyeDfgp20z+AjDAUBLe/+aX
nmzqbBC/yUX1HsJ5hlyDwwHcmvmcMFkTx5Dit80AiDY3NmWPkKulxEan865vZWJVRBGH4xJXx1DJ
K0PDCmyKdiyaY/RcVz3sB3rXOK4eTp0qd6VATBnS/lufb/g7m2oIbO1iVdSMo+webLiAgkORRYIY
W3/it2joMr5DpU3feFj2eNEhCJZ4sjfXhGCpAOOREUkkhPXU8UZIO1WWckSX9+2WmRRQzpgC45tI
BSoF3wTp/mZ8FLc2UWRKHcfi6itxu3erb8wfBnsBcHeY7XFxvqQUG8QKYIHQhCNUe4AZ7P4bisf+
NABX0bRevJe7qnzFgBbDl+H8l00JPutFBVY/hQ+L0hWiFM64YsDdgyVO/hcbNFByBFWXMBHFhJW7
RTU1rKAIIsFBVW1WY38/suhGiEZOgassQbI9gPmPCQeMEyUlGt2J+BjJOiPQ7xlZG9OtYFv2IZ/D
jl8I+h5iPrd26KDc3J49tSOqml1Ch2cm1/I57kLwh8nuqaNXzYgSRmijZMH775WyJW2jjTJfGIUT
PMHHuYOtJJ9YV0n86s6PKBZ9bu+X3YV4HCzfnmebjtBCEEAQDOLOci3H7MvsC4YZ7efYjaYKzOZK
VM+Nm2zVCu02R7mnC45wtwU2gzrtZ3pyg5whJyqLVhLwZxHafjD8TT5TbGxXiL9mN6o4p3pNkpT0
NusmZGHAA3lDBOlZvcTkA8U0aPVlTkklS4IpGax6TmG7i1G3hM2gQxiRL9juWpJC9Eg0NwQoXewb
Igby59t2I/S3vDIWFQ8SM9f8pREpmbX0yhGOk91UXge1bSMvnNyiuU8AYSZgAO+3BnPNMd5ZO7Za
7tvav5jHJ2UGi/XeYhf0hraw4bOoK3CURlOoj0NHa+XmNBQ5FdvFgd0ME9xjL9oZPclVEBNQexZe
V3UWiLBvqbye8bPjkpWE4b/y7TppbXxoKhmMO3V/cHCNQakL4eje+Z29IjVxokvFD3vvXtczwJdT
tHxjpEn/xsQlGc4rLzO02K1lnQZ/ndNzwbHu3mEB2kFMJKRl4TI8OgxxbPiPTeK9qcBiBEOffSCl
BAHP0rGqFssq5kcQ3h+hviDKhSj7HRmLdnbCE/Tchr6Zlvt4sB9zLu0RcaEQrrq+JPTStQswdVvY
Ba8ftNZ3tUk8n0jelrsqfTOBJ0gckBoh3JYOpJBy236XbiQJ7jFQNHr3bM25VzJ7q0QWP+KFPT6S
Ad+kfgJldrTrMExD/43d7wKQK6TFuW7zpGVXN67UAVKLO8AZhMiPfEgb6JcgOmNtm7KiI+JSSfhn
KBVb1LIv9urVoKFHMJdTftIP25eGfYmynGIqNQmbFmEt1Fahnn+lRITT/2/ty9RS8IBgeKSWgVZ1
WR5VsuYqPXkIsWzXdNlnSSl1U7OKYd56Js9tFRUSgnQH8Hptc8aVHd/urGo93Dsf+yLDRZbKXxmV
vLEN2XAsKlOVB+0Wd9Zl4MYMEqzTeuTA9ZXZuLeCOQHucK0OViyS1UGLoD3ioP/pNnF3bAPNHccY
cIwpXfiJhqTaS4InUwVrz7cDSyhLMuAcyAceDx/K4ylfk938h2nMDl3JjC1QdBtV4LK2d7lZP69Z
bN2BOu0xgK5pA4A0ju1/TGIgzoB80IcyZ3tOZAuHVOB1EzLHyEc6HoF9XqiKs59awVp4sSj7/S61
IoLFvxk1RuRHlRzXHYYirNZuZfRrBQ0SRkVZZD3UrZDiX481MFOFO2buKrfGZhVtcQ/Lc9EjEkkm
OaPf9RjhlGrrXLquEPJMAt/kU4DO1QR16Ci+ptYTK703k5J+ONT8Eb59yB7Mw5SvZmE4KcV88w8Q
IzVyBJxDGfsytIl4QucL4RzdnudB4zKzazV6SVVYyoXtDbkSXUDNI0wztk7hAb52RF5imw4Q6bk0
hRR8CWeIV3zpVpLib/gZRae/T+Q1I4itQJVVEfAk+JRCMQRbTU7YKIvrNq/LcqgcWUbiQt+OqLY+
Uf+wZhFZ3eJ9/QEZfBFeqW0tk7DnmnhHo4rVJzdZDpXSivOkDZmua/A9QvWjNOARsGBy9rKVNxWk
sBG7zKAsf3mhjh+92IMf6bK8xOia4au21ot2Nz+Cu0Pkh+WK9vZ1VrDCNVWEaUDCOxo0pCCbvr9E
ShQLpEo7wBkKlzP0Hwn4yIbXtsNkt4TtukYrSKP9Ufk+SOKq6OKvLYS8FoZwc7GfPi1RlVen+zx1
OTxV9wMU29FZ64FHw8JFuT9iH++x+Rc2N/wirGzshQgQLeuLdbocNSeZC+2ZdnP5kdh6yI05ghGB
7fgaZ7HrT27xljqZsUi/6yL50LgOOeGJ0S5v1P6AV3YLgRcWftDoanNUy/uMN9+Z7Q2g/2VMz/eA
I4vuJONTLeO5I1CERH5onUC01p0BLaHskXATFeUbXfKDjbcDzTq958ZOx083RmfHbm+9WI3+h1Po
M/h8x6drs1u5bEgNWC1fuapwr2QLN5GsoryUMVb1Q6S/fEzz7Z64lwXx/jmEEKgp3HC/TaXQ70Ax
eMXNYY4v1yA7/n+zRT2ralk5+Uo8WYEzjy2MwKZ+k8UZVx7bnSsZcytSM5UoQlZL7pEhK/eEBwkV
e6q64uP8xRtsQe1mdBl9AD9yoFO4q4Q9QsY7Lwye/4LF2xtlEb6D8x2uEl4WkHjkIyVbpffyjlvt
4/EJW8aUDn043JDn++S8UVQ2cal9nqx2lknFCwwMtiI8ipK+7ViCUdfPpHllDMHcUHjunwKVdPil
IZEczIau/YHEc/GOGEGJl8arrCQf6ykWBkvVjEXJ/N/ijZ340T/v9mmwxvDQEx/Jq7y8A+3/RqfZ
M3BkCD5aeZ+Rq8GKR1kuE38qsGSKHime2hfECf73SErOBgUWtuBuiFlH6YpQUERJ/IL5UXcaswpP
dQllb4sK0LDCytHyevoLbi6IMvrEbXZBqdyO43nRSuhGnR0e/GEIWJ9KLa++Rp2f3AZHALoGGm/A
KYAcRD5goTJ1c8je6TdazvaDA32Sf+C4BLFtBDG0TmHJqR9H2QnVx1GtoeDhQeHXCPZMVYtjfLlZ
VV8dcnaXkz+jJpGv8agKAce2plpNJfk30Qhg61TSFxzhif0lH2+KJOnNUnwEU3tm4+Ouyx0p/+8/
JOnp5DNBs1PZaTaHbdzccqziO5796lYubYYvq84I5H4FhqKgiXxp1GTt2MVrcqEI2T/X3FgiSKP2
FTcwBtxnG6/YDeTZeo1ltmqghJzhkckGMPDx7wUkyhxl5HVH8ElCQ9DXVJ9SJDd5fqN/Q8wrXKVk
1hZB/071WeFOAm3dcLVXVsdhc5gPc9M7Fb2E5Z+ao6p+0ftpOILzOCjm1QNY3M82sVPklEcj+VrP
UEsvDnZSvfJKGxvWe8fOSYS26HXA+qLQHaC/ge4WIVJJDOxM80PbbOxW0WE8ML4QJaJXKaFNfIOt
O86ZlU/zzh6/6dM2S0dXOvNSXSWIfZlUYO4wZlsDjd1KNIOlv4qufe41T9zUNvSdU0aVbhFmfZxA
CTPHgVvMwliUIeMekcgnn6K3WxamAeF108vXzzAM6VyrCTLoXPFIKur1NcMcXPO2JwO5r/larDaX
Bk7eUcptm1gMmcjQ64uF0PCV47xf36U7RXK1zCo65d2o8uh1Rygg3b8VaIvQW79D42iB4f0kH+Qm
xJF4qfSl2GrTYn4Ip4bOVObBqPKT9FW7b9OfAJGR2N0wEOb7axtNPAPBuSRsOPS++X3M9olvadGS
p73Cw458tNswlcq9jWYP51t3BXa1wGx1Z5RBn14N4YRR6er/qqB4KxutTtocKVdLLGFODt8hSdRQ
JzMCGElMwg+yawzfIzXpEYdBIypAprw7GfzO/E5QEX23h+2wxUFObQ2V7aBYASNkf+6ucGGN24YF
W2bSzS4QtEmTrw1KJnohZHLIfLEXuvcWnrt8U5vWZctj73EPCJqgCtB0Baa2EXhNIVu5+YKS5Kx2
WbQ10l3gQ7yMH+aP34sv7hQUss+I9o5t+fm2aDG4aP/HnWcb9esa9omRwy9iMdk91XXiIyXmWViB
vWc9rCyBL3N79a1nfpWWAu2Ko7QeObWsYdT7Bx97Zgr7xh5IBtXz/WrAruZa+GwoOVnEcDJyzPL8
5ufK7cV4uO+0R08ELk+Uk5VRVKkxxOlVvhlKEyUvyFjgW4XPQtf/JxKJrDNxLZn/GQ7+C3ylGWnk
kcaZZadch0RtHi5WxmQDILd+Af+pePy/pi9nKCdb7kNxCLLmxSP92wkk/NAIO8lSmYG6ncPle5FT
vCea5qM6BEYUMAkqesDQBON4XNBlMMcbbdKVKoSyPRG+r52Q7+m/HcK3r7klP5BBjZu7NzMCXCYz
ya5Xbvqv+5AQCoYSqtx9SQ9AW2e6b+4LveqUnLI9HAlc6I64MMraC//XF22/mgZklXUAeEASfmmo
eB2d7RlbzHqxXf19Y8H2G+hgPkIuZjuJXA/jKPpS5SGYweL7TpH4edMDaqM+43h4xgGusWk9kux6
upgjY1iTyA6dH/1WznwX1iR81pnLONBdinE7UgAdC0nooeM6OPRlMdnHMxNxWsdQas92v3dN24MQ
MrSzXnXIBRSjTJ6nOaulcprr83N12vRLtf0+yVxyKU3Vk4Kdm492fkY0H2r3V3GDHAe8pnhaJSoU
FV1/JeLFlLQbte8i9M+iHXMbmKoD78nLLEgslNLY23JTeRQ/VBWpOq6aZDOkU1oQ6pHhZAV+EFQG
AcHEv6mJHRGMtCfT8HzrjU9cbNWjE6RtZkpeP0QYkXKugzKMatbdTxeghFkiacWG14td+RNTbKT+
ZiNs7RGph6+am72iCVC+fBnbtyjldgwpgq4KAJumzf+QTwJHc+E8kM8YIybBcoYm/h5URxppCoBw
jb9Gmn+3oVwllWS38Ij75aDlY/IDenWYvHDbLL5q95bNcfCZ+cmFBRpDPs1sPX5rmuWEd94JDwLu
0ORRE5d59u4Xn6Cn/gFr+/8ba+f9EybhENWkY1w8nKuecPgYzoGnKusxi/kGl6Wa+KtefBLxDwq6
tRuQK07AyHVfJ7JN4BuvGlSfeR4QsduJaD9bRNduPCUiEJ1fhjELfileHrgiBwxb2uFbeiZiaiZl
uzxoHvTCMBre2zBIXGPWNVIUiQRHQzEORX6sIk+KMJndfP21lbJycsl9PgLI00WZSpqFyBMu11S9
vi1OaMn6DQ1/659JJBE4n6QBZL5NUi8fAMWz7QI7x8ug8r0Ife1NTJw0EAacjJCJ+aQ36Jsc0kzA
ilVa3KCOHXjxrFCFQLsbp2Jgg4raYAnLiudSWQoYjzHHbRNqAyIxzJQihv++8pYswUP3QGzF+0V8
4YdQi0TzLg+3zKAMMY+yFsySAXHXHtTC9honX/GSME8slU/q/7PaumWzrWQSBqVRiQIMQSYhEY7q
7z3cKQWSYqlLw+vgwG4hfljvZqu9bf2NcQKEGUZUkzNoNQQu6Ap6LF3HQFe9Fb3CTaCFsdkj5lZQ
Rwf9zljpl+khu/WvKdvXWpAF/NeXHXXUz8m+cDVLkA5CVGH7N0CeNFagVP2YkAW3O+XFLgGX0SWv
7BozTMdDtSykQw6CnF6KapQnMhsX2nd1T68Ew9iF3pDq7m3ISpWmSuYCZ21gS8WFw3NV67mVA6YA
wBfNbhDfdVNH3aQr1SjQV5UMqwkWTJqO4TL4E2QjDQMG5dUKi7bXAlS9T5AlBcpEd//GVS7fWMcp
gjqs8RV80E0g/o9tTEgl/3BDV1Yl/gdT1rBqXo0hdrCc6k9RDEoBLlV727ZYLxiF1Td2MNR0tBte
4GwVydAi7UKxamLwajUBi/KLxLN1R2e0fWGdAUyn6J6F2rshpe78w7Qzswwgvsp7paQIGHmH3J7Z
5teJ/Rj3X01wsE7Kh5bqkcrjCAP+6GRX9uRWnTETtRQRXutQ5V+k1Br88yUvq4QYOPLmrUdEVeU7
E7L3ST/IC6e7YPmZnhXNkG8cStRO4qGJWi7XmaW0Y/dY5GBXmQy8OeLoO7Oa48kITGvtaF9zSWGn
6vI6wRPakovyUJ/3+EHPO5ARlKS8qpc63Bx106mssbXvSuCrEaRuxKfLXKWyyTpBCmQEjPOjIp0n
LUNur04LABvDb32AcZfYCEPixX/D//faYku3P44OcKPHCKZgM1QGU2NS79Dl3O4BknSLKjCMzoju
q547vwnDhk84MlMHV5erNn3sP0nVfvq/xzu5a3KUEowlDMXcW9mAtaSOe+klQwvqsIiA3HBx9pTj
t7eRtmtD7gceYmnP5eNLdlK4fGbfAlGyHd+7yyJiyB51CajKgeQOJ62kxKdrREGjBbslRMClGtJs
kNLOyoHQBdfSoPqszUb8ME0Ai95C2WhpcqFH0rtyBWojXhrEKJAe5bADG1b3svYNSxmglOpky3DN
Qn21u9OA4QR6HPxwTHWyYpRitL7wLIsZbt1IE0ByZFPZLhmgPMDgxtSsQ/xCkHj81EcuU7SVZZE9
nkchEbzMRveTGiWj7FO9Bm7kN1OZMy4BC/pM4kemV/50LsPUVU3Yfoq11SREidnKuffb5VSXKdZr
mdgOSWyNgtQztP4QxjIWiy13/khT+eh4+SYv/CZxOx9RVwb4umgQeGR7o+ltRZ/YrOT75XxcZIIB
Jsu38VaNwnAPbsFYpAzl1ejtHXQySLJe7WmrAj1Csn0J8Nc1qCpr4a6eJIT9tLPbDWHSQ+1EN6gC
jeDvNWXnYf67sXCp/1wJg8iFR+XEbMNGTXDvGCkjyrHTIRVBlzhhW0VzJZc7bN8mmqOzKrGk7HBf
Pzt1FB0U/Cu6ycOGIXnQa4WRAIrD7hj0XHZl4fMe7tZNH9CxRrmb+J4dl2q3rHVlN1r4AeiquVH7
Ro6etliWOfJlKJZyblXEJTiUVn2n8cIuaur3xVpqxAu2IMYLV2CC/dDFdeDuALdtLAjOHEM/CZIp
Q/Rb1CWYoEciM81yCIKrQAY5avDCHfKIph7On3dcQJxaS5R7qpUVW9NxA8cafFJXGdN61zlyWPjY
KmpH4eBSSXdcCVBLyxCXJm36y5cWgQszIpnqui0LeelQxcoVQbihPCuE/5uiQomDpudz70jxBYSv
Be5iTWK4T5oAL2TtRTZwKxZs8NqmWm2zxBlMFBlPbwhZUVBfoChawVhH+YpICyKkVm2a3Km2guhV
pJMIFVeeVjs6TCWHx6CPSQGC8pzXFT0SKM0xDX1v1PNqDItchgGBwZNSzVxE0JbL0qOua/wNbSDj
u43JD8+lhozgl970tW6ZvEtWYlCRHW2lJLhTNeouk4WoU7G7edytV31LWrcd+cLNliFyX9k2fw53
Z3/09mRZRydei8kHyue01NpcFjZBt6Kd3T9sVvtV3OVuZu9CiVvO+vsKpElpDQ7XTP1rAWQRR98H
xo4qdpjlQPhrM1sRHVRmp+RavGmj9JTSFhIZSEyIP0YwR7kILDSdf6aDk7MN/JrbjwgZkW9pm2EM
Pef2ROZgkPSo6p7168QYEsEpXLmhZVLiJTJ/y8v1mpZPr8uTFG0piNZPCJUBlTfx7JCAykBj6f4r
Etz1mm8IBTScc5IQEtzL3x8E2BpYIdG25qEaL/KPpnvphg0wS8sZUBwa7m01G9OPsHwumjQvSqLg
c1Un7EfBMhhpqiDhqyNaIoPVoJ7r4dMpHp1ejl4ztid0SPPFPHv25Ph85U7ugyCfOvkUNOCfC1Wu
gOFgRmLHDguAAQD2zxmAo6RKF9XWNBgg20laukBZLaOxTzRlz7i2QCgqjdnFzRGlnyC00yN1+1so
yOKs5lDYdehz9Vg6ztyOEbLu0NeI568yG+X7/YpAuC3nOnCLlVkhI2zjgKtXHamPhHDDiOz13jyd
DBwdVtyZcDKOF+ZSW05Vuqea5gFlOp8NqjevnCMbcV90YaXsCYHadJYxo7Vd4Ro2a2zIWlY16khT
F+fce9sq/snTEQfW2sDFZ/VoIqd2lsgViP6M/4/sGoygQycKPzA5sn64nxSJxBXd3+R1pr7vo9mt
MNe6h1tU01qJQpm34Bwytv0MXsSJV601zB01maS/N8Ed/5s4IKgVDAFeDnJf9lIaE7sWvQxWAxNJ
7FXubGCsNgiU9i18COTl6GrORoCfPDGdhASozpYivq0LME37gxOwFVDcif7V8QrvTgPUSXswXbXq
18hEKcTx+p1kcppKgsyfdfmdIyOawsoFqoboDBWR0d5X20DsTnpUAV8hvuPnVzdtnsoBJdcdXcw7
qu+Yz+aM6FOS7lqsZd1UyoCnkf3HrVJsD4wynDS4UdUcdAlW1iqGfeLtkG31oQPeDj3r+Q6gEmrx
Cg9c28VgIPP2N3AFZ67YrysU/0YYgG7S4SWpK4EhQ091l8OkwS4e8bDsAIHquMcUYohXhymx0Aiu
y7TH3dcaG8h6rvKEhgaIqcf3XzfU0G4gyZNJku4aTFgPZjhYGnAeF/IgLONruo9ywDDTfM0BR8QW
36gYjHGqU/9rATkBzs32SQjXZpVqVjXkUJoAYIGLY//fs90vpwVQoGI204dze+gB+rs24874q6GA
tEBxOmL5s+BGfAJtkea8TvVm2hy7lKgYqKTo86L3J2VAatZ2iBKitlOpho2dOcXZe6VaeLDBkyT+
SkYGGi+O5jJuExlzSU8f09v9fskOIJmyTI45Epq1zMb2wI2b/4LLSZJhtsliP/ylDP1ihboMB7rd
UHMWTuP7lZ1TlYD71KW0Kt2FIYBZ3fO0WzzpjmpvGYE6DpufbaIecrJ2uIeRBTKreLl21Sr27eQ0
D7wxUrZbzcIwLC7KaaJ8etvGVDGN6b+RtarDv1SzTn/uah8NTAp/rG6/il/tiPUvbZHli2uLizA7
WG9v+mIfmXr0g/aMPdRMBR19bXOeM+TUVMZi+PxBkr9gYRol2Q7T1D+8+u/Sk5/iRejOJLuGDl0+
IK/I6WHd4tzTz09E5Yc0aVf2Il7ibSRGsQcDafRTSWfPPIRitsdRiWECJ/Iucl/XpZFowsUmC9LC
77fEmMz7jiq8v397qWf2YJte2W1SJ5UgRqTuczyao/sNy11KHmdoueLXUbrj9TS5yWymdYsKHDiM
fUJWyntzUviIgd3STYbJl+mXywbGOh2rn4rQ2BkskvTiwnQdjvbcb+CmNwMjF9RTF6xd1GGIrq4c
0dvJY92JaMATab4Vp4jRWUDurYYSzE7J1GZiHMhHMhzn89f7QxHSywj5rjnRN0W9CSXYqMqyK009
IM67Z9LQLFGHLuVHLJYMxwYtzNx1a1aMRHEf0qQBGykDeCX0mM/GrLjCoMiydIG69TjBQY5IBxM/
uUvJ5tWMz+ZvM4RyzAP5LMkzeyEIL//koHDwRi+nVwe2ok9Lb/ef+A6OBmXo4y4drjjv6gKFQV3T
EhZbG57t98AUTZ31F4EZdyn02BsRrupTV2+w5uz5VyC6z46UOFiPJwHR6BEOkKIzaTq4haeDRK9n
XF0IGoCs1qFg0U392Q5sRrIJpUnLwT1a/tzj22zXAZj6V0PlJdIp7VmLSjp9QRbN0oBtUjuEmK07
KwpnwDnbBWuUcIS15DG7zO83VnRDs/tXrgkhv5mDVGfcPCeUkMlbNnx1VMCXr7DKaVrOgqcxy7Jr
Z6De8Etw1Go/JguJbb52lWoMwOxlvbYTlZCs2ngvSzV9NFIQgDjo6NPT132Br53UqZilnp05cij4
VFa53RBjjtNqYPO0KU0B8MYjGC+4fm8kcklwfQ4uhQbvxSEMnpFExVnrO6sz1YkIOz/L/y6IKHNO
aSSNX5QyMgNQuOCjDFRj53nD51lwfotU4oCE4K19k4tkisfzfEQSZJXuUEI3+0gc3KsGjso1Zuc8
UzvsIDzBYWAuSvB76X2OPGIEXFHTK+qj+p5pnJYuOigtzGqWNwfiZ//jztaMnR1slPYmluOKu/fF
oonJJ62MVTraNnHjzvFSvM60ja9xR6nTo8ndG2nnl+xTDDvpL+bC/kkVDhLdR29UUPvkBGr7IAUL
63VKLPkiGA1g7PS1kp2DHhyZq7Mjyv4g87v5wNvodLZr5ljGiUTAp0UfejE7V2l6UwO70ke17pRO
5J/1/CTh5WnoaHRZa3NdaxMkcg4RI8SnshoXPLTnF5uyleSR38C+IPiDqcMNZ/xO6m9RYeSHoffJ
7K+RdkZwio0h/sCqO9FJ+/k6yHnLJgViA4KrZhA7Pey6k/9uaOn2GUVikfppXDV+NIjQKGKC6aMz
m3VfqeUfR47xHq93RwStRUmUAiIxjaU4eJPhxv6KRtP38MXuO9K9gvPAL/ogcd2Q3+VShikIKl35
fJlS9s/tKJufm6fWHgQoScmttIuGKf+hQH0r0uQJJB14U5Uoc4F8lov2/Z3J7ngDh4UeYsH8/9F8
GRzPSWzvpMa7P3ulUgSuKfoMLyGpqqa/QKNitaxS8e2SVJWADZxONFLEirg14C2XHhz1NSrjGAKg
QhSUU5XbLqRfteCSJztwbj7D4oZUdHFlXsm21VFUSUT4e6gnFcag7dZiysefK0j7wN3N9wFdsbzh
H9mtyca23s3ibDLN4XTUMfSS6s3BpfqVxJ6doa83b4p/Qmd86NCHs7WIZPm2Hq/W5slyJAdE2+/N
Uw6jHh9A1s+V42efgBBa5uSJzL63Gekby/NiHyPCEyn4GRheF1OyUacD78w2z/InE21yYaSwnqB2
Yq0atw+oe2Gv3Nnen+3Mu6mPZ6ayWkic1CWQhhBDrBazrp7N1cL2Vq7A5w4iF7hSjvEHnuIpAt7v
VTkycLAVuc/+l76DqhHAPlP+AEnn7gL7nB279ByAJ/iPPEJX7D1ye+GyNYU6WzBD+JYj/cXARKN6
DNBNYDL2TRkUYZ6uMq2z9N/grO7Re71KwL0FhoZ/ckjD7kfLmU2MVcLAKpRJDbkJ1fJga3/JRkJF
nQake+de3GKo5jExSfB0+RFJ/QbZRnTNNtnWZAQ00EOxcwDAcv13i44QTh6qrurZhr74IgdjFbY8
ucOak0OJDGJHCLOeWocAskY1ODmZMkRhDDyTfJGk1nLZ1g2gqIqJwCMMssGgwH1+tB59Ibbh8K8H
2Mn5P0GJdSHkb/Z+RHlMPK3CqpIKbZCuFAFDj/kAGILaruPkpum8WCcGaPFFlFTb4gzuhEsBYi+M
vpiV/AvyQIpMJkitFIwlmLdFC2znjgwX6Wh6LNXvUKSI1AaddhiAfGuVk8O5dVI+LUGjkzK+SJnD
HLULY9NP/D2ejWzZgcVDnCAurC5YgdkWaQGuv8x8SENXAH6h6W3IccLIN8bZz1Zq+g1HQ50Ew/tv
zrjPE2m666KiHFGjEdEsOIMGCrjy6T4mj8B8wxHTN0Jo/xr4AniZHNE+MmNSHD5OGDMle+cuwWBA
CuwaA8SVgjUp/pJZI/QXXH9Zjks+p9RYuepQ2Tb9Hyijk1R9DGeqZyv8SijLXHrgsBhCSW0rXtiD
RnAJ3IwpaDl03IM5DGURA81uF9zgEd0u5FwJ1KcjqgDQMzgpZVaTsD9401j2FZi6w3mcOrzCE52F
QLCw0E2DN8TxlrPXlHU4jQyIfvzZIkwSwrD3Hh44El8KwJK3u9BLgkXnCtklJA7JpvoyrpH0UzFo
e8XlxgG3ovsDZqHLYIBb2DLTL2ojECgrI3Nr6zTuwNLK+NSAGqqYE03C0Xt/Vs4c2BoqvpeGumDG
ixslml3nxVHLYeOl9mxLGBXP3d0E3i+Nhkp5/7RN8SFRhFzdZwB104EN6iq+RqBTZhYAtX+UQrIn
SEFz7mQNCGJ7Y5T9S9pZBuSZnxTTyZHCVSAPV3XnGq+9u2kVA29o6/QA3rfYw+yNV320svlfDZ5J
zUPhT61MqRaG6TemaSEggZ2VDRrIku91gz2SpWmtLgY41EuOhsyq/5Y8mNUbtqjzhSyyQlHwd52H
n0DOY4otd6bIrQftspBaE/65etLKVg73werTZByAjwwFlDO1YMu8dFrCD1Wulcfm8yUTNOy0leLf
BOIJ6JtPP1LhF99MEipJ+GjBsdNXhx2vWytnU1c4WZWWa1PQVdXrCionp0XVCRuCCgKDMvnp/57A
zGU4J8JZSuGl+gh7XSpaYof5jB4i3poc8GpOSh/tuP48/5R2Skpq4ilw2uOjYzTyBDzJHzLESwge
HbEP0Jf5oA/yEzyVa+cmSdwST26Xj16qFQ09HPyc3vovwSdoysmkNO2Gsw0idhAvUideAvbBLd41
Ub102nz06tFyGAEo4eJ97dS4XAbRe6OR7lLsQKrJgyslkrguQUqQ5rBUXvUlaoIO8+Y6OovUQAbZ
wOLANEzjIKDH2r8nCxCpxfofhjTpzpSpBbZwo38nE5l9yq9eCwN12YyD1/7mcCJrxWSqTj2NVl6V
2QsLPaQTkl9uXVa1KqNKJ3D6oFZddB5ZNX+EMm3PPXbUbvZXX3e1Lx6awm0pMn6KYoFctgoXt8/v
wNrbMB6Fs5pXukIW56gm4z3Gw2+0Eeh31LNlVlpKX9NQXEDJaSOOdkGr36I5HMvnO4U8RqTOa57A
KKwz+jnNCgadnS3/tYf2FnQqbPxmLMUWg54uYdQmRWM0efmwRTM1VNdmVkCrB7gnP2pKHy6O28vr
sbia+nxuUbn7fDlLpyT8h6i4e29YxRRoLjHUGSc4xyNtVn9+jpFdU/L8t+mDo/h3aSaT0baWr4fg
pfKNCOdlTbiBLZP4+sRvcoLQvATis29p4gKbppC6rp3Mskl9P8DlRNCSMY8p5HX+2cuZEOMmWChK
nu0d90OwpJuJRNUWvwbfk6wMKtkmLwXjsTDC10vQv0Pnn3dfbrLNb6nC5tbVWxO/m5b0GQ+vVoW+
L45SjEACn7chFOZ0vNnVVoAwjoUo0J5t8kXn7EL53sPedJDhWLPRmL++lvnU2vn1q3JfqJsxbYRK
a3h6KG2kGcm3YgXJooyP+eQNHG2UxqAJeJJ/U2f0RYQxtCQVBP2izfy/oEIDd9SeLKHDlT258RHI
/P2+3LWkwoay580QB8OkZpTdd1tNDo3Omrt570Kf4tjs4iwM8zJLFL7F8rDRUxH0PTG+7Wzv1Tvd
/cnGHYDv5ZMY6WU6ncFBuJzeES5175SWYYURy0gRbCpJG3Mjz/HYiCuO/g+PTSJEKJjpA2jdMdoP
lQX7nds0rE7Z5oArKDpJAcbm2WQd87qkH22UB+Q+bmRAQw/Qb5C8pdfUVH1AwxHfmUijqPcKQAdf
p+2Nsy5+YNy79k7KQxQ2p49gXUcg9vQzsHeQ719KZq2Rzy0GM1MagpJL9VYp3T0gqovHsAS8cfhX
DFsz2HTe5PgE12frZI3xCvIku4nE4qq9StwPNP2saZ8bHuDSYJX50TjLEuDdbTS8xsi6UPU5rE3g
BLsg3Wu9mBNKeV4xEbQXpxydrpROMrCGX1drTLfeTx6s1Wkg/eonDrKQ7GdQjCR3DSu7U0qQ5WqG
12B7RGTLDsqNNEbIyycXgvRSCU9IvoxSM6rEjADHKpi+4DzBbIz4Uv+RmiudU39yUBEMiIhGXy/n
1bigRtsDqXmRP2fDcEke+e18VPPNkt6R+3jnC0p+d2BQP6nS3dplvtJfyvtDIav7bvYZK5P5bPdy
12ciM7OcoDFTh718KNdACNWRskyEcjs6kQk8Ks6HgWaxWJkLPDvaLagsTZo5T8SYLszUgQFgyjNH
Xv0xkdID09C5qFuIvYd1sGv8FaozkLl++fMDpDNy+QOvKomA3xOdQzoPVo3PW9/pPUUIkebjxstB
bnaiqfy5tp2tqb51aGr+OTu+qi4p/Lk2ONiaYWPam0jbe0BsOkjs8PnvmxH1MPhFWdwmAljap+mS
z2+gdkAoisTWLb2Png/ZLOg0lEzu1lhQz+kHedkCr+n6F1t26zzH8Mi2QBJeQJ10DbWfucCvn7WA
g2Fvi37tg6eciNgrVJFMN5iP4sD7Z5PVOtbOo2G5b5v5rSaUxZZBneAxwflmIIDzFKXunb/QvSWT
qqfqA29VkTJcGvcluRy9etvSrDkpjEbUC89MB4Vm2QLU+vcMELibfzWYJUB0a2JSAgSovlL+OXaC
qkMIYB1zDzSbQQv96vLNuiquy6/0mhE6kJo9hsxK3SFe629CJGvFugo817BMpdmxU8dD/Aylj9vk
bQhbqbxn5HsMSVJzbXjQf08212xodYa3QuQ6f4l97VEsDnoywBUR2351T1JyhV7QVyiqtO9Rhvm5
vcFUNswhywRmQvJhrg9HCUZ4n0Z2sjvQfbSlwDZ2T0wiI1OLNi1Wc0PCJxQxZCDqLvRo3SX4Wci1
+gzyb7OU2RC8wFG612a8wElmg5WRpI7UJ+5fp1Ms3AIIC1arYhyVpFTUHJfQ4WhVUB+0D69p68cz
rm0m7iZvs4h9OKgn13NcF4e/BuxsQK3LcaLQpFO7tAQP/BKncS4bbjJjpnjjzzZbI6j9JZYuR5gh
eQys1aCVW3DQXo9WpSgdqT6IRCTx0ayMLy9rz5/MyZrbhhWktkHaJCvYBxn6fupH8GrW+Ll03Pig
WG8MRmfpewQ2Lelqw2slgwjdNdQ6kGzFD53e1Ig0xQhl9K8y8AJKp8wrZBrxUA3Bw32TjQlEsphn
BqQYysB0nae/nLDOf7sQKf+sxegxVn4iGXc5R2gq6FDK+63S7RWLKD0dqB+IEGeeGagMyZcrOTN6
feA0BY87uTzzKbVRUDJCH6bXQ9avz9bxdt5fP3f4Wd125RsVGvUfxHC6BX8gnejvmL39MrLTBFHk
J60OneED6HcvyPiln8maYiChScPJrpQ4UBKXLPMcBPRovv2T9RE1aTYb9/p/5qhrpcn1XcoW8SnK
eJqzsnHRu/SBRQ2g3Xh/Y8DN9gChvdLDIlMolzScC59XFQprww40NXDrhynKATWidHlunO8W2+uJ
6XQO/EN0bjHEZkVA+60AqtS0evW2Yq1x2CLHV5yne2hLLSRJRuB53H8yYKPxpvfoZuNGLc2wthHK
FSP2txh8ojbQN/LpKWslhhg+vxghOoaSa2hvzwzSDs0g/qP+9YeQZLFi7S2SwVn8yT4QM3RSpXyx
P1GXBVTdOfITGfTT20Wq3akK80ZqKneh9SMM7Jm9zUusbaRpC+yC4x73jngXr3DxcYPr1+chZoPK
K1suModqYOWIbC0uljZhuLlmdGkDpcZHSu12T/UilM+obmNhoy2p3prCqSp1/kRqe8ksjvyDi+5Q
YORyYf2P+pWa84XVHoNzNA7AxOH3P6Ze1wvUQ9yrMj99YX3vYfnBTYuIymH4u00mHzxlMHgUT6TB
apYZ4svK6Djpzz9ZiJzR1tugZLxvO7uD8UhvAzVQj4UGLDc+Ws0Z5dbUZT/ZAvkSIVRl7wk3HjZu
TH8b0mxkL4xqKhWJFAh5IVb8BsCCgbXwZXEs3w9hD17k7fHyHOROJIEggfvIi6qzRWWUCFLe8/48
fpV2V0gYnqBjpHGJLph0ZFukPCF1PiD+0B0h1vbwlW+C0Kj2e0M0WD9d20pTG0UjMoGyKH1ZDmTe
qyGFxmeYTNFp0NCAC0Q8qpWbNURU2ha0hdhs/UKQ95tGktsTI1hwjP5FEmwETlwBVfIuLxMzGayW
Ld0Xctlrjzwo+eIf5NfdtPg7NDrLnKq54YHzKKKQAPgeHuzOMyTiZjcRfp5a0axcrKnEO/qo98JW
+A5a2mYhivU7JgOJLMd2dz+Tei3yvxJ0yI4GFPFoo/yRk0hXZE2NMZ/4GCdbD58MbAUi5idK77Y7
T8L0oH+NmtKf5Kl19giw56tOgIqWhBaJGMpq4vciWeNW2wkhropXAdLyvYR6oF3SNJRi3QlGnkiy
nLSUfWub3gLRgnRRZ+B3b6c5epWlZ5gWQHHoQn9KSwCJVtddxCRW9/X+0bHpXpsLVXlg3SD4spdY
K1BNntM5UDJGGcn92MNpa8wdMSjgcTRnsUo7BIl3fmRnHEw7yAj9hSvtVT5N5Cw1XmOJdFzCdWv9
e+EaJ/WbiY6U0Fkt9rFM57+5Xx4KOPkPS+IiNQrTo0WdmLuBy7XBnpWvBlVO1uvoXili4JxjNbTF
sH//a+k/79021ktio4iDPcQym9dvkVbbRj4DM9UJUBd1wwS8ukMzSYMMZvhg1T8+hNcaSPuSF9dg
JeUUqs6IiCuJ1t+Flfdaa913nS4zLA4f/7mfdE/JSzjWpQVU4t+Lm2hdtt2DnAF+Ie4Ve505SZ3q
JAaxisXzddtyDNKzHhQkD3SucACb2ICglVB3JkA8saL/3bGc9x6qDcXOjWE+v9mY92o1QCb95+Yc
5liXX0ORQ3VMMU7jcvhPEB+oIHGlGKL2IxwOHpYnV++MgBqnmr3ehMwd+oMcrEprTzi/ljJ5f2iK
pCzjGfV9En3Tb+YCzB/Udo52WMvhFpZ8tZqpoH2GbMDxz7PWpAWkKJ1FizFd4qlK3CeTKJvKjkok
XK39hfdS8ESc2mZxwydIwyfy1504gee3+CHOjD+ehy9T1p38xAM43mDAmuGDYbxzQWvG4AFNwe/I
tOcmInLqLRvpLV5cVt/PtnlSxyDpVP3GCDREi+599A+MzqxxrqzzK370V50i9umQASs3zMiNc8bx
Bvbmuw+vu0vDmK6aPNj9QFH+P0Kz+DkHeJo9jwZdEt3I8kq9X/qgrwKUjnJ2xZttnI76qH8B+fyF
v130Bzl088oiyEnc8MCJjIQn7K/syNWBjKMokHVC8jLHdO4axopoYrjWrYN7zaZlEKM6W3a2b/9K
wkaRHOmex+MHrwIirKamC/el1XXXXHBophFdcSNs0Bkl/cov2b/xMRvwQ4Wasy+GrldhjJ6y2ZrK
LKfqKVfmDykJN554j81v8yxExLDpfwiCprawL1sBbxwwViLF6CBctWGOZhO1l0+LSB91yZ15BhvF
7QhHftkA/zISWjTdBrzjahfRu+pbBV8cH8ljh76eDvaIGqAadd3F4v+gpnqCrokZMrEgjCInnlWe
SI1zr2YEbrsBnjgYwsnN4JIvvXTBRXPkQTaTQi97y4K6ZM8/RqWYtdE4q5kQbOi+wRv3lAtF+mh9
4+3Zi4DFBzOGBbnBsT8sX65BdXfzxNRoFDj1Dk+1Kh1uAQBdNv43OHVomIbwAMGMF3B+RF+7Eokd
5oUi7qozLUAT55fWkfKRTlNvwa+3YXW+NJay9sP0bvGRTKTW4sweRtgV/8GsdoobKKX+OXjKQsGc
w7Z3TxmI5r0lEqqVcpc3aQq0ez0p8GUVc+76PTwsnMQMs0dzRecZKZpHClvqTQUq028jdYV22pQx
x0DINgLstqTrRmPENfw6YQt3jX8kLx0AUA+dD3zHvLUWCVFZ+G7Hg/4dLiLzS10Kp9X+hKWbyJYV
AuE9ZlJuck0EERjn0TULmrniZSEtICAd0belh0UHe0IaM1GLaGl3Xu04pi6ADTTVT1jNpJYE1fTB
L4MWnyyPd5tallngUR/uRKqSnSG1buttxOAzawDgmGw3DavJWVD7XgDKgdZPADv51vzEoMJneaEb
GxIDmlmdqjORj81u0P8/VpMkAzjWyd1a3QpbkufVcs+lnqKRs2nOl1aMI5lxhRcB7kO8Qln62CGs
fEnNiV8MZx6/5poWu+aT0m6UX/HAzHoI1DMi4RBHDR4PHJs9q5gLhhyox+Zwe2sBPdhB93VbqkJW
9HKHZHaK2feWgRm4aIqNVK7seL+lN5KRg49R4qi7skvG6FX9xs2b8ryaCMWfW/kpEnipvQi+kSdF
Kb08mrErUcDTua+Qn7/YntaTqZV3c4tSeICZSWOzUHoyX0KhJQRpA2TVHTQF7GStYhCQvAONKKED
gNPpEjcBYeXNxdaUpVQ0KSi59jsjN7bECECtJ5UvXvuhmr+MfnyunaPUVohX/9o9aczOD9HNC0T9
iU/JoZ3maRYqf++/koy02cN4pUvdjqgrZDgwots5ynjYLbC04f5bm7kZslg9BHiA1sYpveY9lpai
sokxf2p8Ht51xGraZcXwSonXvFP5PJa+XyQQBVcjo5Ou+pT8dxWsVGDFfxyYxA8KSCDvxLsqvsNi
jun4b9C/DPf58DL3wyh3xdMowPl8IpVn3ppGgsa3hVtOpRKTS0icamg5Ka9YY3B6aitsvspHI4T+
S68lTZfTE+phWq/U5hSaHsLtPDuplJ54KqkXSYGBY/9Mp+Y1o+zoyaTPECg1k1yrgYt7a0/ZsLZE
JSwmJzzmsNVk5rIH1+IZxim7wM0wCfbLwb8LY+hnBL1gieLjrL6YWFjAO02E/KK6mPdrTNjCBCYu
meV6NWDHXa3Pnhr5XoWTKKZK9VmqVMGMPtfwVHXaPXMUkr2XblPHzGlWDhnfTZ7G1+ukTen2UQ7A
uojIEahdjK7UmFrpci2z3qsXtXMvQZpEb4wDprQIBLa8jiz4GN/UNf1DWJ7fhWOzaL7Ft9n1SREk
/iN4Hg4B4qwpO/k94URkq/bG1QEUL6H/rFuMSOK8zsVWtfvsSsRhaQSZATBvDYjgMDuiAVBazeno
t7liVa5cHJjoe99fbP9gkUTkjOWFTGcCZTXYUOSHhcshQmj2A3JC6DndkOdLFPpQi9ccM9vVmGhV
XpUz1NdwmE3VRLnRT2OQ2EtfpE7XsIwy7LEG0QTAM6+JabT4B9YoAMT1VrSYHdCg1SpaSGDKv35H
3i9VxcA8d2JA8bhB8A+NsuBuiIht0nHU1zv1C+NHYs/4LA0KPDsjy9RS58LVdd7vlF8ImlqNGT+v
t7GBuFSkZ6Vj5+cl2E/FDQU8S6Ltu756nkWBLMj7+YVw5Mt5k5LFsPR6Qq1bNaRUPAP/wKC5vhGi
t8s8FZfAkQwHnI8HN7q7iAxQ2Nq+xrRsSgboLFcYuliTw6opvcBrkKD8vBFe8wsJki8ZgkwCwBzD
WiO6A9zl5auxS3gIQ+ULhWR+139dd3J9FoA2gsNoZfzK7Wa3H8WqkLaT9Y3poUXzckvb3XBQW0b+
lldVJi4633cFZdDfMK6eAKjN5utC9MMj4yokrceJjm2QQgJlPvVhG97ja2BHVskEI6A4nv4gAPiv
z+NFk3K4UWXhcQqTnwJEoIf7KUY/Qbr0OJ7LD6kVKdI7SDnSQMZ1JGh0sewWGpq8BG/yTrsVK0rY
EFJVhgnkbr/n82li1VfwQoh8rwCy9poSCMwTDgA7ff0xJAVF709u0soMttzalUySZtjhvbJMSMnk
gA0pz0FLdtw1v/NkVzwhUdfkbSgJ/L9p1x3qH5IhyzF/saU6ARuEQmmUWarUpcOJY8L0myV8EW2w
oLyRwToJlI6r8b5qN8u/n5yZQ4I774IOwBSI+NYD/w8Nk3tuRmfVZRvZLJ8AYLDCvFJhlofRQKQ6
WIcEQEI7bkThIHTmojCA0VAtgR1t9Y9VWEXEjME9SNiOV7ZI0Jxzx2xBoei15Kt1K+uaWsn86DpZ
w546IOWJV48KW1/slxHbpObpEwPdPVAJ0HS+L58onAFcNAneTFKWyQqkpAusoHj5vPyFh/MAM+vD
tEbSIgSCpuFu19vk9BPetG5n2fmu0bWmJEObgcovs5+nJ+Cy50mtg6enfxlO02tw/8qx+LMwQodB
XeYzyz41TpY/2+NFqCubWQG7HLd9sAuha+AJJuQvMVSHAun+djLBJAqNwDGa4fC4Lel0EISOTAwH
IeVr72T2Zm3MEULJUmO8YgYJbTbUUd/RzH0cqXFSWX8VaZ/PUKMWHapW5XyKfL+3HAKCveDyXNq9
XsZpJJjqS9gBT0Nsk92OJaQe3J064bVMDPDE3GWtr6MOQqIf4YXUmn6R/RLzKTmK8rD37PyHTikf
Gu2wgnIw8T2I8m8Xb8zoT1ZIeL22h3GlEfb4/HGboDxxw8f43fsCYdn9zQ5QRXDL498t/cE+UBBz
mX+qjfXxVL3dhCk+SKQ+htnKS2c6Dadzl2cagKu2fCqtxikbP2sTKqdYlbnEgQ+P6CtIiWjaJ8nl
wfCxEauamTTRaoPdoM4kB4vjjwhkXPUgbuBxu+NlzR+9blmz2Cv0eMeyJJ9yGL+AJ1IMNW3bp214
/oSVgFFM1EG4eXk3/kHg/GAOOfGVf6xbTk3UPQLWLaG+lYqzv+/zC71N9vkdZ3ch8ea2L+n+6//d
JNPGx35/PlBz5AQcRHfeJPLms/HgU7gRDdt2TrmxgDKOBme+5dWjQL0W8QnabJFM01waW9R1fttx
19kDBTgphSAYiFOXRcJEjH8bvZFu43ytYa5gCm7CwSsM2sISwNt9sB9RwsBiImoqNlT4rtOo2vt5
5cKSHccYv9+u3yF1rMNkIHDypzz/+YEUggild4tvNh2f2i2eK/2e3d848yYmQX0IT/F8HGet5u6d
bNI44UNwA588utGFmY3FjgfVx3Dcw2Rf/3pJ8ykI/kChJU2BIsxSzhqK+/VnlhJxht9zql/XapBS
IidWZ8YJrEjmv4zT/7xS0+4QKLjGt/G5uFHWQOI0AHd4ke7ZmD/y7Mh62Nm1pJ2RparuNpPB8MMy
0Xbf5N2ruFsYz9kp8I3j+GNl/gP/5xX+1vi6Gy2EkcA521fMvJAhpnTkQz5n6/tgzddvoNVkR249
tZXvH5qGrCysR7dM5EBNaJ80CHJXQ3WPPlUTrFQB8Mqlo+RWeJ10BHhEyx2gPjZTd7lmqIEctDdw
W00nEGqFmXCtlJvLCkNiWPc1MmUsBR/jkhVI/Aj3/2LMsbb1+edU0csR2Qz3NbzEOXm08gAPecgD
6QHXHJLzOViZTALz248aCzQdq74n+9leRPf2lv6ashDoHYU9OVR/t3eIppw2jtt1ON1z1bn1Z7no
mdZ1/wzMHAjeRZVHk3Ri77WGesq4PqRYWo13nLCVoe24d0RPyYu2qij9WupMMZAc4tFAe3ANwRip
xXfHAIPj/o7jrrQGnphg1Czf4x1jhTiqhGBhnG0sJdcZ9Z7p69W3HM2xk/4CH3RF2P2jLaNo2bBx
9/XfSsklE0Wp4zhptyqp1fIUdwGJQV8YeFqvIyuGnyZp4JbDvZ7ucNWJAgfjobIdU+5ETtLQF0Cx
IzD026M/s9rs+fksyreHTF8YLZUJqVf4Cc2j55UJVPkbQ8+h0kSEfgEjFI3C1LqvsxjUs2Si3Hj0
9d0CZRAnHBoCn0qo3rV8pRSLVhutdlw9MxU5CWVzEHwniaWhBYjhHhoGlhh/uYHsBYubDBRes/Hs
Lmqeck+rMUWayqqxTYVmBWfsUV2O7r4pQSY4xb9QIPDSniNjP/L2/tGsKMBtlmcdu2CD38eXPa/o
AIcLh7X2GR8n5K38ltcBfZ4YUbbkPWbRuGyewtSbp0g3BZIuOTux4eMGxqwrMrx93oR6HBOac+eT
Sj1PiGOwMdwV6Pg9MYwtlNK1sxaH7tJLf2kL3RN2pqTtctDdtG/1EMhD7bNxoj9YokXsxwFwAudV
451uGglRYxYgRpoDyJEAZMF44WuPZ2/KBGYNyjS+qCmCpnuZLmA6sQGdlnpiUSftvAqXfbPvpZmK
vOSj56jeNUKFOh7nDq2ahDS+fF3dLD1YuOzkQzHBoa3kVxtbMMBdCpYD+7Gf6G7cHZqer+Cjx4E9
//wqarGVown30iHbVGlHwuGo7TLP+nbNxM0mBRHta70bwwz6mgmCVvhMoaKGZG6NLCNDxj/IYr7P
3psULyAINCBJUT9esANgspbjTa+BEaUW161/1CH80JN5LU75Poz9F06TbtHtc5c0WIuNjdHen62n
/60mvXsN4Gzlwf0zqAw14numDADvZ8/xIOdiNcxEoRZ5llbtsrgoGMBhH6H2ke8eA3tUBthKUyGn
i4ZYnGmeaGHy5HB1SOfBJe0e/FA+5KnQyY/l/ZRsr+Wnx4/VFz9EJ8J0BWYPjwFrL7M/+x2P7KE5
dWt3NkB1K6/OzrMBsPU3bhMRLrE3p0qIjyZFsHFP+ZAqxZPPTvNrE1W6vpTZ5CuiqtLcF6mlrmW1
anKwTLKqpzlWMVnDtHE4twby8mkjzOYeassaQ0GmLpiyR33uTS82+coIsnOzkl4EZCzkdlBJItun
BWfOojo9OXmrcuYFsvALXPRWCqhvr2DltRVd2m/ad098zYzZCwGDzOokL0uKbWo+Vu3C/muD/Pq4
yWJK6kFKSlUM7c8ncdT+lTPjw2ePMf22CsJYgPJ3gK5aoNFBaiv2dVC61+Ja7FjgM/x0y8FU9vU3
2t6ryciiTkh4WQJ5Xg+NzQ7p/HvcnCi28lQLNUc/G2ssiH9z7ibdewRffZa5F1sRZ1Zb59UNrw+Z
Apm52FB/lku9B1byBFglhczS5PVbaSmO302e2i+z+iCgUATnmqKzLHlMidye5KOx9+EZFQ+smT3F
jtbuS6gpFa9SLdYJHzXAcaRfbnXK9U4ss0dWGI6sH2MqUoQLHP1uxqxHAIqgqRCOiBDpmqGyAfRb
TCM1Mi4w0GZ/kjrrJDfXbMYN+CNuIxOKLIGnwM0KJvy9s0rJ9E4fSdUIBrUEl/WR6kOj66Inr6q2
yff7eQ/pQLPEbTAY3JcuQhRX6Vqw9/N1Uqs+e+R1hNhXVHDsIR5RCGdEXQ7hrwDZjujXWiedNc9g
Dj8KBbs3GVTt2w2N0OIVS90l1Wlr17Ngg6D5j3R67OHtxYmHG+a94+3Wsl85Y6XsqEhcDzZjLPZX
A3EhJ4SgMdvILGFtRBsqF4g02YP/vHPRsaB7np0s5PPxwt1MmCAZFEkl7xzCUiX67VhcNTyADaEQ
3B+dE7dqAu3aPXAfKp3FBA28b3Ir1RcTTtvnqXwwOzR8bKMF7V+JEouKThPlHBTUTTyIIOT6zOAe
RlvCUIHNgoS2cWP/ERQhs8/W+PxBZCaLdBB2+Xr+5wEopRzZAQzR62wPwJu5huciMFS8Cj8dzLv+
Ma8epjpP6ftCsXzglUNx4/AzTALBye55m/ho6JWv+x7eTsh1npp4uxePWR5cvFUIqEfTrmlOVzHF
eM1IhP2cuOjfYtxa385C2HcTy2HAD+OKKsX93SnqHJfY+8POTI+CA0iO/gsJywO2BWn2C49HoeTB
p5etQeEpHn85qPXo+YXZBC5WjEevP5KBg0iTdCAtCD6ey/0sJVYmOprgVkTKOFBksQr8aYpzX+Hb
dIX1F9Ygk0wcw916f0DW+dIukrdqdNKu8BDMHgBEIqdtSOn0F2lD994EqTZ7TNungCx6Sr+3fEp3
7J9UKlgokdDAK9AUxAq1GfwjIEAAI7rPcPblm3wTbxyyGW87aQLm9sCUXUr3pCzt9fldv+T6ZgPU
PHL+CcBY6NvEGW/Uc+NEozIiE4EKCi04SOHICYDzMp/4RLlcHtE3MixpIxmpLxanKmYMo7gPRbsg
5xc2iHqfJy9dSzJ2597E3aMILSq5oMlkESBi6G51Jm7O17GpszlQtKbDwYZBeSr7vHcI+d5iu9ng
kSJqJVvd81Y1Br4lV/6A1k2JR/ROkdJvGQIXjRoBQJJ0uaDNBO30NAlQ6I3EOq6nyO5RQT6K8Sva
ZE/o/+E1ThpxJNPQkaEPas3TCWWwhwWRQ+sSgWV8398IvYKUsDpb9mjEsWAPMvrEhBOue3XMH1zn
qhJWq/xBGOyR2/trQvt9nMtvmMK0ZASiukf4Wg6DZFyrUlhIpiiwhksiwnaX0LwtxgVLS3GeYwsb
ByXAqtHzPdJ69Q8gkRc2n6evF0xiwlJN9wSoHWXXl3hA/4yYtmGdc8VvjuW/dSnjK676rceHRfwj
sd0tIdNOxM+H8J/3k5k56U9o2yo5vLYyN6LwW4ZMkSs2gI3EBFxrHGPIFYRIzoLGYb4lOd2W5tpa
ZlfjHdtq8qszTfN5vnhQehsmGsyyjOrUugVz3XTAoMdIvLTyYf720oDnK0cGY5nNBjjv+ndPYp5p
oe9FtOAsf/s8OV0uYwVHvGsgdhavbZ17DiH4PPzUBqMqlara/y2Pkc6+iSCAwVhKgSHjWIbuLdRL
vqxQaKqcXHI8CVJ6rGsqhjU5h6gXhytjlRwt6JbhvlVHFqfe3Z7KMD/Hqnn8ECtCAx3FjpprbkDd
O714a8xaZh+Eog43cAbOgzh4wp4+0/StBV/HVIq4fIyZRGSJbIQ7A/1IONyXneb2X9H38lCEAU/2
BIcRBD/T6Mds8GA5UJzRGyp7Tl86IypzAY3qDwd+TDSspEjZ6y6oALo8xiaNgt7y99BhHFCQ4lvL
+x2F7KMnd0Ihv9WdTYbbF37IQyKD/MvH1VqYoOsFsA/LKo+RjsZg5uK0H/1C+4WxFavv5tLGjvkI
CvkTfWRGrgqRAo+0tNnrmaOEE9ciwzYuXt8jCzb9VGI0WE6cq66wP/Wnz4AlOmQEX9Hl9k9Oua1+
2hdKHu0fwHiEcUxyqUndsFjY9zCWBocSI4PTQfMDwpdLkmzPBBgbohkEJCo94U/gTZ9n9JGfjPb+
mDzgvr+T2JCIvEvOnU2AtUKWQVRGOevJcQ7XQAiEVP7O5+K2bMOQObToj5JukSVr5Qh1efWoKt8M
gAzhezQ5O6lI5QVwAa1Go4XKDcX3hOEyvo7ZmR1AD2V0rzGuumlrjWKvneIv31jm3KPB6vO1zp6k
mziOEVZjyOeBXx1wt/NGUQ18huhJ5LF/cmmlBBciCPEBJBVrzv+EpaIRZIj/rD4sziMAd670U13z
ii5gozp4r4NpTLPi5Lx7KFMPYrRyPewB4bxxytcaUuzleZy/ZawJc574nXO5m1IeO/XkdC6JUs8r
kw6RJ0bq7Tkzjcb1ahc4dtuF/urkVEN94A9At9jVJrB1bg2Ol5cYqiJqs0nwczo7igNjv4Bmqjq9
tIijeyK39NTHv7BPB++b7pPCZ66GLNfjNd7yVCgk/wGDZTHEdLvzjIpL+2YsV2zTq9vgKmOJkLKB
1Gu5tfoRrpeIhxH3VwBBnpo+i0rVvSQpedijQ3rNEozDhXO+Thdb8X4LoRAxTKdikas7FeMQqkdF
U8OoBQf/qS9aCLX7+f1LFA1oAWLICtpJZyAZ/fLrm9z3IF7doG9kRx4TWLeys7/qaXhYPYAEjXmu
du7occdX/p+YbA1SpBQO6hamxH2y7pRI8K7NJwBZikgmy/7hHrKtifI+m1OxbHnuKcv4evp17nzZ
YcsCGy8sAepufPgQkH/RO6MuaoC/yGUuZj6snFQuAXwaQBcCO7xOEiCxtTDNBUo2wfv+QCrGhH3m
Oeegi58K+DRH9wqySDm8WAejG4rmmwC72Ytw4bqiJaGZ9QK+SiD87IFm9MrVYCeyKoQcpwncTTPg
Asas0xIs//1RBHaWeRo3cJBUYXTjBGbsdtgM2/jIgc2PSle2SJDGoDD0NwT+UrycgO0cCxrOaKRb
juI7/A+dJOENm66L2ux6ltCHh9pxsyl7DRJaAOoaOAdiGhxKFf0rYdGn+PKcU29J0zsTVg5DErjX
FPTMau2J/Gz+hgcYBWijhX29cNrDIAHd15zNS1pRbHG93mFK3KE3d8nUv7VlAO9F1zuPkXXIuh/d
+7O2agjLZqx8AstLFFxKCJPgkcElDu4A6LU0ONwRW5nMT3Q7MPD32ummkEw/wcs6pGHeok8H0Li8
sHxAGyWyD/oF8p98eZ6WUJOcJVlzI/WECttW+GM0Y49OWyKnKupgBV0R78dMvyj++NIUdewdb5la
yniUOmCqt8P54kubG+jg3AnXrbI24z/y6MnUAEVrI40Lwvefgr+1fT7/OYcg8EkfaxW90wqb8lAu
vIEUB3aFh8quapbSYZUpjX4Onk4mpQ+KEu7hNGNJYtX1+wAgA1gUrrsU3PTr32k53mZcowKxF+lF
dNaL7pYUDogCkEtT0lBiBynMDzvhC570wCeq+rwZnQaVzKFxaayh33P/+53rh+K/2EMvVbxNzaeZ
I3DjcETZhVTwCsGFPIEeVnIqNWBJSYulY9tMrBdyfFVPCzFKl/0SkZChOKuY8ZaICio06mrvEx/j
NMQ5bk5M+08/JbBar3lLiLPF6piqO+dnCZCOGnna+sSCz5Va49FHgqJVuGakiaSsiKlB44qTKttg
FH3ylvw4gNWRnXvjWdvzSpd3QxLELI0js8Eq194eOQOQcGwzgTy2LtCk5ZnQ3KHCIx9MYUk/gBlW
Rdq5/aCAuJmLs7C99GfqKNEDQfcl93nCz8RMJeLdHUZJ0yvFjVmY+wumcSxGRouY3m44UVa/kTsr
Prepv2J/Fx6O0rN/oAJeXt6Lq057vl/mtUeEYYpjI+Yif45pByPFL3ct898NicdF1uuORA1J70ip
7Ra6so6Ku94hqKSvD0JgiwiUW2enF4mfkI75w/J/OShJUuqIQgEKTWO4yGqincnHwdAMvH1gOcOR
onFb7x6qD2JOlpv6/Au1fSKG37FndIGT7YczsQ66EAR4nddcaaMkfXlLzmRVUwHWJEpwop6pEgzv
/FkCy3sfeXyFu136IFun5W/VBgUMCc/QC6OJ6bflhOoe0bbN+wnyJhGwWwew6E5+eLE6yuGij4dH
tb+NC+o/a4k5/RaE/vwpjCTX358nhVU+twgUDT7UVYnVqpnySteAg99ldNHJe9GvzP6zcA8Ga9Ub
/XgXwqGWCQOibWZFjogR9NJG3zcqHiluYk22IfVVgELig0pI/U2f5pTR9ovDXaYUoPUaPhbwxsw9
0uGk9vFMN1poblfnUEHaVMb2Az5UfaOIpD+dEh34T7Mtbm9TTBgbrTP3BGaJ/uOfoEiJqHWYMK/L
69eh2geWiCEz7UL+t+GBAJSOZ+5dAAUYr20QgFYU0bbqREcALnPkjYhWDjIIiF0BsfvWuf2TV6ja
PFkAyLfdppaM+O9WoVEZ8IT9edk9bw9nfUBSxPrpJY7xqJ+1k1dXHmMMaPSQ9MsQHk9MLqNxEizo
U8a4PTRiBG61FaxA0Qh63+8c3M7lnIO/iAVb77Bme9BK0e/flo8FOzYj8BabZpwwKj/hrI1tiquA
wcESDIYZGogHB5Ark9SiAEIEcrPlkgC527z5X0cnQvgPu0GSS7RebCjHYPQHPHhichN63BvM+Xct
GtZ7DSm+9isxQBhPnLwvLuZjjpKTRipdX6jpxBQ0P/nIyp7AMMjVz61hEuBp5/opD50hXXEvXZ5O
++VMF4dQFtfd7HnFJMkRhXbY7Rw/Uppz6xhE6G6pe52WOjCiL/WqFe6IloEek9pXYepO72mKfRjN
9fmalOhFjsD5C9gL3SVxvk7PRiq8F4qGQ4MabBrYN0jiPh4AUrhPjNWmI2PJ+GDFYNJ9ufHSYg62
EtFI7L2RO1RyAQhWO6xtGl9FkVZKcXCb4Tx5uz8ng9cNfPMSXf3oub2NevK+GU0M14DGxbNUPVWz
w/BBIEKUIfU1DMmf3cOHfZhEYMX/EG3PVSuCre4OBe4CsQw7kdVuNMXR1YBXgqNZLN3mYomJ5Lg6
3lP/3MQ/nAcBM9ccEaJd2ObZ8yiCXcKeTgS81PngSieOwNbGM3nGI/cgdrvUqSxg/FB0utmEF8Yi
FerJ59AKkOva6NKGMdK6LNSyrZSrI8s8SoxJKO4QeC9D+brXcfrb6Bm1dlmHp/U1RbMxOcN1phfb
o3gcYPwtImp27XMMn9RzCbi+hAx5C9v//yOzRN7AsfvkPEnptsIMCYxE55VoTrTzvoT0ck1/AAEI
j0y9ElhY2mC7dJD6BzKJ18F3ueyOUBHSJ7ek0bu+O5Fl6vR0rh4qWh1cuZ8lVKAfhuI6KSRDyxOk
wjx3b5ZjEwrf8QZGZSm47JXcUtmy7yhjyyypkmlVMR3EovMFnZ3R1U4oYF0JmeRhUpCIUetfKU/Q
LTJ7zJHG+/9FaWse2+jX9BNf5Wu6C7l9LmLv4S5yu0b3dAxgWSbP59EC/JiGQ/YH8czjIckrpLC7
JPIU86SiEsDMOvyY6QRPlfZr/EYZ3g2DyLwgqsYkO+0NhOPD0/fUmlRuV00VB+NEPJDqAm7vyzyE
/AAIt7BhcaQ1ksbMpN+JFqbyMJuiOnhyo+XxM8Bh2UDY3CxiywT2BJoMIypw7X9BzDAXMfGViHft
/hcdeazkyMgJ6oOorZZIC7hny1bmQTOGnoFigVlJ/JSwg9gnXYOML++euOg17q3bVmQIFduQZDg5
D06L9foCsYlvHQgDypzKc+5A9tMCobhrt+l7BylQlM7lACbiAaPishxVpbNGPYDongvBef/cN684
uG7pIQaHd/VOZ296xQM5rKNKvTqdikR/+kWPeONY6VkPtlEW2JfaYbCFYbHBpGwIu3TTsMdyYqZ0
99keMvPuzuClechhyEIzVJGPRRtEciMk45vAyurGHfDUYaXWWch8uXTY8N2ShdJ5rGdYejA65v4u
bSK6+0w4B7Qgn7hQKesbDoZxn2SpNvdy0NHC6Kbw36J7dIiC3+qWhHTCp+Mx45ZnBI6XoCPCa5eB
4B3s5xpdGhPPgPGQpopPVG4s5f53NHSxF0ez028yT5jhrGLwx3kgb9JMZ1y2Np5kvvTAwhVHFSmm
WrscONTjyxyqy6dbYPd//wv9nvK44LkCpX7YIls1Aac0naoaPiKlmWETRE3SD30Oh3Y5RbmM80v5
mEbtbZScPVxTA3ilQr1acxQySDODap6UrBnAT7Z42ucVK/SMqWnHFIEOsdVnmFNCbs+FaeavWAEm
wUP4hiJBiGy3Pg1RUXfjrnzmo5yQ5qWm6eBaSRNJcsyA37/u/On3qulCRbYJeXAbdEq/kSIctCbO
FuY5ZnyIhBC7FAxlpiLH85uvFm6JD1aGvMxRaFDy1yuz2/qY9lbWzORm3P0Z95MPvprRYjReoTXD
yQaCefINPQ0iRuc0zox3zU+fdFLExPmmdWravVWp4gtjzTzCOJbIQ04Vzac5XXWeYVixIAGa90xu
Cz3dpigqMWaiJjwmIL1vKpBxBDwgPMw+nkyNhDArpzbIWrjUFxtIb6lFxN9JtSvnNfFKQI+UDajU
iTqAWRiJQg8ua8i5RHZpymBAA6bzA8DSIQLWHq/H2RKJ372HXHhG0fH52LSnb7kKTNCMtBdBgGDq
F8CnT+NBmrfRNYw7QW1bqNZqaZLB0f+HegdJLefzB65P5/kUZNWlbXvDozyw+/vhhfj7xuUjY34E
UoN+e14lYNsK/OzW+JB1rzRUO3z/NkS2DqyjJuRJ3uGJFh2EYiF75FmqiOeJmbQ+jaxBp4UUPwhj
UVv3RBKg4fF9HMmttEHISCzj88/PzbYxBcf3uAgSDjspVKbZk50pmz/ZPfFqXSY1ZYKht+lfgkg1
vNJRVmgCds+wkPnd77b1K+6HoTy8AJlTUMhAtjTXh0TtdIMAzDXoBWhS/bZ9xAt+2NjePyyBV2Xe
IS03DnkzVSvrhP4ISFXGfRJupTSSDNS/kIkvhTTjJUylDWGPRqpMEwiS8FXwswmpqYjfru2ADMQ5
QrcpnLYfYf1QIl0LWl0RpJhpsBrYIAVbGr23CJtPed7TnUTzyX9h4wOPhaaUaxWVDrSWtc7J7uMI
N6v/zKFU6LN1zRlX+OwN9V1tCBaOdnVka9YCCmTBWbdVfd6nd2vcTbJftofh/thUWienVNnbTph4
V3tzlmWATWL8DITNvZNrpJgjVlTvpUYMMQBvCvRpvakuCxCWLlzJoI1WAvLfZdVG+u1pNlw/am0M
TfgjKb4lHw7ZkRbfE9C0PXJgrxK4eezJ/XDwBtIW3Hdy9qExCn4nkoA84HglJ1arhLYqyPAhIYcN
cJQUl38MhAAj2eH6C4ANizuuaw59ZEnXBo6KF6lrowT/ceQ+UwhQZ+25VtS3TWwcEkRBNlqaoykM
0DWzB65Z3zua6XonMgZuM8/ZdlM/KdUYNJYoyFA8+mDUyg91PsdYx8cRrLkQGtgxfNLINRA6HeB1
ljUAItyD4rh5VvCyyYBD4LfVHn4uQ3KBGqCnoRKTRn4+Ttxy5PdWJFDc7vFcryafl7o+3Fp7Q1mm
49zC8mMQ9F0EGocy+ovcsNiPslPpOKpLPJBt4pfMYZ74Noopr8my+XB7Fk73SK+gWwLjMjjjcp36
cPtzdgB5JtOjr+7jfBRuXoxG2KcojpxQo1ArSIV0mH2pg/33zYAM+OEy9UMXZVI3cO3xqln+UDPR
ho/WgbgfNcYoN94NjsqsyyHEQgbwDkNyfxR11CQsX4+9FURd4K1VaPKt9hIKnRiaO9cju0z2bcsX
d675Z4ZPM+3mzlJ7uXAV6SLH4kMWqZBK9alDw75E+zOk8hh4lWXD17S/9fcqizrjjvzEtETxfwyQ
6C9WUHMJ1aAcarrXUDAN69hNI+zTY5ShpyUQeVnTArIOjtsQ8vUOMhdQ9WFrXPL9uUhrjWKXUkHx
OLVMrrxflxIrk24BQtvw5cYBpVQMJi1PbL8yS+FjtupTcqUg8BjocmntwDsmd6bsl+o9rPqWhyKF
bU8XOeAQx4PJsnG2W3/uAFJWGPcPr52tgwrRfwUi3NGIwCaPWLrlROTJ1ELKwO7E91N3NNs9Gpxf
hucXrue+zDqjsJnsD0yFRMSeJvja8keTIjuknM8Vl8L3OSUQGn9BbjBIOGdeDNzuQb1JCmch3aiY
I+VEc3Du+jvEGuaHx3RX50Q7TPsPplT3h1AHjn3GeavEORQLQm8XKwZij+RTX4gYUnlvvcZ58znX
mOav4QKGEpsF03KXLKhEId+M+uUx3rbTmA9GLbRlCShmpkGw9XOub/icw5ePhav8Ff3+5giI2J0c
2WIwfHpCZjNVH6iQrBOJ4kgRvKafdF5/Hr5G75xiQQjU0UNEaKWJRwQ+oDOeFbLLpHLoo7gPfBoH
FpsElJrcPaSaIq3j7qNpIuFVcqu2mrbjSyzyAIR4Dy5aJb3kh8xqakETuxeSRQ0TJrLL42Ue6gV1
xwjyTJ9CKd/7KUqicmpBviFxaLxW0FOhgavrkclgqNWsC/aAZimFEG78ssvzJBniL+FhVWIJflDK
Lm/UWGE3f4WkeFLYqwmGlGlgVkfXZWeohr2C3ByxO3X386Wvzns8HCcizvJViVSFFD9RxJhdlx48
IB9Zin2Z09MesujXgqCZey1I0gtcOU0tGKwQno7JRVqKAU5GvSPCLXgoGJqujDDHE0DHZyCFjZAs
/9mKiyCIcVCFlHxrCz9wzwozSxYHBEyeBoknWxh8pNHUhGkm2OY/25QAxHP22Wdt6+n5u3uCGPPm
9ih3v38+rN0kiWtX+XfO08nu5Tg7ha8V/18S9BeKB5+SUhDQz7rQ+EfxnVBUPA3iaUjFLHnHkATX
DUqTxgc+0apwxYLwh0FDfjAlT4CvW+eZhWfBjRVKz9lDp3PLG2fY0nAV5/+4qTX/QCmOjxn/zAht
NUVaIvn4npZkzxNn/fiAxj4EV9jpfeNEMujMlcR9zlU2g9RIyU24sVsZVsh2FNe3JwPH24BI+qcW
P4wwnENvzNea+Djwe+qT2+sFagEfd3O4m2Wp25ZlF4UwQCm3pxZpJe9oiE7GgKyr5dWHo9rvXIUQ
F+WFT4D09Le0j3g+dX/j0LjW9MQrcKu8jNTXFFw/PLTelgNVaFmsfDpHenC6dKMzXYbZNS6ROXDa
YeYS8wz2okqn7NhQZiJ9DPA8122lT8Y7M8ShzFDF78EsUqgfRaH5Wc9jhcv3eOhptn4eum2D0/2J
3p+aZm3Eru//7fzNr11UPVbJVYubSP01RZ2LkvTwRbP2C2lGW3w6ObQiwAVm5EVhbtLiicvM0o9I
mL0id42VOy+ZQNMO73w8O8QVSKciYZO26nOgPpGWrbCEjlAzWHHAOtNCePGt27cFasvny+ZZDw0R
dBqVph/JO8T77iSTL3Pov97w7iXMvScvM6dVBlxSFzzTranSPi2bkRpsfCYyfxPoxOi2LhLDenMk
2fJ3n3aaY50Mb+phi4sOQZz9bYqLu60884jUznP+/LsleQTPdGLe138n7WjzQksns1UiGq/EIyIs
vBx6fl4hOPaDiRraOsgjZzuPUvF0vVivYM3UiakMf5z2rNf30YA60jKVrH2JX5xK2kZj9QitWLI8
NOqXxGNTJQygd7hBZXG7t2w/AwaS3RhTLQQeDMS3Le1EjE1GfNBnIkm4HNeRmVZwRMyu/e9nPucS
0MwzaF68gcvSq62BXYUhcCsqIHV/6hnGOo6P5pJqkg1TC97wW5bvlx7YI4k2WdsrZt7KQi0AbXKe
szSbGasiLjHd++uRdSxowm+yEcjDIaDpHCcM5Y94H1YH3HuUCIFJ92FatXpElMp/MZPLo/eIxDiv
5Cy14xDrM0K9C/dazTLf61sZIX1qrEj3l7gn+0N/4hKuFJRPWmG8Da8cggbOsj8QfA3tpEttO6vt
zyIDjdVDI0JzdpTl352v/abLvgWBCX88bHIXRrX/mIBSszlW/RLFhXGO1SJiNn03CaBuSJLpXSGs
YWRg5eoRmERrFMq27gIuBQPC6svOE69l71W9eTRCjDC2AS9FFjR4+hjo+7Fbe/2wujKaXNz8zHZT
nWPLGy9ZvA6UWuNkLV8pMgOq+zgq4HpAnVJOhAYTgWokKeMEQ6DYSzcJ5TqbvDmRl6FyG7qBMyjs
IxH47oN6/1KnivVWU0TZUfz62FR5UdYeyF2TB7SKItNpdW8KXPnwC5PInbxYHrzRwrcxhuKImbTr
FN0q0qEXXLklJumBQfZhmomui02B11YTVEDoMq1xu6CSDzhdslMxELqT+1vL/JGNohz78lu1jwCs
rxdD58ZgkT296SabiTK9uuR38iZyA7IxEovzq9nmVnhhr0o/fMn0KLuNerQhal4xmQkbYUhedWYR
0/dNhDY31p3/R5cORTN9IIluKVKMri20iipLQDl32xJluppII2gvIdYNEDztjDvQlwN24IKD5FNy
NBdC7zSZkHEyYi8JqAgUXMTypgdnxZvtmLd//4okB7ZJ+orUD/tUqHIICpiprWndsOMBPRsd14AT
oBH+I+R2QwXRWYs5BONHNe0lpeq4C5PlukrYCzHnHYkoeKzdKIlRIpC8AtZaODmZ5S3WsGPsXqp5
uBE4weeD0mUapsWi0DMCk1jNKb1B9drFELhKBbYHtai/EigETIwo0ct/xOthjOdx3pZqhL/g3MRE
//d+rS/Y83yBjla6XzhWjoIAOVWUBLd8eB9X6taraPL/wXh0WWHL2T5D99KFnkI6vVrdY96iinOe
XuHglqYDPPsQTncdF1f+6o1bUTwIyqbdUgZtbZVK/JMYckdjdgIrIW+BRIxDF3GLai4Tdbn+SiCS
Pe2TTdPx+OAQKjvSqoLhIlmmnUKxPIXh8KgBpNIChhvdE7Fmtur3LBAfWajhtjettRZKSfU+UuzT
OzQrar4MZivOzTFkxGgC/LxhUOVFEJJduooYWm02A+uohDve+bq4D652yuTxSE4aznW1B+CUmtSD
ZorA1h5D75U7BR3PA9RgIFM/tZaZXPZeGxNGtMT4bB/plSO82DrLVwzMkr5IQpltJlr7SQXW619o
BZp0ETIukxxPoiWUXScDLeV7kzrlrGFNLhbtDbRi5ntYAbeU4SRQ5jihfAjflnspkNVkoNLN9eia
lTQHdrh1t8tKX41gRYqTkM/x1PWHdFFf5I7oXoCDJNQIqwJKdOT5DTMNThE+B4rwWIbJVJPGUnAY
9A5fz5685VnYyJDiNbA0INMgF4XuJGaKXkG9/DeqDWFrXN7lY/GMzPsBPwavONGwPgiINkFKpYKs
qki6NACuZnYo7dpiA3cOh9wy+7WNDyUSje77KKcPRhR7CXvvOz78MAfCfiaW7G7+AeAU56aYS3gP
m0/eolOHkaUyn+Tz9yEWe/5BSfseDdLi70zcQqJffeZY/4wE7ByVdq6ce3kdikJOIHdc9VAjrlDN
nJel/xZ6to7U05Iwcoo+kGKhOfUks1taEXKix+Dv5SeMu/pUU7dXUROXT2gEQFD+ilj1BR5ocHM0
mZs9Ll8d1mmmzvCnrorkPOUuhHAqRhjtHkpYPliHZMieZw1GL6bK5BPtaa+w0evVnA76AasqPoyx
5QcwF0iPEN7nbg8MLXShCk5XCnInmkFlVlLSfmvYRC83Mwy3yLFsICCeOqap7TJJeSTcnYtMvkxF
0mjmfVM1q2E+GdOOyThDRfAkxuESGQntCxTJObZR3Cq0OONOAiprigtmCtS6i6fmug1NEwMBk8g0
KblsQZA5xqBOxDwFGUOQFg2IlVYESgrUdLm+hU/JuB4VVIUtgInGCMVGUoXgN+2YsJHnUeZYFyoU
QR4ZSfn40jqFg8lUn/w+ltbxSDuTTeF4p2hY5ZbnjnupfCd2YbrEKUeDKFixWzrXsmxdEXcYdZmq
Bgn6QULuZOdPcUNdx7irDxAHP/CNkz46i7H6NvQJHgPlTuJJCz47GfnkGbaLFBQft6tHpaMSec5X
Qqm/2S2PPC4PYVCuqX4zHP9pjgh01zCsC9xH5AS4HDERPzny/EadEZ+iEIo6AiGoQ0M/aOMv6Ukd
DJjDrt4Z+IZo7MFDWJfwHMMbXh58pEgpm1xzml148lJhD1jmbgt8dbZSJDtZj3QV4dDC7r+VaC1g
gFZCGvp4MNneh+a7BH1iCKn0S8T1VoHd/F5LvvuWkXfXXdoIWhijSQoCT8ndGTvFs4R+BOyRIG/h
iULn308wk2jetn1lfSRsAlHaTpez7bRGXdEteqrun0pntYo9htN5V0tiZxxsK4a6jpH7rAft0EHL
2/Ljx+WFBPJwbq7+qzf/uyLvuli3n98NCLIjPgD9G4plN4bBf8quHSiIR3uvDHIBPG8FnrzngUgU
LyFlYS6IRKyV4CE81Rno37kjENg1sOzhaUwmJEid5ZFDX9ar0+w4dv7hvND3j/XmBuDigvZ2NQYU
wMpVZvBJ+0vnD3uXMieCOup1qL7ByqR6EVybDpjIeJ9C+xpI8MzPdBu5WjxDEb7BJCnx/eQiOJ9l
asQHwty87y/FQYdFTQOqlxm4USeEd+ZjS01B9Cg+C4ltfLHhhSQ7JbF6ZACP78DCzK7QWl8RIGn3
NLfpDU1vrhSB3Z1DeH4rfTRMnJChbZyCFFDGVRYad8zaNJPH7W1sRSjNS7mM1WJk0s/VPE498lB3
vOBTGQGZ057Y0DRAXBciClxcReKOnJr1JF+5OMoBQ/vG2YZbHqP0GysBJvO6JumvN0BskQaV6tUU
S3lZSJsycY4qmBAvnsk7eGy/yB4v19HNCZ9yD+nTuug6o4Xcsn4opzlxaxaJbLfjRDMUs0GE0JFf
zFu0Au1EpRI8rPJhB4UP0c09Y/UxxjBan88VBcmUuWJx34aNyQd9I+O8QRMlkEE9W0fm7dK2yP8K
XGkLALYLWvJ0kTtK1OSwoQgGbjCqYKmQwQ/mG7yK2D8ukk8QECHFB0yB4sqVoGVO63B6UWeSKQTt
O8qfSH9IJNHTQNjGZmdOKcOapDRUGTMDnUUtvFnNMlpDnCM3GeO/GXKOwTZT+vYB87R/saXI+oKz
mwc+Id5oqYXdIYWnd0Vli0KwEZNDAEGQLnpIK3SVoAGfJuptd+Fy9Ne4JE8CLgiNTYffUxspuFkb
2c1ZIm2o8MhShnih6w0+tx/8J0nCBy2nm2IssIEZ9wkIQl48/7+jooaqgIHFVCUp59eQy0QBeRbQ
noEtFgXpdIgn+niznRiMC0HV2T8eTS+77EHJOu1vZLC/GErGojqTfctnAxuN6SRIAWODtrbDVtxq
qaBsjTReWX2Yhsv1TNdymRFFDZad8Ag/mT88x9gj75jFYOv6JYVjFAUHXUi+QBMjGdu9fLptNus7
FROg32hrQenugOoWaY93LpOW2ZmgXA5HjCwUoZJoUy8zI+J+D9KkQYn+awVdwSJPsz0j2y+EAYm0
2URoxEtnKkVJZWowy0VTiSPvw+dh4/rKD7tP+SWwSTyFHFpQvVq4KxA10sH1zTOXvivMRZomVuT9
5ZtncLo22Z9vriNY/FgTvcYQwnjor9zgtopPTw7nut6pgT2TNKbl5Az3JgQVY66J2S3LOjFMb6Wm
owUgAtJLs6TxUHgLXVxzXSsz7l0qUEzFkNJ2iBgV0cmilehvVC9qEAtqG79texpn3KVqbzvDg5EP
Qv5DEQ7lv2yp0g5PNzN+0Tsm0zYoQwPrJ+0HO7VOST2V8uI0b1fUDN50YQjD/zIEs5QTlxkRvVk3
URggCJCbZbrg8wk8ignEfq/K6ztd8R9MwZXFD9JYelwLS/GiosqXWmgLM1P49rkKkGP1AtG3Gi/U
iplwFLIBBDmSjj+5VRjQgIJcBWXBeLUBxavzZwKKh12vI07Rllj3WAhZH5hijioo0XcUfs+8WpWE
H3P19Xv7pfaMNkqxKqbn8eVi9ApVpost0ag77Olpmy39sUiofh6gQmx3A+jZw+VWAVizGKsegN2Y
FhKYRMPn2/K1seHFtyhBYv7pMXiU/XWW78g+5YR9sfGmAhaWB4gQzEONFilU4CaGzR9lH5JU25WE
CzRNRqlTnvMJz7wEJZ8pCu5ycnXT0QhVJgBW7/IumGHSQ4Ue1corzATqS0H8we9wsUv5vwL5kajs
YK2mJBc8yNk+RmHSYJkQjbyLGK2kdawyh8s+g7X02c4Ryb6LuoL7g3yLCH9OsORU+JssKbN9abGI
JQZhegvNogdWh91AbalGWwfawcY4lckL0YfJEfVLiJNxjFwAgPF+/NGgdojXHAaI7aKFTwW9guW3
z1I+SV6ZoI/jpnr703NTk2vx828kFj2i0N35mEK0OoYNM8WWV/T9cAJTVl8wYiTHXgpxXmPuFzbG
c+m42F5QoHlBFyUeE6JFZ5g1+aka2oTpWOX8p9R3/jOI9wEcmZrDINJq3eGYJuiFvvJG9OxqZ6vg
AtzcfnT7VCYDwPb0QARxXePQE3PVMpExOyRHLAcWVnl647oLR1lEvNmzdNOO04/+vTofnbiykShF
j7cSTicOAyeEnRC5PsDsbJK2auvcuke0JgCj06Nxc9QdNfXHp0eWTHvl1fb8qA1NWyRCXOmFNOHA
/OlHflad0SFmBL/oKDspo+Ukvwyy0Dj3Vt0odCWHeSArB5m6IKI32VIXlKTedvsJflqU9OCoR9GJ
4JeVFNr6BXHB0hbpLgDQFWFq8W8oBBJV99W2LuBtTOcq5SHoT2VIPut3z6CTfaDHBlerI6xgPR3m
pnRtgSC1yeUTu50sR55+4tCZLr7B+w7zSaPv6I4qELXQUadahGar8Z9wraqcjARV3P+/KiUCuYSE
s5YXhRiZpBYJmKAWTpH1ItEE3zPRWP7oIdsYop4+P071P0iEOMefqLAU9EXoJb+lRtemu9yaDl9g
RQnQ8F2hbmqEzRPZ0zRz+MMmXaxgUy/Hu5I/zZf0ethtDWOS7Ooyrn1iWRpuqi3ZXKBTDfkt2vS4
sGs78e3iBzIzTETPdnp5Q6lc1+CXPsJi0MZWBrmJCWVRHEnQuUVjRBbXEg9vjTCSQgWqTF1Onh3w
fduQz7V+fK2ZJhwniT9IJk8nbMqFSLgmNmSi7H5SGAFaYLGHF6UHhPaIZKildQiKovTWWYRKVvlX
li0Rb5jlayLlfq97z0LVac/oXhogIN8Jsqc5YAPe+M4ezo8F16st5s+bmyOlHYmllH1VzabbkLzi
Oh0f0hHY47ZWJtWOUIquwdpOLv4ANOLBFNw3slLvWQ3jabDYW8AXv0O5bqVXhGMzhurt5COqRgXs
Eoc92DN4RnJejbQz+zZr4gnNW+CoUtFGF7ce5v664m7Z8GcPiJzhTZBuX9Zxc0c1+xDpvcsK8c8D
EaLn21NvES2fIaIWr2PwQyN4QCvXNHSlXJKwUg8t39jmoeGA50T3YVF0Aq6MS0IMM11ez+anKiq2
kjN9iff8j7Ifv+T0VRwLxRsB/gpK8X/8XhLOSD2muAWrb+xEEeTnq+SKPKFPq8+prGCgFbj6uY1r
YC+f7LVYyWNrEDGZsZigreZagv9AqYoJeLQYE2b2xmlEn78r6iEz0e7jWR/cGi7eTwxZTKt5WJez
SFaPgl5fCDWpTz9WaeLtZp07Tnd573YfQBMacAJ/n1dkNH1TFUCwJYOIEAJsVWvGWF0XxB09KA/5
NbhGc5gYeXHXsHYsyjSkxZOq0q8EJf+7k7JIkv27loxKK06D+R5DYVpY8bV+SyN79i7JV6HaV7RV
DEcapgiBAr71AJca7lPsTHVqCh47JFg5wsme7a3ref1AUf9k6E1Y08Z8J6fs31geZM0cCx4oF5fG
gUBZOd/7QATZFSJKloqC0IIEgTFTIrlApU9HpeeepUctWUP7u7L0tymYTU/EpW+57zUZodEaj3C8
5cX1KtMpH13ycIZbPCxx0tzrzg7vI5MG4+eP18/nohpcKTiM/PJVWtReSqFbVLCcFaNxXHN7jjxg
h0o7fQ+LylfAmBwMI6Tf2o5+twVR1ehF5wYru68NFUW8i3WhVS2P2znX69eyGiCnKxf7t+gSokfh
s1d3/J/dSh90HP6UjNI0v5QluRNkfyRp3ajvN0EHwI7UatyVqvITeX1rbSOZkBKd+JfxiRbW/9s0
gCKz1tEtDmr1I/4P37xjEwEBgC35AVURdxHdM34A1QQvua576WTicGNqPPahnWGeplFwbCWCqnMF
iT3RQNx8aIg2VyiPKfwDUJtfa+golFAWIWio621ZCA4d/3jfFd/7AmT73RKmDtcx6I5a8iWgeECR
aNKPvStmI46NQ20JFF1JxmP3LfjRhwoZCJjRhRPptmYwrAO6rzbyGKnuVT+6uJVVDPr28UA5ke4F
zQHZ++FgQCY2SJNiWG6lvss+QgPo+DZcEUdMhURqT1oMVk9nIVDpQ37f1l7+3jU1HgkiGT3do1HI
jPWV4C/6ppaNmLcShtdlIYTKXLodc1thBctWgHFrk5w9rG0UWb/Osamjx6ZlrVcnaJBU0rRUXsTR
hmOqgCDAEwnzE50XqSfDJUDHUzXPcUD55JSDIDTXjc2ou1mlczYv6Io3N6NlGDU4aP+5hCw0aQ3o
hnZHzmJFemdrxxdrBzZS8LhoOZYAi17R23cMEv+P7MuSwK9m3O6NUUmcJ64QnhRouiXID3/rOG6F
zO+GvMMYW+E23ZmL+kCm4qJmCqg6cquHtH7Ah23khcDYpFA0dsjU6HMkBFP7PGq0ZhMWJKRIY7Mc
HBlYJ8BLX6NyOKpqms6Uvrcybhz7Q0Xap0uI83dXWcRaO8+bNKCmro8zEtPRBo6709RbqpCBZRuu
PyCgJsWyP78Z/yiFhGpBf9GzwSmVOSFIWpGq1DVTtQMcgg7P4CPS359/U8sSg5V2/MvwvIqsf7+Z
38Kaj8ruQdnOFiGQHbey/dTcr2tOHN4Dva91+b2BWj8KaKWWu22kmprGGLmK1WitcEUV+ZmJMvuQ
/MJCen6Lkbb6ZYGi9xNto3gDzy9+HwK7lm/k0Km54GbdOZ/GBMoWLnwmBKPE0lpScIdiXQgCDZ/e
JLcG2Ag+DWNYJk5rlTXLY8i0RDJcNFUim9dzaktUSHgpWeqhBqKPeLkV6sq1hyTudJr89FQDJO+T
eFIwYrrLu+os6DgDCxpmfmfWOYGjpnYxEetQSpIqJNY8Ff81jAay0juMbECyTOQ8SUEbqA8I0u1c
vHNMKgyTnFYcEZ5l2tSeagylUzqRIgpFyi/zLGFvfA76kk95kGaWLxPAdpC45HDUgNebnNTAVQeN
YbRf1+yFqc3MkN5U2mTzp8b6zZkmPxLy/7mWhyQWc5P68j3SSxwSQVxp7ot7Z5xI5RIJk+Jc31pX
b/uSuf5T7I7azqPau+oODD7azvgEznBF2VtYFSRU3cobFKouiyjlyzUDbDTQuExYMgn4vVtmCm/c
gj8VGCQO43gGHrkrAZTu2UOwWlEw4FoMTuVLqr/UNem01AZ9Tu76X7UGOsAXRot15Wxq2qFQp8sL
WQx4YAib7rJpL3+Y3r5dnZyeuAaiSx25X27kuaN+/yyRvX+1xM4EJUgdVbj8Xh0kq5B1Gti5wzBx
KVsotBXoMiMOJZNOwr7uBckD8A3FgZFH8o0NGs8NPJire7sHOgwFdbujKX0bRZpAmbeaqfgOQvnM
z8hfS5/b+fbjxDHjWf8wUVYYduPIM1P/i8OYIUNDxBMBsB4PdNNToSSDJ9a+4Nxj2Seuv1f3n4wU
eodUao0mTOVVP0vj7j7vEDOD33sJQQEB+Uj4xOu4/mpucyOtVtRoWeoKBhxAgDq1+NgIknWavRRC
MRHZyW+wKZTXxtrmRi2J/5LV3egBbrjRwlBP5bBklM17bUwKEHdq278hiGyhW/UatSS00sVaeHYH
/XXEtUmVGlVBVPvk3CZY+0V5PXVXALpuhPB0BJZblwg6c+zXSpQJfdb6YxiC8AE6Ctlv2kNPPPUm
5G1UGG0l47Fan1f7PxM1/eT3uNwPoZkWEAmwGGpBDwmgPd8XbiMfYrZtZF8PWqd+8Tq8qcB84NmZ
RJPeRZlL+4/V50s0YG5MLBJduNVfx5V5AJYtPhtrrU+ai8HR9uYjmAXYXHEYAcDmxHKYa4fe90pf
AruDsmZlLig6Kde0oHE8yKWn/356b4ogVaL8icUGQVpHmldkBnw0M7W8HyLbJnWeqghaFLFyBeLQ
bPPGki/uvyNiDZjY+dBX5A2q3w5vOs00Dlba0/5wcRwaAb1P4UnRNmGobLa+axXo570JlKifHdfq
vpIRW3oDx4mAPWe2TBV32TAZsVhy0Dc7JQiGNo8qeX2YoHMG/nRv55GXLxgeGm6WMkOe1IyNBMDk
CuM7PQwov1naZbPRB0/QbNI26G/aZ4sQmz0j6I+tgDkouyBoAKtmQ9fPt2tqQZR1yuHlETBUhpFv
UXI3B9lRWy931WOwOOmBIaA8Mrygg9cKW8hZ5ySEi3x6NEFrp2nG1tBSkLc45YKBZdTpOl93zOHZ
+LaCeuglBkrOifrZGRvwNfjFD0QZQMxAzALM0jIGbns+1OlYk6tJLfK4idjYPgp8czs+YvLLc1xN
p3pWU9az5fRsamLo4+uqIVGoZQW6bcpoR1B8WyWheo6UIBcPFRV2dK+lsNj3rcaqJmlm7BQp+blV
R9GeYwB2HADAIl4G9OUwSWkWMEwUI/kHOabCOX/ffGxHY4ghTwsTWVZWxM2qRzKQ0RVUocXvtjtB
/644giONMd943pHiBGCuyBJGPJ8u3Az/lfdz1j0AAHep91sA+hHRLE/McSVRJNC4ROk+M9w6ni1N
39iHcBsklschpL7xCS1/xdMh1yuu3o2mxuwkx6zd2fl2lBwp0GpSVsbgtcPlbJjKKmS3m8Qe5oAl
CNWWP8WP5vcaRO4X/BFnWHaXT5qDXNvoJVlyqxPbWQXMfQz8rm6qjP+FSdmnCZdBPhBt90/WKDOu
GQjlPA+4JdPrvglb0Paq3Dsj8XhTILAIqx8c2f9FHmxnpeW6O8IbBap5W9y2qKa5LBLlZbAmRF9b
Q+HDGQx/EQPT9sj5cNOb72K6OUt5pioXOXJnzvUK/ZPimbtue9KQYAiIvgALp8BxN8XqZPBgtO2T
93wlWa8WtaGKEWx/1X/7mvpT5O+8QnwOP+K7qDLOPdNcPBEUb3PiEx7puk5DS/6NYUHTnhqK2K3v
1WtiQsEhLmlrnLb4UoA8rDJUgVcQtJMW56zmqX2oAR0A/a87Nzjz+Yq7sOKCIqMeiii5vQdkQBmf
+GdDuKHLpScHZYMi1q0ZfJlqk6Iksl8IBKqsDfI5zRdNItmGUvFVykfrbSrOJASZrZ3K0lMiMgPo
UEvDRa2WBjpjTwfqEHFvL6Mhf4LI08UV5tFlmFcgb1EmLOzZuVDqLOlDp7xu/a+MbW9LgsjUQJX+
kVj37qGTBbFykcRUIQXE/TCGUHyMZqVt5MXOFFVI51MHeM/geE6QX6lqVo4+JxBsLi9FcVuY/eUa
06kAJ8qWKPTm+BPybIVrY5DtJL12jQX7DW2AATYJGQhGLCyOo0Q3MEsbC9R7tiv2eYonzw2bm6at
5GNnHHBSI+mazYanSG2s6LpQnwtfs/crjUtNKG+E/4U0uhrsjNBUMCgsPAXtMLXFlvpzXjiQCSRR
0EHXPq9IIJJ2oXqCK1SJcOh3z96VbBV0qJtclBcNl/PEsmzyhbEy1VUkme969Boi9hdJ6HZdWlMz
oQRD0dlJ7OZ+zUcFObCmuba4t8ukbVWpE0LEIiESi7XX9vKsC5cjXVuXh1jJ0cOEST8rLFEayOIP
9Aaqvl2FeqlSBxmJiMaQ1RcfgH6VhiVJWt58lKqUbOXk15/nwTtPYtlnfwxZUZrbdgzr6fp3mDWK
NWg3qJgl4LkZWo9+VUNTP+4Oxanp/J7l0Nrpp9olukTqofCYCF6qTDhv7DtILb4OLbxcLcqYvPtv
/EuVlZZv/Q9xdsWlMs3qvXOvG4MZ5HtAnZTxvGmKXKzot0ViIhiUdHWt+iei6LwVbeaKX+VCwJiF
B5wjKxgTp+WVPAMFmZkSvZxGQed9XEAJ3kz7l+8wubYmwMwTYRlYMbQzh2ZYK3Bn6toNxM3mb+ml
FjELM9ODKaeY0mltQFJ49RAMq2DsQ+sZB7VvTfvtODdElUg3KVFwB5i2O+nUyiwPgoxMejwxhUwx
K2q4oc0BDMO3bQH7LD8kmCvXQSg5q9R0PYn54JfroWb2Iqro0jP81Lit+ADtDf5ou6QLcpNf01UL
4ieqcKICMSdktkKrpAkB6Y6yJzgBKXkyiJF+65orVq15T1Fxhzo46HiXrsJdDRYf44fjRB+GoKon
rKWpI7cGZjxx2KXctcklFvkDLWJ194y48LOD4x1cbLkllF2mKzQ78O+XQPAC+VOd7ct7oMl/7ebi
D3P57gRR49qCoF1F9JMf/BJJssjPg56CFRrVlHypmxRRwKqTN+OHrAMNTyo/or5cqHGfW3X0994s
tEOTEjHuqm473+ywonp6IaepuY2KdLbyVV/IOL5zg/XyidLAn3LXkPzoh7b2WKm2wIbGWuJOUx4L
E1QTApdHUTkuzqEglBWo2IRTJIywUUq4xSBjRj0VndIatbZiiFMBoQBG2SpRlOOghLTfFFCxwnSG
ZtG1+NC9vsVWKdhMUqN3kNV2U8ftM3XB7iUf0LiRdAfj3Z4fJMTs1t9cE0wHHm2QcszlDdFDe4/R
bNEVkwc01qqXyw0tSbtg8g8VIHEYpDM9ezRfjGEc2oN6NZdh/J45G5PuwSkHcCgTa8kPE9C0sWkX
xwT8XaHfaNXaMLVzjKCbvKG6sfhC7Y167L2wppVpejVylg1jqSwzBU2c2vldV5dbFW9dFVxSOofR
FHqCwSgjNMpOFf0/xobgSxLP0wX1MgFZS3I3rg+HUtvsvQB9XZMu2Uhx2KaOGBVYAMHkml2Ea335
nlcvfG4NjVwCmPtnBoW0oU+lnDWWR/B3LGM7shLPb84jQCegwGB3qKESjYfPWu8EzW4IosdXdcfn
sSEeG70GOcfLyKVZPUP1sEseogTlisCbMZ3/BY5KdlzSGZe+H1/81TpkV8ZBZoNjnq/qM/79TLjm
Fn5NnQXzC1AxToyKoO3u+L77LzaDX4wtlzxYQStzpPu37S3Qvt/os6k5KyyYXfhCi3bgdrXxi/1N
c+jsQ1uJSGVPnEINyv/drc2Eis9tYKiOSlE78VqOHqRgAa9vsVglz8GXSX62tsI8F1fm6ezBd6eu
aR3HxycTCeEKDkH48GlMw5zbAxwWTw2Y5s2gri9KNzKVw8+o6rhO+yP3NeMdpIXH/eLTXJlHXH/p
XNutmOc+amLE9BlW4bR40sqXZkqIW/2k324LQKWJZKxnyQY/0I5z6up1nvoew2XOETPlNSx64GG/
ZrBlFNJxOozbpIW4jgpitNukaaJUeGxJ6//y//1pfs6B0E1cQb/e46pJG4QVeh6BDLNFVMcjW06f
F+kx50owm2kaX8sk7Rjgzwha1f15c9TxQafdC0tekiICr3z0HU+uygdH4J9q0pEoP+hpuz4zTD7N
zNG/IfzTi1fEV2PXURVC/dUaxs96Wo7h/SCNDwQUCwwSEJ43t/mS2yZ7UO6/WbreQcwrueGhpU6Z
wmajSQiY2g+f575SC0fps2fx5Nc+X78Jvy8Kba7qYvudgaPsT87QqZ3OB1BugqbtBQUyHEF2m2r3
u1+YK/DEAnHyx5nVMO7v2zdxj+CXDomMQTUxn2a+39y6VCFYBBOyBrcKIkWcEwgCVjcQHMM9a+lL
co++U541rz7OfiqmYmUQn7+s5tnvAvry+OqTVhjl7L26BRKH+SLW+IXhFPW8l/Y6/RkwxKHZujkf
fGI92dHiwDGZpNU9Bf+6RPrrgbcBXnC+tGTi/3DFfuykHspfUp2g1op3l4bgmk/EL0tzuSQIRAJd
pbIyy2E4RN3drJJCy4LQrIF/8w3VkVuIDW/LbPVRAvmYZYYJNFFAgUdY9TmxOwV+khVLF2dvoqRP
7b470ewwd1az0SVKDQcMNqjCI2vN+QHzvWwsBR8g4de0v2wISYRA9SN+/q7irqvJhz7meC+EKesa
+VLt0Sb4NECCrEEBNleaF3B0bOpsBuxCcRjO1wubDG6exnmaSjqtjtWObi0JFSF1S8jsc92MQFu+
ss32my8+/Eq5Pid3I/s4aMORONxsGy/Y/JXakrkZ5utxQtmN0uOo5VEWcAuNWxbvCE57GOmAdTTk
c90X89T59y+ebMM3PGZNuGj2qXVLd6wGhkMzVadopym3+Y6e/gc1VaLkNCRIznfbjiAmSsW6B6dQ
6H4f7EaS+VWu0Rjz1i+6MdPAGvsx/dh6+A75kHnyOe1s9/S8FLNGEJjRE6ED/Sd5uL/waWffHyAA
quCnhFaTAelPK+pcxMS8Xj6+3A2cOzbH6nEVdbQRG2r8iCHGuZBJtV0vFyzP6CFN5vtcdcMDbA08
EgwRtZ+x+5uAUtVxSlJH6edh/Y4Wls7lCeSzbREABdaRZ+wTJQJq/YU+IqhqhFIuaO2qndOsuIcF
hwmLN8FzMjZBm5unArPTsGBQ4ZV77SE4AJ7C1AgvPvD8Ce6lJQuK3D8s2zYDXiCj85JxliQ5YN4y
Av9815KnM8yXUF07C8t7jOe3l89rh0jDZs05PtC++H9HTMP6SoWFQN461yNVPV6hmvUFfAe6pzyp
GcNgd/t8tRxbQbITL54AGJviKmVDh4gHVJlUmzSOWNKy5LDDbprUEw7oc9Q1AsnJcNboD6wIj9C/
x7MKuCIEMR70nnQD9W07IxcdM+1RosZlh/lw323GvJu7C2M9ggn1v5qpYBWOLtSFQGksG6wOF0xz
zDgJDI/veYeOzFAfMLTGq/tyfsSE3Ffj0fXsC4GCZR/MKCuDbddwTPzQEX/WWqPY0o8W9btF7wER
k5/BD9Vybttxsedda7jpqHyyx5Ez5kx4BLQWtN0N7LmuW0DGlAbL9Zn4OhZCbrV8RLkd3bNg8Oqx
C6haGqmhsVQvQkxAraWDuKd20Dsq3wh5mKg1THStkZ1XKzC+WqEutkH8GimbOuO7wDoVOU3OoeNT
v93SbXwWFKZeE6OTuyI0vIv3AddhViuLt0Rm6J1NILsp71aEX06W/7f4zz15nlqtEuwQc5I3pIdM
TAX1hM4pMOrLH0N/XsCdA4M54pRuY+gxOm4Lkozf2pksb9YsgIt+Nh/2b54Gn+kcL8NwWnlpbdV+
/wyuJMP/OW+7bu9T3vHg11nitxTRuiYvOL93Uq6rDE3vY1K0vfWrS4Cd1v5TnPSoVW++oupLCpPC
DgGSPdl4Y0qpo9BvvrO5agnOq6QWquwESl3wcy9upUxDpIv6ioUSxFGFYENkiU0HIzR4AkWEWi+w
0uCr8GCkKci5GtiWljlo+kXR0dDNl5co/9raAGBc7zknVLcMaRoGAw2cBUA2b77YN17HXpVkm8kl
g1MTBFM3GSg4TtGRsYHqU3m1pwx0XYQ+EtYvVYDMjR4Lw1ornFYuDrgi0GOMjQ6ZTcTHUXw7Sa/6
zKope5Z7Y2HSEyzbspqBZJVnHrnvgyZ0iT4A1RPWHOTh6NTD4qNr/SxXSpYfWxoJgavSOSwYZmMO
IiMQ4kGseP/qg8le4FQs7DWPVMbnFhxxlEeoN0xCdgkhSxxzy+OWxocKIjfhwY15P+QMDuRBraqT
TpU3gcCJmIZRK+FQH1yEH0yOro3uXCwOseHJLU121H4LXNzCn/L+WBJd0rTkQm3+oKdTFL9SgXs6
WU4HdlpNVDa1BqJonV79+xERSW8vErfUDwRnduuDUG5EO87pzGYMqBDVKfi7J7zcPEcRUs5NAYVd
6scpqoqRGuaET3TvmLvnQACr/nNiP//7Rq5eD0DAtVikeY7F6OgzetPD02L1brQp9OmS3qGJwqln
CpN073ihOUV1Lop0Kr7O4fhIcHwzBgtbygn5nDFt7PusNLgkpd3jtzC//BkR+X31Pzd+G+BdFrLU
hed6MH8V/egn0rfB+4169YbGsYeQUodAl4bVukHAu6pOGjhUZNmz4PqS+oye7XBE3GhHVaGFptdt
OkKNkk4FyEL5jeaeULQuFMTbc5Q8O845UaKZM27PkgLwKbLNBZefCoXuNykT7McGS76dRfJhkW40
gK/hdzTZXSWgelXCKK6LV9pxkTVSavsUDNRhmy/UBXZgL7Ll9XH37vS3mOP1ZXRJcK5uEo671fk3
OAIw9d1b79iZkJsYkeT6BXK7LOPE2gNI6g7TLQIyVz96iytp33Ii8tqufaepp200gvi23E8UL3Yc
y5yWCMKZC7FXQ2rKka8WnjC4Ab/dYNJv6qQjOk4UkHwobBSu912h3tsTGr0lym57yRss7O/U5cLp
0CTUGKrF/hAGFLbEg8eq00/8I8ffZMqy1luJfzacad/Im2eIKiBAn5YJllGkJNWKLPOdYBRX6jws
+5tDzEgO6bdr484FqqC1+1bzwjz05hQ4faWc4YSrJG/uTvQto67ruCg1QBv3U6I6e6pW6aj8Kq35
kFGOYdea6uqCqx3p05OqB5npskitUZOndhY7QX3I0BIQuOQExetXaIlglFdbFDs7c3KNPjihY9sv
x8ZexU2E7Z8qxiU0M+KQ4sa+i7qMk0/hV7KD0DzUqs2m6iSaOV5aQeXJGe8bk0LQ/yzQ6xN9Q4jQ
8y0A5a7usykaFeLQxxat4b1KS3qqsMClv9++BTSTYapIFnod8/eGGvQ4yqE6bftiI6ME8scn1Yno
5mc+7u0nPwSv6IMhEw+ENYprQeoQTrfNc6jDbgtMbq3/svAlSRFq6EaznyjmItsMjhV5HJTYxcDA
WOMWb3Yi9eztEHKih6pyPqCW+1fMcYjRIdLUHUSum/aIMcka3stdsvR8ftF32xrThPUNhaR73gAL
I1bqN0Ltsqmiydk3mRWVIdLWmxRj5ChTwelNgpqH+0oMY66a2SHha1qXLkIYqjWq3EhhHtx6uazn
MFe/fhpTE0dtJEV9DC6k4H5BXuMuyezMrBriBGZzpsnlQjwI6hhRJUj/q2e1WyxtxIk3srhtOzkr
rG17NcNKB2PmTdxQMYRRR6WXfG34s+YGOQvHS4TqS6jMTBkBKfTlJ4kZGct2JH+Psqm3p5kjy0Qj
iDJ8CFxU9yLy4eqbZUEdWhjkKm9S+75hXW2wZC5Sc/1k1wYYQCbLihyAGkiI9iMtHgJRSwqBbs54
83O2cQUHKVlJVSgnXiGudm8R8biXWxs76m/ARH7OVOuaYxXHOiSw9LOfzBHO1fE7S985IuGHVwZe
2aw/gAAAy48U2U/0fwklyk6jrqV8p0YYUcel0EXFj2S0kz0Uxbu/dofxXEaeOkFbkoAT2cO3I47d
hLQssxLRKd96YT0syMw50EuudUePC0LI4PlZNq41C60U0bCP4H654fP4KSUTiHUa839xF0tDRnKC
DDDvI90kJJi0mmdIJyP24DSnS4QCLKYp3T25Mrr2/frOGndEF1fToF5n1+l8OMwoJCdKwiCL7ej/
EztItjtVCHH19SjpZelBcHIJ5JU70LLo2TiSfWtRH/haJshUg9cUnSPgpKuLXZ9cnl9vz1tk0lHD
5ShES5xjS0YLKcg+4Ee/4Cjw0siaPy0iloeS7xki8ILjhXXHwD/TI2DQo+KXY90GJybGQGBWtOW6
ggiqXj/GLRdzWr8P4aSzC6E1xW2+rGxwoxLqNJmaESGuiXt4Fb9olhbPIZNEJIHBowMjGIYyECDt
fu7DFqGuaB9V/5VZB5ro3/xkL4joYPd54WHPkFH3apXxnPeLQ2LjlOcFpklmfJGpfYomQtd3fXMC
LGZBtPIFot2UnG7WzzXta55n2ewBcwmy6M0vrFoLd3RnuVUrulRL+al6H1cJKUBVxUWR4OkSbbCE
Aq/Mhf4XLun1hdK4tGdcVuNw+wEdojci1j5yBljtg5OiQUZzVoGT/PyR04fggygOLUhXwBcutjva
rM+gJvRXOJTj0GyxjaOwLS8zLqpIE5CceEU8V9AfsrhyDjqGFukXR3dPhXfHSlbvD7Ic5d3arpo0
vif0s7jlY2c2K/0Aft1HvtSX65FgzAupaP8qwNKcrjV9/lWmFud7FgxLj7FsAh0stkM+J+TxmKL6
FtS0a5L7Ti24FV8kCLWQEMqqNFizJ8jj6jXeln5YoOTDd0cMdfwD3u6GKUphh4RgTPrD1RwIugV8
1/Euy/sbWd3X8gQu9CprIyP+X+5e2NA5jMT7Z9DQ9oISNWr+nHeuhYWO58mLj2IjVWxoYOguBtpW
Qcgx+e8wF0XVdFa0Vx5KCjRipeV7mviy4TT4KT7eExpIUoqN0uPsE+/ev8B6ttXyQnA3AM5JBAcF
k6exZ+8CQI85u0tErHRlXBUiwtVa1JMXBLUDW9w0foKwxa5hiZVrVSlPiWhO+POwTjiMjZS2m6QX
Ebvv6X0GU8HVr9GsBMKERhDj8TJWTj0LTQZ0aoysaaPM/K9fdc7GZLSyP8K0UKWtsc28CuX3fKgn
08l7HQA7SYuv7n984IX907H9jPTAiUJLqnL6JWIgnao1m4SfD3Bgl+Brl7T4HoDqsE5qktREtU2r
nWf38Q2rbhFpHn58jN5e9FMZCxfcWs68dlV4zj2AletPKHKyALu7FBE3lyRNnsKhH35dU4ZUcKvh
7+br/OxDKnUEUJOuju6t8jMZ5DTPjoBwE9zTyqmqZdqBEGbtrFdgoH5syNjFTCVBTZ6qkPkjQ9mQ
b2BjTkjNDse2mLApzufnyg5L8PO47C6lgsS0NNO2XOhRgLVPZxQxqfvZFsOkjhG/mkihNhQ264+O
ZxywdBHuZVY5ipVJsNPTJCZG35VCNRz5wiKdVv8kLQpYkV/6nuVlvpZULSmjPw1HBHsuP2vKY42q
z2Kc0sxUNvNVCW9uZOVRQmS5VEX1KgeUQP8/HZikLf9IO4+FNqa0a4aPl06+wOKBbhS7qxdFxCT6
3sRH6JQ5JDUeCZhJyQV3bDYlHthyay8mCprsWVkX+kz0LWWwhvI57vP77LzzVHr2GkhzdcnbL/iz
jFzJZime1+nX6J6CQkVqgBh0Rta/8Nx0duLBxG/gzgh4s5hNjVQYaZLTXnRiGXF2iZRgDeAnkCs3
9H/Xp/L2Yr5iokL1vKnGd1PwYUcSh7efQQwZo5706blPDQyPaX96zG74fLSctQAGWQCy4cdxEVGp
e6fwd9ZG/gxlm0N0NsXF+QVe3S/Opj7JGAFEP7oklvWYsatYMLhYQczy/Grf4lSoQ1OWPpiL46ax
KNO1Dzs+VoO8YJS77ElAXYX0MRJS7mdb8FWEWqf25XgtSkn04qvuCVU7pGvciKAj8i7RILYVSji2
EjU/PbSFDYXT2UWHmMigQJFuSkEXZhVwxtTKg9GxmigXYNGoqOEyxk27VMJ2teOSSwpfokVf9Ogb
+XmchKRYjE1Gd8ImTZ9sz6BU0pzKQNjITiIdZOAYmmx8rYjqdKIrXgWzDPx8iywO5kZoLik452pQ
WzhsK830Ucx2PzOAwB/rjCx+JGL5r7PhG1LhRbdPL+O4DAwuEMbcxWNlIBSOz1girzRBy2XAFWxQ
OhzelbAUR843H93mED4N7zEhUhjzPqe8+tWKCfjo2SXjmLFvzRG+UIWYUdxO8oF4gwVn6tIciKib
0+E85BDJ52dykily7ADs0pvfbgY4xTnP54o5Q7QyKeRZRLtJXFUD2v4wsSiV/NgVE12aiZzWjvZ6
6ctQNfNg1enp2xyZqDA3s667njMnLyE8DTPJGDu8CxQ7aCmKJ0Zxpr51toAxX6gdFfwsfDJGTN7G
JZu2QfSRN87uppSpbV35wJVfnQrBXcrZ09rc5+QZkfh76Nxqy8kg8GfWEBdoaotlOFyY+EdcahzH
zpT0OoJ8QAsUGJKVYivtsQik9qyJFTA1V04WWn5irpbVbIURhY72Lrx8pdGk19hDKXzHR9YUTx7L
AEocg0VQZz4mqyTfgUObIPXfuGrqujDzpfDVoJL9K+oYHazq0xi6A3USIziF6HWYCTKPUqmB2cSz
tCb7Dvj/3MPznanydRi1M/2vHJOgWWe1fLpOxFCVAz+AFxwCB7L3UVOnJ49CfNBcsLw3xF1G10/6
UVdKf69ZOz6zISvhK+D9uUVkXIZHOm24NHVhij/WnQlCTmBFQctimwjb7yWpii/gDSqMQe+7wEeS
Ayb7faaGcPwg2vZc+vWuQXjKUptTuyRbU3g//fD0vAZVGGjQPDBl/TGeQfwXSKn0/HTwIECoQ1wp
H8lQgn9DEkLIOYjw8ayh1HDidAejaNSwdNPLX0afCLgY1TOBNSyvVdGCC2x7QZRRtbIK2J5wg+VW
iDvyeGyqnT2SKt2YPozJ1LQL3KcSxMkiOppjuz0CIqylVyBo9ALzMu7aHDMNOjGvxi64e+7FcM69
skqjUyANr9cxDPyC3n72wVIYCCuwuYDhJzL1LFWPMfuxpnjZixNK0JyTgsn4d4As7iOo/XPVWLS8
/y58ViWCMdb6UoX2EcKq4tqF5Lw4nReGe7zSHUWTTyO0I+OOFtTpMwGKrWhFld27i1Ou6helI8iV
WIBgVmO+rgJm1VMbNcUJQO+X/nzUnm2cjCS6VYqO/MKAcEcOfohWDCaI6UzpCxVybwTFGCDBNxZB
JYT+oIeG+kzRbrPteBzHWq9/XI7xwBFaclGPiscPqCRO+O3KEeh5h3fiPIwzUPrNDydHlbuQQd5e
NuzpfwYMsr6Pw/zxHky8yeBHHjFgeofSHCMglie2tGYmPa2TNRyVLnJQSrJ1tl6mPvsZ95qAfDKk
l4s1us97NDvKvfzu977mxwXecxmX6uv8SR9/covMyMoiAqteAiozqquWhskE2s3E/Hskt5CEPcLG
UlvGC9Trv2olrV9OPAH5eBIONjl4Nhgg0AfqYonzqHPuowINqF25mICauwslJJwKy/s1+rxKoAYx
wjgUh4EBRbLZacXRGVPRvU7/rDNOMK5tn+HsoNlKwpw33pj60HVjEBizFKjL2N8ApCezWAc1qp9n
niZBfOc4OLykkUJDImoiolEzvbKZrMKUUM9qONxJJcZn6tfOSelQQXUhfUELOlFhSgfJziVogGKj
UD6qMU3qboHZBBou+D4eWwQzydQlwStw1/PLy48d6NXEVtLHnFPuwup3dq0vyDeyiut0I6aQ1euq
LEKr/S9bk7J9YXkU71teS4g4nX9lmiDCQntlhJ5Db43kL8X1fYjDyBFL4KKS/iA60so4wwe/OlmY
LTUvPhjF56X6X+J/VxOu0tQ6NtwhYJBWloOBSlZFmQCUs+9ABAbqb9Y1AU75+H2C4P85Lg1E7C7K
/+BU8g7v0lGbfemk9v7N46MnL8ZKwpqAyx99Y8xkUijG0vlsG8X++tNUgTsKj9DtuysmyakfoS23
q1ZiFXBH6ug+iZTNZnNx0GTVKTgpi+DchhyDPVW5xG5GYQ0v74ex4xYi2L5lHWRZZQVtZPRetZhq
L0yn87fwNoKD5635xO5ehYxZ88anDlKZ5SHKwJxEWKWKNJ7lYbj58e1z9s3YCjN9kR/MRODB+hJe
ilksHYp07wL/3rQxwLBjYX6XwmLDomP8Clc4jYJYdnf2p7uloaZ7VDja6X6/Fv39iwr2n1iQbKHU
bMCKy/XMwt+z1tEUmaEehDF0rA7wWB4C+gIdf3J7NiF7ZJmsxewm+q2IUu7gFKrSb+lVKwlTqsYQ
IA9Qc+NLroeH3L5RIWwmNZyo8VY571I2eebkcnpX/QMbNFZKNQKAlr+a4QedOXLfP5NW2fEsT1Wd
2vWKDdmLk0+0uHFQJ+FZrHLAD0KVSn/fLqT5Rm9PCKJefGQ3MDm3huX76sbfdhUrbutoBJ1/1oS5
Ptxv0sQQktxD8z88f8jg0XbbbKl+NRa8MRob1ZjvN+yNCYsPAfuiZwgIo2dY52jfngezkbhQTopB
KwdiSmKXxG1Z7BzoP0nNtSjZbs+wOXw9qe7JA5cR6HubIwNRmNsiri7dwaE0CEkY9o3rr8uT3GtC
jWGO6yRycmOTNtnvVDqj5W0URFF1uvYl+3VGZpiPORfQlkdUcdT0HfChfYu1IYMRyBGrylzSsYbr
U4NoqekOjVGELgr2mbcJ7pnpI84UUJW0WzhlDfhrhPgaRSlcYuY/boUeN6N+U9Jbs2YK+s6LHdKd
6NoKCczlql0PftFlmu0CNDy5stYlIPjiQNoFceMcAGDzdec4JWUaBOi2Pf5xylJuZPQzUsO2zw/z
C+e0k6k1iUdm1uo6sx1ISQCe02sKIJv29GiXKV9NGirLve2Mn8gAk50wS1hrwUHgJRUTiyt++O3r
LVQ12nBn47b/wctdo9HHBAguSj4/FPTi/J2rrLuC/0F8IflCxFmIgwdhgKm9c0HJG9KlJYsLGLku
pNOEC3jbwH3EitA2itG2fxzA2SSEeB6dvOhCHBGy6nwysw4OnttteSGux/Gc/IVfBUzy/oukyiaD
7cSVdgYqHerBIuLuzl92xKxr9Mw75Q+qtKs4TptNx84q6sqOqiwA0gOyZ/YGIpyaY/euf40+l48R
g8mjuuUQ2YB3RUeFm+tNzTwkViesIbc5OIIDVPMtZceddLQpF5761xVPU8Jt6ySxguA5pnc7YH8z
BYGAu6suwsCECyGmYnA4xFTx/1Jb6O8E77A3kmxPNBS35keizwOsO0giPVRxWJptvO7PJfptPGEA
kHrwYhE3S0hqlEqsE+hus+GAW7Rwf7ZBuFw8PSbyQS7KEPVtMHWoKQLJzrEdqjwgZkDhGcFcnHhi
WWcwlTZpfqS68oOPDYbiQuutnPFbAsySzbZFgTshd7nJkcl+s864dY0X7uacvicwtF7mcqb5KUH7
64a0v+gZ46LGjdZanoAsciZy2QLD2HuPzawwPgqfw7hMEt4Z46XT+cMsOmp/j6zVfM01iYVaHVia
sx//q5//tBGiFmWJYlIxMIEX1IrhLMyAkedCRggi7P84L0ec5uYS1nb7Xvyr2tc3EQsAnRKGsioR
t8DbOhSX7NadcNunKjjtaFLwRlkQsJCoYjbbPrLfnBXHSsVn7qe8w4njTl+gXptTI3GUxMdspv/4
1xabnoG3CtkIO3Lt+GUdlhE8WA43Xt9OgqSifmlaq8I/dBYUH2Nrdnh/na57SHpgq91vmfavEKT4
YfMlDBtRMAY5dcystdeV72t284eLZXpwhI2ZkKqxOIUgFBk8BmHydrSrg8m+3sOf0zs7mEZwtzcU
PCQIiFSow0DTLeXDSCtHOfkuF2B/RgnNmLbIMDIWrT6n0McJqwA62GMCAoFDyya3fP8rX6eEazs5
gWPQCzEuL7sBj6/KgdzCKviwz6TgR1DWPlr5U6IOXKlgJbRudoxSIwD2JqsAScI587Fnui2OJI0w
P9Cjr8ix7lUChBDMr8IybkGROn1GrNtk9YMEvOreEYUvtb49dMH1yK6DTxg3htErK8kU1przjyzJ
6wm0pfO1swUPUPVWHclxXhnZiiEJDXiFldccY0l5Ci7fpE5FQiq3kd8e2qD67N+eW8zBQBM531ir
EsIiUBTskIUXCOLX7wAxBGRwWv3oZuGWxYCEocDSX/XGmiw31NXwfZrzRkEZaEpmGxKjyeTs1qxy
yQ3fFhZ/coRunArHAwU6Wn63C5yeR1vpKz0FeHAtsXIbwTfGpvOpuHs1kYdytTCFjl0N823DIkDV
fSRXiDpwyUaOB8BTKUme2Dx/YlisIzXRE6+bJ7jSGz9HOmHuZ5uOmfkHz3GCa4L/Dhy7MOBRxPQD
W3wTIoPdhcSJ/ORRO98Odzc3Sbxi1vfaMD87rVwtQN5BrRWMvg5SmHMsI3FDwBkjeLrYGyUBAzb2
7OAvCU8uXMJI3xASOOg1ocr6V5k3JbVCK8KRxita/6VdkvlId4SKQ9qJy/XjutZ/yni/VXWpUIuQ
TCalHGkbt9MPlPD7nBS29m/anNkklR0ZOCr8zxhx1+WRWVRz2n55jJquewInzWfPLUGdQeYgNsVP
uNg0+/HDLvCdGsKM4Ry74iGPApuhD5r3WjUdbH88x2pdD66R3vTykNpL6nZzr+QDP0Vd6fL68VL2
C3ZgtY0bkrH7LEzY9fFXCNwL1969YZlloFnKGMwbRotzAQrx9YzlEZsCIga8xSAF+daBGKj4e8Gl
LkXJtpuP2ye4s6T6NHB2AqOEwSs/N1ZhHzp6EG+Oixpse5XiLgSJpSzDZwfLotCQMldTkcTYQBQg
HgdpWRlFkePXx5eyx0rTm0OnDqfHuiRkuUQBCoVKDlPvYQzPqWjb6TQJMotFytKQJPHIdRZd/4Tk
obiKbv/JodvecRIV/LX0MfPSE+64jJucS5aui/Xy74VNHxLN7wnoV1hIPNKUY+0KViEXzetApnBF
fusi+DcvsXE71D0XZYXnUiMJN7F8+bw2mGA2LUgLmBNSrQbXzRnnhVP2zkqDsuJUh883tAz41BRk
75EKjXIRxSKuFaW3iESFHLohZvL7s8AwPaKDQIbVzn2XjAb+Fwp2aZ8/YMaPUAZGk3kKTFdNCzzq
Uedr7HR0UEndCRfebk0A08nsikyrBL4ys9uVPt/BJiQyu+bBYWU9f7+FfQZqme806fnB6Jv9fIMF
w5OC4lPBeNTw1MC9IDUGRhgg17Owm0XMCZ2qNNkqMwah6SDYhEIrYBEmN+HOg/QC9SZXks3iwDFu
Hvudq65BwbNgxz05M1jSeRJ5dCYto41bzBERYfvVjwXV8cXf1zmX42IgImVbg6YpRMZj2+PblcBF
Cpo2jcXTvFnhkagJZzzYKWdY2iYY8pFcPgCzDN7++ihUrUmRXQbEiZkVaxdli0kfJV0G8hEH/kRx
8M+A5DYrMcGlUElXQ/HYHZ1yo6TukiTJjZPYgtS4tGYGhIJdh144jQPjFBotnLfrkGPmZWsgnNmA
IPBc+lL1gQH8XnQOe0mhzCJOALBCBN+Iksc8goaRqr3iN1+PR4sM3zi1z+E36fbo2QANrlV7nMtX
dgP3cEIMvBi/T9tWNfqeq8uBmBO7F+GCd3iRF2aSXbFVFNKyk2IB5JbMMkOACuMpXjatk0tenuhb
PNtg5gZPldODf5hrsgSo6WtvNMAIC1JuBegCP+/mWj55YxtdmcBrz71W/EIuAlqlVJ5NknUt/x+b
x4ww6qPHbVE+P3tIaG9zCSFiJlA0guz+GqSlmZU2cLbPIZ2sH6praiPUtbLDBc6b3tlbEb/089vq
qlNI2RsqhFrBUhxRw53vqjGWxaPAhwTRGLjm8Bjc/dz5zbhy4ZEBlZpypVIuqiJe5xuBk96u0R9a
cPUs0xh5Afe55E1JV5ZoNZqjq4KkvTdeKWNyItRRWeAONpwbhzen8vqbmiUiAf0wE45Zwv2sTf6t
YvUnbL405GjSVVOXE86PbnB2bHGUHs/vti7VcfLDsx3sL3TFD9Ngpyi/deHZvQniqpTxkuGr6rw2
DLYqRoOCRXkWetsOaOJyEOkBmxBQ0GkT3a2A2q2TL0cWkedsFiNXNsp8bt7QmFScoP+CN7vp/EDD
QFTFQOBF4ym71uCIfnHloB3b2ArXU3AB1CEc3LFxYDgUP3KQ+HYn4ycN1yWNdK6Mm9eh3Se/dJGP
M9ZohO4w0IiIOC+IpdmZOB2+sjyNwG+q+8Cwas5GxmcI/6m+8Ys5/3K6sP/+7DRbheb6votaSnjo
unZF4tYW5cTb3m/pEB0WjYOxp7sW13zmLcUKP6XGhVI2t32hEktcemY5Vusvt3PVaXTQuWV0KX7G
X6iOCW3/V5WTiwpgMEZ6nJnjcqk8t8U+khYsJKapcAFLYKFLGmrDZ3dks/UIFEbUeA5Ny49vJRbA
HxoY6JLYbV3I9b791YeyLkSeoibQVsnQy+V6M48M4Sv7/C8yDfyOuFn2pFVlQw5KaGQX+5RFB1i1
9EkX/BJjupVE1VbT2MS33nlK/qDXFB1rMWu0UqMFUpqT3+6H1jNFYguNXCgyfpIx6KNSPuErWTtb
0sPbLbs3jHiaJOzRwmnlmpe24oUSOPHa56wK2BSnKCXZw/L6Mlk6b22CXA0wNhDlTZZpiPfGJ3+c
KgEtHWXHdla3KYYjO8dnolLowb8NAuwgt5keh/gxuAoEnLKelbR+xZmUyRm4mjiiEIfMtWC6tOvG
47+23W85tivtIlMbPP09rlitLRVw+1pVchiAw8oefatiBoEAVBFdka5TB801odqkwEb/FhuuokyY
kzdcIuMn7RZj0jfeu2ocf1ycIJDsqdgI1+cYP5MIicsHYnsgFw6wJ9nTu50EeM+OVWptmalTfged
QLzDzMo77slxUWMFmjbpxWNbRQjErHAVGWDjBQRyqWgGbJwGO1ooyOLZNQ9xxE7V/n0s9kRIL0Yi
GY77W9vVPVOjSL7Juj8TQ09zQjf3WHw6RQ3WuZShKon1xMk10mITXKwZr3+bcFmZ9ApomHYPdr95
PvXPf+fCFJmuswsjzoyutxxPZF/QpYjZ6/+zsok24r351w4rnZOm9yAByxvVzGtUGw9xBKuBeF4U
ygHjZ2ZQhFzOTNW5XNEIDb5K8jfcVEOFxHcMoy34mhOH8LlQdMO50O9ln4vIyUQCE9LltTNajQiG
Q2s9YaTtjWm+RadaLy31yTqkTm7cNVLpZWqge7vu9xsMrYgPaiejg/+YJQrJWoKxclOFbh0dtiEP
68zZQNaI4N7wDazhgapBcbzlzLyNcPCOXn4EkLMkHPg812N6UG8TFbO90+BUWlwFLijTO2AULGR+
VB8+GHcXNhiqLahyetrugh20fn6k2BRWmW6kZ8/tiaG4DgFHHKWvsXLvlPgmsdb6XAszjfSq1iYS
hwaTYPRdTm7E5q/nYs7KMbjbbR0qEWzot8fYxLvY4+L+ow0X+UwclLfg5oFHcUPAph3ypYh++IGZ
U61zqWGP8noHBFlyCEoB428wg6oeXaovFlSIJYmAyWFgr6/9yJC9bmoxBdmJMIu1CB42ZJmmOrsU
ECxMs51zHdDQAxuiFvD/Fvxw7ncsLs7M3r+N72Ao/4vpVkuBraWzHWsZw4VaoeBa64KlJwtQBeOi
UMbUAiieGrvQXFD9T98pVMFLatifAWRoDLqsEasbr6hQPaxnuJD5dsgXntj5ay5I9K5mkfuLgJQv
9YblXU993fset9vtCx+JzAqKLxmJisshLn4+E4m4Vv43iEWyxqDGJhvLYl8AcDSiokj7u6c3gXaQ
RVs0Fi7TJrklcXLe412i4WJRnYqSDSOYj+I/5bm40VoxKOPIfOEbPfDQJpgML7KjwaX+S6OWLpjq
Zm7/69sIhnOwoiSzpp3bKO99FpDwSIxi5tbT1stRG/k5x53+9pEJc2VS3WjWjekZJIDzC9qBA8el
yRuIF6VhmGS2to1WSsYYqhOJ/zFzGVvrOp1KdoAxLna/ClzL6usu4xvSFe8nKBJuAzOzaQGwUGAy
Ya1iFOOq8IT2rIFWGeYnhdJWIyYkUzKZv/Ny2RJ/8FcNJycyX3AY/HYbQQVnJgrWJiM3iMHK1HcM
JY3nlh656B+ix13M/U/G9qNI2+gYjrFeVMmbMZMK/QubkebuIa6d56vB3j9C+vIi93WdLuOkL7LO
n+xDqWWn5XSJ1YTms2DFMWOL1a6IhcWEwwLcp23mo8vOQ1HeRH6cJ8UyhNKle3goK5M3+snUE6GC
YBk2mZrE/5El/JCuvgWlhV5ow4LOuf4FnIYU+7s1RpwCm7taPEknn99XyUQ6Hhdz6o0PA0I0B9qM
oxJpXlSgE3NDtQnTZZef3IF8idR9IhPSucdXaiPKS6f9EHxBafnTIKXEmsbCfHbsucDq6VYXnmFM
NEGOiRUvX7bsue4hjZKFcIV5I5VWBV8TmfN6MykwInaglB/RU5+ch7jLFrZHyfKMf4X13MxK3iiK
xslOagvSNZ4f886brHHHW4B80cq9cqu/BBYMCcWAQ4gfl2ge/xvD+PNyO83gr1+pJ4MN25tZUCsE
n9VXQ2N5xvO2/OfY8KNSF4mc3DpSj2SQ3dT9scLqJx5Ea50Jg6K8dCH+LVHeQqE+b2o1fhfmvg9o
6AAl8FsY0NPtwMwVI3Ncl2ojdcaio6qs2TgH/LOoZ+RU+Jpdnc9cSAxATVUjd4vi6UH1K8h1qhnO
zzelM96o9+Y65QDLnlThPsMdjsOwW+ZNkMdGkGOPQMRaN7D5jONzmgriQMdcVJOuN/ARq5rQ6z+s
O96sLZySP8/gpZRc6p4ijZyn2Y0in6bTjU2LzK7u2beOZJWN72SoV2SnJ4JpCtav7tBtBNtX2qrA
KJwSPviKyPg/1lkBMiLTLfAXtC0qANyn2CN+4PgRHYoxFROFyCbjGsZnh1aomLrn6JZGuwnI5tTf
+0+LnXyhesFosU9chOibbm4a5lt+8b4qPSdh8s3htjTKGGSwUIMGeothiEfe10BHHEdVLZbQhnZX
9wwYyqKG6fMlq1FMCb8aLKz1ttZmho5BxKP9PZH5trLFkAjPBE0nwiZoNrRedbuwVTkmH2b3Iuxl
DMx9P8VW7Il8tSa9MkMZVfOhkvtd0f8xCWAXzgQ41tRXnd4SK18mBF/0f47Tvd+I21ZJNfS4hIav
0gOWhLx9PTksLVd92FBs7BkvexgqtBHJZTLrfBDyuAtXj6ULA3gy44EVuj7e42I646+XpXNZPqtJ
uCq1LicSxzGgihawY56D16iEFV4ypjX5Q1BvWA8D5aD5G9Nr26pPVVb671NBUIdyG19F9/Jq/m44
7HuEaTKvxTV7Dhq4Ds//yGN1IOJ86VNSB23gaONe/pySqOStktTkG/JLvwi1i5Z+coIiRHzNHe2A
iYZW+mUkF4KP5nLKaa7IfCXuxSsAiwbCHeRwWHGcuXs2dhKnNQH6Fvbfxg1d+FuB2bUKhGeLgGSi
K7Pz6IKNAonCX/XTVCu13FQ+x7YiyQc8jrZU15YCtQhSJMHW1Tov9I80up7/047puWcb7/dk/oFf
0NuYF9K9C27VG2MW5MjqSuiaY8SjSTdcPtNKFw/zWSu+qfU1SM9F5KtdJujWuZaBlkLmbtTC406S
ikQaSl1h9zBQGkS6tmt4JoPnLB5PUV1MbaAGaXMrZXsNWBpy0Tih2VfBeSKh8g2cqyCFUw0d9O5i
4OfZ3HMtkWl62H9nMprTpmx8YQbKsimGGqnA08PEHKBbzY52NuZu7IxmaETyF6BB3eCFWrqanbEu
eoVcLPb76PwbMqMyygW6GFtYNNqp0wosvUUnj2W5V6lq8XKTkVh1rcKEroXBV/8G23oR1ocdLf0A
bh+NdrkI1fe8BwvsGzlXLpbJLc2zSieo//jqnDG+mFgKtEzptXSlXOnaIfZiDfzebbNY+YLMit6e
RmmsAPxF2fhg7mw8fFUiHiDzWUWWUJfERrbwLnW5NMtJVB1AWTyzaa24cs1zeK4vV7/8I0dyqiyb
mLpV0Jh5D0ynqHutCP8HuQnVDIjDhI2pWmXOEqiemIbhM9zPqMYQSCLKP78ucY3+3EhylG+SaJmI
h2/aiLvNQ1wIFOnR2zua61pbpvOpuZY7JJaqeob3CKNG1ju9JW1IOU4JLdHMqCJwvE+l7hcISzLe
5xvIq1BumePniWZnRbd3NSqBvkWSF5A21ZlcN/EtY1rjdVezfSfXOK8SSvNeuOvimagEn30818yi
5FxRUSVZqkmXIvHxcWvRIGzxLqYpzyAfMy2NBLgvbEH0ASNupmfZJzGAavwDJyFMzAvJbyq/sAL9
TqXNbPvgGSfirH7MzGZkKrFWTwgO2B+pvgGekov7ACzFqrWxO4T6OeHjcnx0t+tXUCPpWMZhw1RX
YFVIyq9XNVIsAIoOkirFsee+/a8FHwr9yUywC/QckxutWahmC3bcHX4ncjKxPSU9WkUrh0PbGD8A
Zr7BwRGpcGawZDnCeVz4fzO755HcUCPDkpLbhMklskvZn9vwmY2j4R+54mUUnAdUlR+ccudjvr5Z
+/6IHRproHNtozoHsN33l+Dnn+Pd5IGu2uDlyxWxswC78jOwLxFHFkPd2S9zDcBIbdNadwNzhbYO
YaUfomg2xn0DjcefoioaxpmVdWBVj2bSg4pJTQNPv2fqBEshIp1cr2dnyJTUTqoG+pP9G9w0Q4+Y
dXq5TLQ73R6E6WHIH54BxlJfnmKIyEQwlqKVHXGV45Y0YXRWzY0jVHP29q1HiEopWTyYN4+8IUPQ
8+RGNhatcoy/hEeeMas8vhR/XXqisOx8v6+Dzkp9joGdpVlw9X9DGv64EzEzxD+fkVS/5/JS/N/d
8cr8C+p0S2E4i6zqjE7/1PDbwVWHwhJPboqddOcE2mGoPnnsqtmjBqIPLa87Xe2HrwCXlt/pTRAJ
W5TcMKv+vMJUD246z9DOdwTLiRYVRtiXwJiocCp9J9hoCL2TmWKAc3x24bbgs1CV8mETGdHkOFRr
YvQ0P2D5jAHwKvBfvmyocJOKIIt2saRM8TszVKir5d1UUdBFgkdi1wtxy7Lq5/UFzYS8BK+yIW0F
PuSs3djq2mgKjZrT+eXOHhzQxJ5ZgPgQOzw3dkgiQ9HnO+Dw8EwZgom5bdPwRQU54Pi92rKuFBOb
+CH/hVkgPSqn83pWeJP1lj/4YOIWyXxYVOi3BDHOlLTf07piCO5Yklcoh9FoWlwg3dgBPcARGVFx
51dDa0pbj8AdD72YcucY1jON32q5S17NX7q1WU0g/gCFFEV+OLbZIk+X4bZbg9cbBD2IXsr6j6hp
vGCe14EIkoVI93f3RKTRnEDcXhgwSr7XvwyMssG+Yv65nid/NNfcOaZ7FUE2Dup3U4TcCQ3bT7OE
WpmzK84td6Yb74/Iw7JGUlnES8L5fWQtJtybTVMrYNx4nLodzVdCatUNYQqiV4qIgOUdhjt/tDRX
/QJJv77wBTG+v2y/XKTHCv5gVdw68YOxq0q7IxKsNFPKjmCG3YA5WCP/zCUgVt4MUI6HOUluKKl+
CjGYMuo3bttQJLB1yauvAYfXvyd21Unj8QSWTzqFmKMYj/z8pZeLO0kMstmw6ug823cCQNBVpHxV
KvsBcaAKkMaGmIMM2Nv8fpt07BkNaBAmWDtfGcWh6fV6n2/tCZRU2wWogSUDnPAwXS80+DKE1xxd
exbB8AIQNI5lAIJd5knjuS2EVwrhax+zCHM/dDoS97bVg1ZqShnz0gnXFyAvJsItaHwKxxjgIwrk
KefpR769CgyVNhjbpfGq8v6RqDhsD4xU2856LqvHPddLNQ5nZNJ97oOKKoMbQlBDuyaq1SKcKUI9
xmjJZlKFVD1FNOcWhJd/DQ6ZaUo7VlgSfl15izR1JTrEEltQJji9D55B5e3KFOvPpPGIBCuGUmKy
TKraJn6RN30fw7ojbhZZOGb7COCMz/Q6bd+JFLINBeJL3XxUX8HNCr0NjHagkG3H6QddlZ/NjLyD
Fx5oAwv835qeym/v2zn8MWSneiWvVs6rVKdb2ZdhjeLEhELRYe/o28X+ueN5U7HRYfvUeLnA+8vW
AFCO+pF9RNJi4GDedvSwNgHjFpbtfvNo60ZNKGgsUKcI7sFyYj8CvmLCKxSAFM7u6FTqO+ZM8L85
ybPqAKMAnLqXN9WMaPnC9v5hwviFa4neZKxKCVYXRVKNo7ORy85wFDou5HybxBTcmyJDa41XC6h7
fspvJcQxIxT+OEPo52TbabjMEKMD7dDlPXlAp4nzfV3JmkbEE7d6oeUjCtiv3FMRs6BGxbeHAte5
wcMDjUqcr0TU9GhiOi+IdH8a+0UssrEtfBlNO5BCh0xWEobPz7x7Lvb2FgEUalHZQoBmg2RmyevI
/sYi9y/uhl9LWxm2j2Q1yGNvphAYrb/WLbijGOQZWqJUMdEmZQSEsrpI4VQ4LdPEnlcHf/QYXJzI
wfo5Qj+aClbUSfRe+udAkz76X1RhFQwwfh17exknbBOydwNH0eDsVpg8OgqnFL5WPd4H+e1yA85H
o+t1d5TfqoMx0tlBbS6KkQ8/aBjqFtx5huiHw2U4/B/YFVEfg5uxnBrm1Bcz/Oq/Lnbit6FiD1QN
IE0iG8j/1wcpbVWvcJ7nYq78VPi2nk/8z+wCBpUENsXUGdr47qpfKXxe9FRDU2vHXMfUv+vprjky
6XguMjgLNDkbXqM2L6fC3xvANTrQkdzdok1I93uyDpJX0uw8mHs/rRADW1iALv+Lq7K8O2tblsUT
us2pnmbKIuBwA6cU8HD33wTDWJSw10fJA58r8ZMQ6y20TZP/5r+Jj1pThJF+B/1CQ5am9c1+B+Pc
HMWv3Hkfvk0SqeOzBnDUMZslZj8gR4QNprcqgOGYDLh7eF9phS5pK4mvyKeb8KAHPz5O/ZA5y8AD
LxLpZwa7cS1bK1hkeS170cD4XilbQwbPnipt9KxRKsIuE5mzvJ33sGox+IOEgpV20e4LQqiwoI34
V14sNhKrAwAcQyowc4w6l+SRSFu5+zNjvazUM7t1fdzxI2uImLvXi6z9FXIxnhuzitl4C/UGA5yB
oqrr6d2dXlEw1wMiCLL4x4kntnYIar8sYiRqswNWTFbwBYvaf6Z2CFKWtkzJCTphrsSQ2iPBSyX8
HgVLrZFxD6l19WhkVIWQCVo+yCSYC3mp5CuWlyXswpK1GvI5cNfee7rIctGs86RJude7ljrUhiHf
QCNSH/WNVuquk3RDs8CWUpv+9Lqs/9mRrlXHaeRksXDD9aReq74+SOSWlgnfM4PYU3qpBCHnSCAp
zslK/5CUOs7T4ETrHpG4pXjtFxI1pnJ0tEFDHpPwHALaOsFelS+9xEfoLuU+/wskhcA2KCGaF0Hf
Iw3OMHTLGIPqpaIhrbQ5/ZNeG+ICnui1bpkxdQbWVwK3T89CEi3CUUCWdPw6EDVwsMvd6J9XJPnG
cpSmxhXSA1txLPAXMrL0ijR03jD4qIH6XNVNbSRg6FkK/VhY5ikjp2VxPqx7M0LqVASY+q1443S3
GjOWe5Th7Kxtpy1d06cmCYCl+ytoxiCzK6LVMoYYpqSiEzubdAtCtnjfgL4fL7KPx2qsxaXOWawk
jotJLxxJnukIajvxKgchISAlQXhziezW++Lnvy9bJLk/dprb9YCpZaEAPnKtn6+JrwOfACZHbFVb
O6FNqsDyaK+d8hBOwvViQo1VF0FrfKLxLt2M9Fn0rkgSp89upCGz3QE1yATW+13QhrFjfnNQYjVW
lR5TYu82VrHdeX1BU8FEN89ydoOSjcsnAgDe/BEncoCPEUpHzRfX9O8sbYjqY6qc7GEzdPnD6xAf
PZxXrEbIjjM8I59ydYK8bNPP0F2S5Z4YwsxUWMJIndXz8ECTQS3URkSaHbjFnoprsdm5fE2pYxTh
rNJ4kc2aCoDJwr3bTUZJtYQ5eKXEYfo/54NbYJZgS4T5GzOPx6HiQi0y8COWLhJtC4J6hAL+Bbxc
s7loYVi1Qhbej0J/oI3awkw87Jie2JbOqs2n4hkq+eU+GjG/6+lD7xfuRHwMH+mMtqC6dmdynHW9
XHU7CtxTwFtSSProM99o1PaiIXOUvX+jVmXkjHjWJJfBk75YUbF+r9PPmmeIdMQhvYCx/VQqEswd
Yuit/BupzIaa537cZ+Q3k64jvUtMddUX5GctlgSsC8sWkudYZhtSryigH3EQcWWEgb5kdVaqHIYD
KOQWbbykpoErJxwC/DH86v4MA8mz7rZVSV7pAdxgOXhSCmuaurCyvvJo8azuoNNuJ/bFGWE/Mn1J
hHkzeiRJ4hiXQ/ZlyYxvoYplQpL/5U9EyYFxjYLHYCNM1YUKD1wznqIv9Z5TvGr+qa04wQKPJ0gM
cE3+387Es0Fg8HRcbqFhDT8dtEAMpJN+mXR6xKqf3uSwQp+ko3Mch6kyxNvbIKzx/5U1S6CQ38Ob
YZEG/cy1eGm+rTrxSEbPRMEX0MAyYxZGM7d/J8q7SV9uXsms0952orqujqHxm463ZDp8fOkNqIhH
+xygMlGyz57fWKn0QZNdaSoJNU4sIQ8Z5Ffx7Qw/U9v3e9jL73Cr2YUNuMVQAL5JlD+h+wOYTvOo
fe5xjWU5yex4OuBzRFhIWaDO6WLyK3EcZZ1X9wulB0IHbqq+1pyAlLb0rg7ma8cq6QL/6SX3s4Dy
Xhi5w0RGzvRMByjz3uMWOd0unYST0WAB7PZTH7zxgJWOPEj4l9xJHqDBU3Iwx8wK18SZfVjbZ39L
aIhADYsbqaMNmNkeS9QKTFNiXeD1L3EFXCdQYeXlUqdrj3Nz6YFAi1Ern1MoDn57rITg0puTFxtL
+nWCrkt9AjAOpiQwH/UylEa0W40vlA2yoiEkhYj9gMQYjaze5GiCwPQL+uD9RSj4hRVnIbgL0W6z
wL7HL90z6KITv7FsHRq+NpPXEIJFYeD/d8XRfsCGf65f8ei1TXi9+FAwfGHseYV5qpQhANoUNm3b
J4x/nhganumyMLAJmt9lc5GyANf07QsUrWvX5Kgvhkw3SwwDe1V/QNHjB0VpbzjwbELTMgZDVwwv
SyBCniPyclE8DiajKp190XS+tXjcScYyy4WgUXybs8VskxeUFXN/ufEseN1n0DtPsU4R8FEGrENh
+g1k4pfaQD51IzfQNMhLJXss/MTY1Mq3VGTLCfXz0G71ow1fsehrlxvWp/MISIC+Wf8ctq6VX+TP
lpm+VqsFKF0qCnkf437ULFIoldsOzpWcmSBOnZ9bfyRNGl7nxCw/2gFeuNwejmvqjmoexM5KwvvN
3pjlS8LbddCRYjZxxB8VktqJ5wsyeQ2cS2JxEkYQ4qkjDUvAimWZ8Dh3NTywaGDtEbN9IcRtEy/1
PtG/JYNbt8EAynZQOFduAtxLhJv78/Yo2Ck1RGG4FZKLljInpuGKbTJP8RoXQMP9mfkQW82rwyU2
pTrHxz2XKD0K4Kvl/LhJPF3z45OjmBV5kSq8kdusyL69lrXesOalExFkJEtLs0JAEOAi/lKhwFkU
SWlwuSMmbVXJshvjREelgwbRRc9RIXSoohZ+VYAkrbyIJT+buIim63itLU1tz5t288wtV5xq/6/p
UKNz5EkNI2LBuu8E0i7VGKJ6/hGvVUgsljRIiHr/mmhafOsqFsYWHjMaq3FKqqsvi/y3n2g49oMu
p3aro/O/UKEg0Npusrz7Gb90hgUJ3WMbBcSjvhh5xDTycDWkIP/+t/AP3Ux76q1Gmp4zEbPTjoA0
QWNJydy231zDGJhYhBLtRBVzPxl1K4f3GnLztfxKYP8dd9bP1lcauW4UZV6+dohwA+CD/LoclWkv
ZrUj+Fw53RCzPPFoyutWrUZ39y08aM1wEWgEIcQGK2i/CaFeyHXcrnCKmFmfqp9QHZ6E3OFav3Vw
O6fMIiM8RMY7Yvx8W075s+T4ZHTPFtXgdra7B0v1jGJmlEsiTNFljXcD4UtpQM0yz5PjoTx6Eykr
ZlkoNgRIY4e6Ye/bKrEM7quFHUoBaNg47ab4zHf/dTx/sPgTT+XfhfduohAkv4atM6S8SY8hvm4J
k/KEpS4woRR6km+qvHmU+NK+4PAtXFXolEdaxxjF0rVmKyOoJjKVMXldFAywDyK9ytETeSWvML0v
Sut2/9TmOY2NzSrKDcNvSvB21tsTCrEGa/lk35aDUz/BLbNeyhlydnq2S/K8Brt+KeYGw1RyjPRR
GlRvlpdpcE6PHfeEak0Wb/kBIkCtU5qs+biq6jybWe1fWycB2tMS8Gxpbcul3zesBoaeqCi5UfCp
zGK2006h2qxbIIr+IIc87+EpMoVi8YV/zxl0q+aX4hPQAsGUP1nwOKnQt1LpW4QuHlmYAbT8OTkM
3/5hzBsGEsaQn7onXDDE9P6rKdspF3ileWrfFhw0DhxdrULUVZKGUyCOTXAqKm9d/Sp5+Aen98X7
th0bpZdfyCpCYajRvcIoEv2DKla7/Zugj1nEOiN+Vee3KriEolZkaV2RAFF0zB6GEcHew1DaqT8c
c9snfxyPFbeWFQW6cUiHVkEshQeM7969ztPKOJ8yiZ+g/ojLVIsrmHAhhzavQoy6BIOKEF5KS0Fu
Ayq9jm5ySfZRECcAGfUjoH5lFWyT0aQfI74qs56YjGXtW9h4LbOMUHk2WSEs7NiccViiA89EfKFJ
wOUKKJ6+6+xCQJigxaq5OpRMYymkg8ABfDI7M2v+aOPOIAhTSGVpVg7EKkfI98M4/CQyxh0lK2it
YclzeoA7Dsax7bVenwfyYLEwyM3Gun+I/Dn54vuZ4rdAgI48YxHKEjE1yocvCU1R6pJ8MtkunNLt
qkBIXsyxdgq3kcq5JPN88p8IMG+0MQIaTZ4ObOg5+0IMoxs0shoA/dvsfdHvHrbgvtMzm90l64h6
vGuTuiYrY/lP6czTczi3+M40o/MAmV/DHOvAp3F94tDPaXfMBoAID4M/0yg9KPGw7xYfxtEkAlHm
sdLaC3dLcuWFGgfLMyf/X3r5lCSx01DE2b0uA8txQIc5YYttGIi8Z8cS4yy7n5Bvk9hlCIPfH42c
P9ZwM5mo5StxYN9E4in75PQR6xCcJgZ1Ay39mvrV18T0gHGN8mSyEUW+9L0wdULf4MjJ3M+nSU14
hqWRbuVEar0TiWV4k2/U2N6ua17latrHXwd6TnwW/ubufVLTKXHUeJq93Dz9uuDPE9PgDyL1JZ/P
bhS8HyFxTkm3cRhSjDI7XN++CczPZtG/6oxlIhdd+XFO0a0kshCgO4zM6dnkStgAmLZMrkMOW8H3
p44hAIQ9c5zzBb2OvTe4IDa01EISikNt7wN7FnWXW12aOnMTXozq5RA1qT9/ZjGQxAgyioYfx/PO
9ZeftLszf+GeFngUpcwPHsF6Ooe8ETf5mr9JK2oxlM/Wqy3MRZiGRSqus0sMhqHUXX6uc4tpnmVL
FvXe6otI4kVnnW5mBwYpKKcMfvCZ5qLvNMqoJovmOSZ4UPaSTeiBHiN7VBN7avhcTNi1R65/Lono
kSdkRUgY0ws29v4uDTU0W7cG4HUzj7bIFeb3uokqicG/M4gChUl385X26YnDhwufR4WyLJKCPxcK
7sgLCW50ZYnwiALCy6DUegYVJsBbTNenEGsAxrr7VJ2KJTFSr5nKsf72vGim4FFqJ1at4Yn2C/6c
9ab1kT1anx6LAnetPAhzMXKUQoNYoRE9oBMB6V8IGWKEIj4gW9tWfeOhQLEh7ZovghDz+iylPMqO
uRve4DbpMGop1TPEgBV9nejK5E40DXEJAHttYxTHGMZCUZCsuRs0qNFiiY8PomZ1AJL9qNLqvLez
GZOF4OMNIQ8fA2c+zZDV8/4LaC0CHApuA9lRLDVGyUQNWVb3B+LpnzgKE+Tlol/ScYPwDtprvKwg
PJKaMtoEXq7Wb2HAKG45pIHNlDHvDcLsMGOz1TIk33/kqmuvhP/U0RsesXo5sg7Q9o3tQ3ZLvwwL
kWZJztnzDatUg1LQwsdBPsxstj7twpVfNqx0ZbvWmpt2qfCwoD02Auo/YYBqPkyZ+6Y7H34a0OAf
U9eBQnJr5S15QZ2vsLKbdqFQujn7lIXGe1NMi52N+I9nvXQ1EmiASmzLMdAEX6J0rdamW1MtCwXL
9GteOPaA7Jx1HY98Ud+/CcDQdIkYzIfX7uqPZxreEEOSMlbZO8VMpdk7hVJxHb/zZbrDKXdc6WOM
+wn7Yu5Tam2AMmgI5R1xLxOSMuP87o3HSudv0sHmtP4xXR79rw6HhXHNIZp4FBCFDMbuHglPVtBw
KiYkdLjbommyW8HWf83srZe4kNTmhvkfCgCLltxYyHe4M+UBVdVvBxuPC1BjUaWXKSrihQXldC8C
8GiVusvL1nH5eCQqkwmvSnDy15BJmGMTivcSQsqya3q7Wfdd5FiJ3rWRZU3I2gGVs2dcJd6fvzIu
pn1pe7XwO+duuefJgQGTbf+t7S9TZL0umygzahDPUZp5Ck5vHnJXynOKkLX7KjtROlkLrxClJ9/o
/HS2tEIlaC1VtY9bLUxsfHz87HmzlE8upBeYwOjX1NfZsLtjO/HP0sK3COBizsbbbJXLe2o6ynvx
mxDO81TafKVmLdo7kJgG2CIQuf3B/DT3W6pWSypotZTtHi4kKzqZ/cZ3bf27I7SgvivpDEE4AsP4
ZKTJvB3KUdeUenuB5tPCcKgfIPz/vO0NEFFSN06u2OOCWPCH0+vGw+Gf832f2eXGYfyjR81tzoI8
XZIpiNEkqvmPMfcnA7wQBzKewc5hD8Hg8esTSZpT0pfhCxvtSMmnKdyfwzyjRxIE9jeFMajDflfu
44OCUXvaz59gAkdEM6bj8izO4Zt1dTuKvs6Asqz9wLioqcFEOzJiRPwWGrqRkA6ngBCU3vgdBECL
1/YLiXvhenUnGkENOzCdXdwXcq9kszTHII60nhJ0vxgLNtq1EfdWBq+PoRZXLxNJ+Sdv6Iu5fVu+
vGRL45od3wOXAfbag01r2MeUhhV3BFQs07OGOId3CI5VZcUuOXrD2HRllp/R/1iu+D8E/mWRZL5f
NJbD3ZlkBLbHbwVY+HhKh4+QcOQkIFwuBlaDS0uxgDZCAsiEYE5RjGgF9tsLxrU8rjV27jYCqxKY
BxuftVHN69swrcKR3t89mmJ3B24H/vko1b/zsEQYu9b0oi30XtgTXrlTuJz3drkYDSWkVKhk+6dA
hxiD2484LBPAME4JY/fANeV7s44DPN7XUDxut8g55puj+JgiLErfrnld9Ec/zGVsEgIY0BzSH7II
eBASa8ywoSvjdN8YUaTiRdstIdshwUxdD/kVB3ha4WHNGVulXD/YYhTqd0dWeuLLfnof2M64chRi
qXUKSl2owDU6jkCXRnHZFrsd9Xb6U3nx7Krt/aDi0gwBOIkA9SreqCQ0CF/abKYV6JUw+tA/GGee
4r4Wx7UXFO0913C7oRx0Hf5WoAcaJc4/cRgIH3aA20Ys1yfjYz7LLKGk1C94lPuAxM+yAD2yXss5
AHSbQEt3+AknLSL8AFysslwFwpk/UczBxwNCq1LZH6bDny56H3748KrV5P6TF20IKVgLHIN87HK9
LqLzv4s+GupXRdt86EQ0/wA2Dr/zonyziOgbI9HAm/Xw1pO77HSYUPB+329eY2OJhT2n11dhNO9+
3FjWchp0SUsfm1c+bv6beymMb1ibbgqnMicVD7ZfR+Doe79nUlUaOSFOfxRdmeh+7ftZz4HQy8do
ef6z22jObMgsKoptdQx4Hoct0glsWxlKFc88SBAaswUqjm49gRCHpaCC7V3dE7lPcAZoq2ta12Ck
gqj2dfNqtGAx40wm0IVCKo5Tcz0E0XutQCC1Z1wuswlSL6oVThwaV+xOgNBGJoTXZkGdsAoMNu74
H3b2jpRNcmOS2uLxnTc3vXWfUbb7lBMmJ1FSmGqddTdinUHaNAhcNIXiEcHYBpye3JeShqacUEBr
aBVW2JVkR6Hb4YjOmI4aeSDdMviHXIM6i+CgHW2dF2aYRnkyvIuwoD6WVhw6HRNFzZXwLE3aBp+k
FJRDFhqnBJ9ZemBkZ3rO5Wk7oUgk+8dDxUV3h7FZx6EzNyCnQkzZshKygbhy1lve/HErG5zlTQXy
gEfn5fpj3doD6xdJ9XP5jDvs1HzOoOVKex7qpa5pOPcGiPwmw1UXPv8kP4Ac59DeqdvWyDOuzX2H
6KfM0WNqPSODtwTQkyiaeSCCoZMsET56iPRKiAZcY31/CSLngIBBC9uPBARc24/oYzkIma5Ca4Sm
yK3N1KPczeUnEHQnv0hBuXPNKQQKAsNX0OE8RvCJKfIN/CIp0ASCJYB7sU37KEBm0fIbt128E7ps
VKWDpwgZ3RJ232BushP9VB+AIHKhzUivcvWJMkq6iAO5mCr36f5wCED9csqHv1TL2D9JruyYGVV1
Esw6mHLdv7ov0YSJAnlwgBtL93twoDethaowPOqWsmXzfykltOngFV6oZba1L1PRloiyeQbgtAm0
RAe0SeJlU4BYaQrO8P441/xBi/ue5PJvUjrDpyVYZ+RVqPs7BZXjjvabhf6mZzkW2l//iHloL1Of
u4JYmCIBB1XeZBd2jGdZUFj01Yb8atFp1UBfcADNmVtN7TV+BSn1WqGAjw5+fmm0hdHlpL862p1o
cndenW01kww68ON+Cbf8XqMv9qblXb66lfjx8OKLXm0rKj4IqsKHqKEE4Z1OI+k/VciiASe5VQSc
2BY8M7FAmwn0rM2xyP+1VUEvDJRMaL1djZRgJbVbXNJ1aQxa3v8Ivcq1mWDRMRUvbhP7rnsJJJ5P
yVFZzjAoyLHBjNeYkmI+X2jAtxVEflkv+OqSVNEK5t2wlLmkI3Lmn5MHtkI/h3VuaJJVyi2+Y4My
5HuzT8IulbcQiFnDELnzgsuF/tRD6HMU3cg8OaJ/C1DQ/ZqF7XAjJlhSxKnYx5bN///o6I/iCgf6
SGNLTmBmNIlzj3u7/BTF7WUgt//L07yRsJKMmXRw//XgD9YvaeZ1kdphUtH/5uuQu9rnS0N7yZMV
FkqYfap519hsT/7tZus3tdf2zQp6JCZ9gnMWoFVFTSc5eRPKlJbqdof1UFoiRWg+iMbOkwD7/eEu
VszYHKGn0K/h7VUUgMyb1kLwbwZC5A/J7GdL8byFg8aBFUnL2Z1RBTG/8Ls7ttwxi2bFFQcg++wK
Ao4OexoSqs8yniOOzG6wsEORR2xXA6qxSeY3RZoidRW8/bS+o7LM3TbJOyEimDJZJfwvmanKpXjo
MJADio3lvM5sC/1HAhXEun4rVewnGd3ORiDk6gnwqAezNPsl6lataFO5hFWCZDwAK4H55tCZdT6t
f1shY0e5KeZyIFlNBRuY5BVGMnwhQgVg8m+I4YJBVgJ+Px9Vyj+M1zsffKYICDmI0PKpOtMzlv3k
3tZpBCNoBP7XOBFml4L4RWQAWQwEMWpwKP5lzgLVbcZz5hQyVzJJB1hycAmjc2Szkl4ZrTJlYBcZ
TwKkm8s2TWzg9eEgDBduMhZ52AB1/AHp3GbpaXOFcYnvK+Ot6TtZ6AOsTDmjD6xrcbRh31TExG/B
26b23ZFKeweH6gGOt73SfgD6w776Umgi67cM64M2so8yss3GKqN3jTQFbjEmmkbrM9Tj+r04maAS
P65XBbC6LjtMtoqa9rBRrAPGmTuz9s6bFOcR1DO8suNaE5E06iJLzerDsvRictvi/JfLRA9neGKo
9pnOvJlv6jIw9rIX3XdwbRDTqqYvWF74mtR/FtRzi87/hOiAH/kd7863/iM4RG/qZ6pl44yVyebX
6xyeW0EzjlErV0zXyl7R44USsfQmRB6uHJzJOUSxgRAsCe4irYGWzVnTmVqkJGQcAaEIiivpAMTH
y/EnhXojR/5TGGH96UR5VSVpv9O3IIbXH46wcodZ9HMI7rLGrAC1k1L7UOsYKmQTaoXcqgJo9aVP
D1FAYLbZFO3hy57MtBt6ISDFpe38Wbch9oSy4YAiQqsGWtZvBDuMTyooRfCto3LQzuRyFav13Z3q
ISxJLM3CN3Cw3nP/JijBUojs3E/BW3v6hLkEXavtDIi3LZQpjbWbCjDRCfuBh4mrjkTIwj7wQG0q
92ll0fP0d7nClt3K+HikPdt3TwvXDn8wO2VG5HGkNBHxJ9kwqS8NSRPyI0/1taZRi9RJ27bKE4pL
CHmvLGpuKnVSdT3Lv+n/YViC8Wv2fGvHsYyednwTzWGBcUI9GlKYkp2xHeVyOBzBSxg5+NnC577B
Xa7YtLNn3+9ewAol6gwS7qd7BGzAKxEZXDZHcHtosPeINLKRAA+Km5S3tT4LCS4YvNjCvkohQykP
3FrC0Gavn8m49LASb7wrqiVx3P6uo1yUGKjkpswnxcXRcRVmTuN3amWt2IGbh75H9NnsHphOkigy
1KxNTi7ALh5O5JPsw++UkZbclnoWFBdWbziFP8JCtV3lmCGwb433qQwjtNmMoCAma3JVe67pzOyN
6ZQkAngJU65VoYxUaZk6btrvuyd6Oewv1JqOTD7T8XVzdsp9V7wpAmivK6JlX8Dze5VG/BNPGnbu
yxghiFDubBCagksHzMFgvt/xElXrZgl/dxslw8I4TAMUqLzpvgegodY4RWdiqI8elFw4NW9JMJmd
1AnHv2iWl9LJTKIQfStq4GJehJ37VmPtnvSFaVppXR4URFbawTAhLNwBkjerC0SwYRjTdOzlV2JE
u0whTDKKtiuypRty9wjlivynV33XoKdxKWSOhlyEn3I6n0kPt/GDhg3n1o5pgnw8VRYVWn6j6W9D
4S4L67WYaVRlQmjkGzeZznYxNkEnyoSD4/C69cVawPqUUcCr8pSgqvNn8XYy1CqRVtRnvzgesexz
Es+eEaHttKcD/gXGPOY9w3zVqge22c3wsXQEa9Nbi1nYq5awx8qnNkJJ0//FPEeEGmCfh2YCpkjw
n2aZHuvZOp4Wl1GN+L9t6D3NejfZO1/E0b1yU7UZrfU+kp/EK9jBpkxSjFPvqRFIJGHB2lV8MAXO
KoyATxBayaXbjQ49f47jeWScLYsA3eCFYfYLSA7lJjF14XJ5QYTMtsJOPtytOOhQcsaeo/OZgEnc
jLX8oA+eS9u8DisSnDqOE1ZmJFMO6Qo4MU7mM3KEoKmILTmHbsyI24fE4PzPS3HR6GEmg54EsbNf
akPtyA6RFK5z+xxnrYllZTg3jGZAxMzi8KdOkfZ2zWOYcyNklm3Qn3Lb7yMRAih3xxCeCulQdjgr
Gi6HKeFRz9I9JptnG1vcNYhFvJxx/LKbFavhulgE9rP6TvZcafW3xWuV5D44WeDAOKb3FvE3iuUR
ubgaOR+6l+BEMCZ7jvjWSvta88UEsEcXE3Lfx5C0vImXfEvYffSXl5j6YaNGPylIOh9Ph9+3//Tv
oq645qHb5fSQhlJa3maSEjo8pCpjpLtN50drmY3TvpKpZJ4B8uiEXsfqXz5yxg3fg9pCv99NaZUp
uxUQECDpSb8IHIlozdOGMR2v7FCXgoKe8TFC9zkp+BQ/p1crdUH6HHEjyN96KWFtn6IPGXhKjUu9
VLrrdFm6ig71t58F1p5tbDRVw/b0YcTl1CyiAH2galuUS4duA2xpETilJaEnriMkt9V39ZpQ6b88
ywhCW66RvVbsuAoBo9yXzRf/QKf/ATw3YqGEQLdx8lXd23XzBxZBCrY5mt6uuM5p+PoplqMbWC3E
jtOugjZ74R0CIyDSKATHTmhO0pjb5C2h9pzglM3bmL9mWzYdDjhQS3MsqHB03JF/sdB9dBEbKuej
rdgU9LNwIooM974jEDBMm+hS6hQJDWZrEHyrurHqK1h51iXhtDm1fE0id5G7PaVv9XT6NChEuv4o
PInJnrsBoaO7VQs70PsLXU/2CQd4R7JWZ8V9bZuRQw4yoZ19YLNUj2FiwI5xA8E+jhX61UEfW4zO
ibcLPre+HYzk7EByDBVOcD9AAOmoXBlTGXvSpmpsgS+5K5bq2rq2ldnCEOoPBo8ol1MbsYQ4DHDH
fHb3BhO8plhjcAZ+tC2+SXaiu2JmvewM2skUiXiB9KZ+aeJ7Z5TTxeVzYlW3kvJy8Kmh5c9Rlejt
se8b6Uu/gF9lzvkH4ZmWoub79BhzyJAFtRMAcTnuIKBRox91Zn1zSY3NCJMCxbVeFU4nhtzqSydS
QbVT0N6SQzGh6GkC+yXGMxanlJcgJ24G5nv5bjViJgL2ZscZyJSfFlyWSuj0ptfuOcGejhgvsHKD
b+HYbA441EFqPQVq66qVezTs7gP1STdg0ynuaUg2tJqAMpi5WexXMzMZvKp+oUarPaMzsVHQz7VO
ZIm6CW9H7oP0SAhNG1X4oIS9CvEUyXTc3Dj23boeAg5o7XmRPfI+2Glc/GMVAZTkx/Gi5M4wi0n8
OOGs2Qb8de3GbrlbB84Usm+hzVXZfW/9wVksDGQIrw8IV/DCHKAi9ar2RetkK5ncRss+pQYmyVv8
UAhyKPdcrapjkYMlPf7OIPs7Lmp6dRH1C4UpnPveZORayevaMV22mvZexOSCoaSJFCEUI9dTMn3G
KFQwxSLA8YcaCzSsSQh2dF9OTLVj5ZODVNChAXxDhZG2k01d8wOKjoTK3mNMFgDVYve4bX5ukpIL
w/JlQiW37fFM+TvM1Uxuf4DqD/gLiZD428RXRKa+77qjHbPg7m28imv/MA/Nyz2t554f3+yWJNKx
Ay/gV4WxLfN/ovwIyVRnxGheXp9nitpmkpUDKFptmSoYCa9xbDPB6WERnlRGvv3EpIOO0XeX8qG4
AzMH5R3Ik/gD8vTMLoYtgdeaZ45pvKuwlBGWB8o1dwqM+5k5sOiziMuuP1oJLK5Xul3o/yLycM6s
qaU04PT0l3WJVsnkCZiyyACk78FUrdJuyEhy6RQBZIQJSdpknEzWmai9g6IF4OyYRkBEMN3FQ0yn
Ke/ks2DqmZ0imzgHnLFHP4cdQ6gdnAT901olGxaTk9y5/s+OAOcgPMk3Q7Yb1GiCeVZVBpqxctGf
PlX7tucOwN+H3zhgePTq36OFY4VJUG1KT24v+Z2tuaaX9D+y8IWZbeE6IxdEtf2KZoeUw+edpibG
YAN9PNu5uasVBM5JvUULXSEjV/IvZMCJqi9Wkw/mf9hb8yLRIXmXQF2nBIirKivuwjsdqm0fK9RU
eG8dH2Z7rn4L809LkEKfTRRq69N3+OdvcaQJg74yPbgrsCfLYbxo0wbdJS8GZhf/PUbNc6Eg7/R3
HZDtyZB9i7Btp0MAg868g5K9/XexZ5ZMpoyWgnVgD5Qrv/32GpjWBtp0aAEIFBST2fOvNdCHh5Vt
yRKU0JEAlpiGfRdB0YdNfZsIcwFaiS5LkilWgeS+d3/99HohQYNQTug6TTjnSSpNJVRj7iTfQSJG
LaA2y8iTNrZWEPV8NYatona9KFratBMHEt7w+2rPVkRDyBVr+WlAY2bSoOCvTBwFmCUr+2tuoxPL
3UYqiJA+n0X2zw3zbh4L1gFj/Lv9KWSf+t+TKt8bnrKoesI5pbRSEYMRkNoGCus1J2a6LA8CzDYr
JqglW+3240enl2a697e3LuSm87H5WiEl92ijmwFIp7EUS4mDySDleWejjHxdj9FemANCwy5XsNqe
PQve+RyDNsFz1u6EHLlKujT+pel2W3QmEimyYNXswRsEOI7AZ7HXenP3PtP+dDRbibq1KLTDujMI
azNHDZiiHP9z+LatEPJxPQB2PcLong+8CYAiwi8WVpu1LFhZObAQTd1vtwzd5iZPfgw2VDgDGRgz
iv2u4tEaAfMG14njT9llOTTwq3QJvSWnTtkmauNDAdYA2KOIIde7FaRROkIzspnmGmrO+g5NXudH
55RfWH+vcUC470x9ffPIniyZTAJzB9eu+eI0NftSa9MEUiEHtCWwk93dYaSLHShQ5+owzAuDvKhg
Ak8AaQEq90daJMVFdLkOPuSRGUkpE489nbtW3JQ1Lcz+ap7wgRYHJ2RPf0gId6Y9FEIkw49hqKbj
eKuJpp9gdX+6SRzSAYNJsTkOGW0GA7CJes2k36sQ8IG1P2jqzR/Jsp8U1j4pIcSTPaMA4uduWFnc
7bVACIf98mvG3bhIORYg22hVDjVQwsxO/EF9HmjLk9ggQqsf+4C61FnzetFZJYze4/o2f8OmdZMD
6aHxbhQofMQwvllOL28n1wXv3LucpfUQeE6BvDC+eQ9i/kNlBLc0k6Fsf5V5HLjco6l9taXDPktx
3AtOuM5HxbmHKwUdmm8oeK6HDhjMUUnldhWkf5qGaWDPfIWxkkg6PBxATv/LNczL7ZGz4HLloNrH
7FSjoxhBz1p8otarYp1fgeH254l3mFRZT+z2ea4anHNtxzQYpIq19z+b7PjqQlInoKK38vCyKkSK
9ZRRI+58CdmVnLnJqUtD1keKBjHNQ47UfshncZgDLdg8ppv/vBVY1Tx+5VgV3fwwqcAEkxusKd7b
qkf4X69h0XsKv5803oAunLjKwWqp6pDstEZwNx6l5lIFp5xuBhgGTfozW06kd1m7nqK6nbEz30+n
1dooSDrXpqzTo0TwVBXCzKjXJCZvxZmxHTZfLJbdTlFSazmRpM5NTsAjRnkbrIgyFM0Ne5/TelEQ
K5WL/e5jeQNYz6+zizhk4Hbzge00P0iSoZ5TL6q5YqqCUhIxHA0VpI6LNw0yDkmcgY5IYR/60kXm
DdaPVjm/BcwL/7tWcfeyHQLeH2tLhXBt7KFekq/DDuivGFooBunYAXK+yPN7BA9HqeE0eTBKexG9
lg3ea1D6cHTe/WGAU9hmBYpK1/z/XbVCpDRAriKKtBHRjel7VqvLRR666Wk/Nw9ngfRDBzjmO4v0
l6Kgek4BpM/KE9P3MW1zy04XJsyGzdZa5Mxi/0mzehEVjZZtdGmGNxPztj6u9rfA+smW9fcGZ1re
H5b3XMuv/S09Je8zqA03nhP4oAbGFYScxtZI/qzAF7SJl3+qET7rKHOWfVY/6nCMLyBNO3ATgWY0
I2BrJzMn1ay64C9jDB5XqUiBNwf8QCirdfFYz0sNAPuWjjIpqRKBaskcS/s9SHEkZa+YBDIsuRqo
5aH7+uEQ9nsbWWZIqMPglBXtHqrOhMiOYF8lsGtHb9PxGxovmwrS1VXUhIsDxVOZtdCVRagtIJ+b
Dumjw2H4P1Sv7sCPnZKfAvnxv2GmaDZY7PQj2SRnUPnIS6/mEVGGHfOkN7Mq40Co9iIEWB75NBzv
k6WFfhsR0BeQ0lgUY6ba0aaz23S/ZUw/TB/FltKn+KDuu0W3OYIfkj8fAMGiL5kp0R1I1DI0BLEM
YUfNHAcvrlQBwINIGiXAljtJGolVfxTw//DJF7C2NSO1Jqrxte+gMTxmY2kFEuEYzz4bQOBmstpt
png7VsLZSXr/r2zNXoCPnUilpxItTQh7DZc2Ao4rkx63RoqiZFtrs7m0w9219m/zAbXmcWQuLKEO
JXdEPc0hBBranPIMo5OYc0aF0l11UouBMrJMuy9/5lmhXexGGzncY+qdWPBkJi2ZqLxEczSGOu+D
5nGYnfkTIjYxGP/4cT+B+VyW07U/ozJi1azWmtgLsWnkFZRTpIjZHgCkyGxbevpA9m7s5LZQ2okR
xft4mMphlhqDj6XJv8EVAcywjVDArzUgGL1+RFJDVzGGD8QGW0nxjAmgFRWj+zvAtY8QcMoVaKE2
ZF2aOWgtcJvGcUnBEI6YACeLMYdGmtD/CIwiX/vTooAFBCh9exVSGEyeV0L9L/r+snjcofO3aelv
zBRG6i9nNo+czESqa2ADJqji3eQ2zdddmYGvAPc3IIuGDa2E42saNOMBNc6VzJTdLJqkf0FGHwmI
3PjdAQFrS2db5ucmgRUNzzIaV/VMoircmXb0/v2rOzlqGZ9/aRc4VtACBTT9kBK1lKPqLSm9Hmp+
77+8HkSDKZdzdFAU5PkZd0h6dkAAlea+ywz+xpBFSv/GjIjrkt9oH/a+JXwZITSYKWcqpF6wUiZh
qa+oRt1WMx3jHiJt99gwP1MQ5rLniGSsZWEx9y4KojBxCpPyN45LDPewOxg/1u2gpiADdVTU+fqj
02t52wTmZbF2CQ3Q79jZraf+N4ZZQCNsfRmw9QmM1rb/a1p7u6dywnK169O1J7tG88/9WuPYMc+z
4BlEHhgXRyLv2mVFUzoonMIf7aQlxsYfV6b3ZgLP9SYK+UXDHnea4Nn4wCgwkT14IxhFJC6jQzgs
ezTbwNIssfidDgnQx2YYU7rC9hjF+bi7KbiTIVYmm1NjvflXiMhvy4FBFccIyNDR2X672dsN+QYc
lxtGcPOyhlCC/B3ZCVq+mpotpACXtRpQ5Og/ssZ7wTz+jV1z6POKqogwyICHXN+I/0J9roWbI+t6
xsuFBnAOKbvNMEsk9FasedyEFMuxU4Q75drWdjYR7UKwzUvPJPKjHQg3m1j80goIT9F+yWM2BLPY
Ia/u++ndfvihnBL7aVg2CE1udKEc0mOaHvzzxAi/PuFsdxROezkQ2KbJxsprezt1/+scOVg6kks4
EfJzTWIRqFG0i48GOBRq014IbD6Jcu4sEZN74XyqEdbzGahwQMHgmMlNP19QCA/Nt0doPxrmbg6g
CX6M7X5NNxILhax/KsrSDkGHXv87ZhsmxcYl4EceqAFkc4tykRwYmiSz2kBdbma77riYA0lUxoFY
n80iReb/ufz4LuD4nNV5TdABbQe0oQY0TY55stp8GFumCEXdjHspw1Ql5xe0hhCwlKNyi27V636s
g/4nuoGEdHXHsjlREu8Io6xlyIDdrD6MImkNDgE0E5o3ur9fmti40yYD+xMqN/LXTROTkrVhSCW8
HEhkfSWGgAbWTO2YrOGYYrRX3ju2wd9hIIB8/qMnVnQUTCfM6NX8cqsK3qQqzbCTirxscDWeVjTf
VqDEiJbxQzH8AldIEJFq+uvzfbyOtINQ3SEN1blK8PBhzQ1+hF247XQDD8f+yHfrJg9Og+FqHlc3
2Ud9muM4o+jlG6XvjhS+RaQONsvAbKsNgGlt/UlYwN5v0hZMOSF3MTTGyLLcHH2lDVgYuuNte2HP
L78xNfCIw6lV1N8Xp5Fa1+FJpiLrnnBsHHhYh1GZ9ELA/4Vd0qcV+WPyQNi3+3HLYFJXRmRfzNri
lXx+HdrKWQRISXAdzZSiUiBdgtE/LtTVwipQGKuxh/PPvgOPXQ3x6dDgaNta5/v+v68OS8wcBh4L
a3WofvlxWcWiBTHT9+aoYkwPTcRLoPfzUSbAvEIeJ6Ou61J6RgJGv+mcANkdUoyo5Wvblpno7tv5
JacgfqRRNx9jyIl2S1ldDprpwEklmJTMz5T6b+RMiHllGafR+PBRo+pkCj7q/Xd0Lotwkt1P7B20
bbwhuENXZv8PKQyZwkbzmqVU6ywNQy1+qTPCkJCDqyES3+sQcovfoWoiMujqIIBGWIbHImDWJZkK
NlQa359/3NatvHlGld929r5oBAfNLM6hoUk3daFm5Dsg7mTZFWw2bI2HZhId4QUGUOj5Y5XsOdqz
D5qm2tJ418c5diseRdVWmiGhJGv8LVTMelChCNu+1mNgz8f1VlwrRI12iNedQVudQWHZmh3ArosN
H1z9K6wLmKkE0cq9dsHKkMwp29jdG3kfRZJQXip7joOuHYUCyl7RffHEYARm1tB/UIXn0gAH3FhB
G2A1wcYmsXZ6khr7bkJZyt70USLfkDcd/lT1orshS/bhsdsC1ABngDhMEMxwNMpZastPvb6noxfU
+oNBUns9w3p/M7/BZjY3+JAq7mDX53pvoX9xslHhQPJjRpfBhmCnP6QLZOOFz9Bv8mvTfuVVD2+a
0Q37T1PqDfzxY0aVtCScn4JVI+LlbB88OWfL371uA8iCuoiuwbb/XEa8v19OUxM9enes4zJ+AUJq
iDFQXTLsD9IgW0xyQDDjrhRtl4QEU/76CR+yEwX0gHMXPKb5sVsMtfRUa8S4jSlL/lCD24AXv8A7
YKX446zkWdAZaWgtPe0Lc6AS+0YnSqDOBX8IgDWgl+QsMdxvt1XwwBdPRgY7t24UGGmNPr+2p8X5
p0gJDZpUsSPFaURsLL8cp80YAxOMHKneBbzJAgrQ2QxXlAfonsT6TxYdvg3uYx3cBC+0eStoYC9U
ntKVPwx+jNkgjzy2GfgtQk2xdYxnqoB6HZl3WR7nStR9syz8UvENUN1o6I5kV/bY/mVdPuf7gfdc
+QpnofS5eGTzRMdr7CKnVxcT2rUMAmROGNNJJ1h9lw7Cu3ib1mOMBa0ePhzeKEuUlIhs9fothFfX
sMoqW3uhKkdzVog4dt+uaIOP2Yzyor5TsagBkvKPkOxOMrg/s16B/L9ceLyDyChqlBr8zRK1NDi7
07eOJCF1rQIV239NlfYwOiBdPkOdl/HqjSIPUg6lUT4mN4byr44/JWRgnoIiQwJn2kCnNlcD69Pb
DRW63K5MyDSltfzTfyb5gmAMVwNYo0FOZYXAbFRD781nF0ux/6FyQtp0bymeFNNljr8an7ymauyb
s+xUg6k5tDthmcupmZK7tmkaeS19UjPfodVvmRMqfQRxRplR969haHnvVbciseh46/sVMcQIm5Yk
HRP2h0SV7McmFistpxqxMhhlSvIIOGPPPuz/bOU+VTJEZO5sYfKMXrkE+JhRKUd62OuEPMkb321p
v5jS1fTIfdtOVxV9fhVKAXacmAWpzhISf2zL8clrn0AOYcb5s39qAZwUmQuOtRkrfSVKTQIc2Ta/
mEg1vsQLD3i4IIwOvMpPaZBEMnY3pqlyVctuHTO4q8R5HbOBT5eDd//fkR7Yze2RxTKEEK4OFXtF
G3pKFRYthE8HItygWS5mA6N+jxwjW3nglKACtoRjpFJgPy8TbxCUP59ae4ksL/M6UVrWEUVYK0CP
fWaTlR8ceFKNQ5MJyCsrbzAO4P4v9Y2MKc17bxna11AwmeBR8yJK1HaVqV1Kkxh1f6RLqo2/VWd1
54BK5hcHTt0f3gsYlxBeUM/dNQhJz2pHP+9wBjuhgxZiTuTElqIPCzT7PRb6g4ESUtNoGTZvsbWJ
ANiItnZf4usMRcom8OWpRIGjWMfQn5RyWwFrU9btkHPbe6kSVcLMqb7xeOmHaMMMBGyYwo1HQCmU
oWsyTd1t/SDwtO7xce7X0kB0YIrZI3wjcEsKdKkGBiAua29sy9jKfxk+BwD+NRKahCq1w0SP4Rvq
mZoZXzHp08hUooTZqhDNxj57NbpJP9ky3BGukQV51YObUHN4ppldGDy2Tr69IiY1IXJnHi5/Wvtu
12iiJsjjol6RXHm+k+8STGAZHQT/eHnjPbZ2cb7upo4Ke2JQ85EgtJbervPYjRVX2y1ZBgtmlT20
FaSi79NFZb0JCcjp/Z/xIi9pHLvFUKNB+WDrEdP1KZ2HTriCdBAcka3KJkQaTkYyTaxZKk/Gsnm5
RInnzrv/znKI370Yon8VXUH8LrYOjBWj09vx14mRd7KjMzK2rUKwRAq8hdi3RDNkoJvUVKtTTxG1
PoZ0ivC+8fM8vERLO9f39w10Q2osZno7lm/KGiEkHqgp/PkeR81M5B/ju0RkhDOQLvkKQUn91Mnu
uHNglRD7YIqjGgQKnJL+m3jpTQcox/yTc5JH9f0BDbkHoprQj4AC2fS38wv02Nd1MYApt2DVyKNR
5DTwc+21beEeSohQygwOZx1d3/Sv1dXBFzy3bLd9eWqLHZ1ZsmrFe2Ou8rv5AqWfgt1DThuEp+WT
Zajl4VnIInvk27FbNbAHVBbr95Sq3Yj75gzff3Eq1ZRXHHQ4hQLD9ReHae+byNHi1B444wojTOSO
udG25ax6NfYW07Sq/NOHe1DUPm3XvNs6D9IZhKHihHJZhpq1Cyy2+1Cu3WMVKs1lJOw2UGguGOxb
SdnoJgQoYS2+NY32Qz12JsMzC7zfmuptXce/uE0nAjqehXmV6j8q0oBV8RyDlY1f0R/HvZipmMno
9mIXg0aMwhuOHqbL/HtY9CDnNBciMXgUnV+kN9VnxsB+y+umREmRxGjutjQy0Kx++AhI34vxqMEI
EBV9iRY04hcbnwZ+UWiXVJJpx5gPeiBYo0ogzRtrECMk0Bs7hacG5MD2/cEyIyHZNqsikf65FkoA
F94pVBa9OnFL8ulq/lGUAZl5T2AH7YXnlokAjBQADr3iaNn5DsOLeAPa3MzgFBRDNbEW97N0nysl
qx7KA6FljpiuJE8ELGvVjDkWW9+z5lp3liDkbUbm5BSDwSytQ80YHF6iV/3yBibgocVTP/rT2qy/
CPaABBDEReT+BGIHW6sCu+bujjQngs4Sp95Fta9oaAppgDuzaqhuQhW/hMrphJc7ggtqTFgC143i
0CtU+PqajYcXKQ21G+O4BNOJOm6/oosPe/VwqVILW5fU6CeblAoGbj9UuveDbsfqgU8O9ke7iyT9
D7aJY3bpH8BIQHX6o8ArfcWyT/3RLyg67JC0w3jGxk4sOLYt77/WCPEBuTypgoPoUe4N0QhfYW+A
3hJiC30s7q6jzcqzfV3hI540gpC1yIDoPh9QdN/OLzXNfE5AHCdhBK5heLQZj9s2pCAugUCwnkVa
6qBszZt8WUMGGkq0HrzeSWfXvr6/9CfmfauM1hQ8I6SlUyPH5CThOkKz9F/Jfs9RTvIUgiFnDFKF
Ss1YVfOAPAh3mHIy1j8Tqb5jQtnIQHxUf1BuaqxMOA6x+vixxPb1wqGogG9VMD6Ser/xsmTt1tIK
PLPrkB32D4pwvnd1/P9qNAWUT5wO6rP56LmcPwi8jw5uQLhr/zLEGpobwr0jp9y1VdOvudmCm9IF
uZ/MRg1UFyNVPB3qrTQTS87Hf6GI+DVVxbundDOSsHsZgBfvsgUOeJ7guwmxDXtEKuzUMBWPbMaJ
iXCstfimHceDAUWJYvw9ndv7mF/xDfB4O/0pNYO2u9VRRetW+80XgR3idq5TlRryH/7PYZBJQAbX
2DNtLnMJPjxPP+ZArd+39hzkpeQpvu6Dur4cavxfA6ef5/HW7H6b9Wy5Cd71oMzrg0PVubPGau2H
b7F6Y41IX/n5Pxt5t+whS21zOZo9riAXefiAOIxdKIPMZpXZ1lRLBSUOx2GxHrHsyPtJdfJ073gg
1SCirUXUkTQrg3Fsku8APFsPwkOplWKSnRl/gq/ZwnquIjA4jeNANKt3Jvq9hhT1ELEmsB2DmxR9
o92L1ppJrfB4N+rCPTKyr00pnhIov8TuC7ctlHg5IRANGr/9sBhplNwo0akLHPr0Cfpu32NwANsb
gp9HGHB2D5QodyVanQleV80Yn02rQGDD8b+WJ3mwAWM2evtD4OGMwJ2odL/cP1o5gTnb/0rKOtX4
nx5MOLE0byv9W4dCAaQKN2UjFEZ/1dx4q79z+FR/JkXTuO3eaixuDWeOIY2m6OuDHyggF7odbfoH
Svmpr6ae4wafhQmu+EykcDI213sDq4euXDgj59Msos6QddC7iU75UZ3J0pJPe5y6V8dSeCZbEFOJ
x5ne+TyG0OvAi5WawbTNINnCeajLg1I+ZPCoZEwuUI3haAqBoN0zVW/9IiFVK0tnKnlJJwomHayQ
zpRW16l8WihUJMl08q/rUy/A9Kb3xUIcW5w4/lFX+XON+B6a+ZGEi7sMU6evLm76eUOQRjvz2Zxq
uX/lFikPnqP1+5to469rqu9qGmUgYrGYdq2ybYTqt2NpD/KutA5DOIuPnaWw3XD8xV7cI/RxephX
WedGyZHLlJ3gGlRvQuTBoHDjGAawfHRTCpOYQSQ0ed3IG6mNdrcMk+aqgYSsEms3WJw1SrzjoR+l
4kPKr202hEtzeBH1GT2V9CHacyfvz9bzVwAxb8yR00sFZgQLaVoktZIA5myOQ0DSy9UW0LBslUpz
PZffUza+aGBDX9bV6Fw0XeUVepkMhI3bkJBaE4sHsookJErzsK02QgNUQ/IuS24JRfiRrMdgyjCF
GSh9uf77Ut8SEBuBBhoYFK7ZOHPnZFuYH2hXmqCzTm46XWWC6Jb29UTQUlet4e+Tpl43RY+KNLPq
Ozmx9ronQ5XDL2fws5+ukDmJ19hlSczGTKoYNT0iykrZL49QqBpb0rFzI0Tj0Nj/NIT+SHs3qtYo
/xp80oSh7H5tXar0t2Uco7s718d1VQNiRNPeBCmVrtvlxzmhL2/Q0BgsokciAY8N3ZS3QcVhlZ4S
AwXOVEmrNB9CWBhF7IH69kQY/WOP5FWJRi41wS7B5lYvldOlvVI+qkXXP4r/E8mrv74jysk4vDUH
jE9hbL0KMXSgRZqT+FUX8gnNKsQWa/K5Cnk3gPMZtkzBMphSd18xPFE+6AI7PWeVkFjr2FoBGiqq
AfKWEyYCZtZGR+I5eEpYAu61RiQwwyVo8uxvZ+wKtHl9T3qQmUlH9csIqWczNaJ+l/+vervBRrJz
oJt+O2uXHBqdDhqysAdsT97LT+7aEt4Ecsxvs6G/81KQIorPvIANfWr7TpGbpFQRNTWElFILiIuH
X3G6gKMWuv1Tv530X5eg5KNZOEI8IhEIpVuqCH//GpUxJSwjCfKhHqIV6V2rKO7R4yUIUDWlYlM4
YyKSZJqeMBQ760nUZ/stxnZYOXDkKhWFl7qy3A7cTiCjVlOZfEj+M6MciWzzj5X4C2+CGTXUjRgl
zm+wKhzc+d1CtTEA+SC7qh71HWAeCjF/kbF7HSrcy+icnP6LJfIQ1qwtzGra3i33RoxWlwQVoH0N
IVzdA+E3cAF4e1/HsvxffiQzDKgzJZwnkEZwyC2m9QlFSW+70v8ryIWZF/QFK5Xb6oCX+xHv0jnB
8mTe1g0u/QvYScg19J+HAWvrzgUTomrT9TyKHMyEKSKUzhx6J+cGqnkMsi8rUZsgR9QKWtLtyHG5
mdHCq1vUWXvnX1dkKx1iw38/2LI5yAN9qj4ltCnn7RPyIkcnZ5Nt4JYWvem/SCkTLSCQzQn15DXr
9mjqVn+YSuTfdVfF+y2Mde4mvolzR0MQ4nTRN6XC0tCUNscHb/Zlqu1/kdkFyZOHO3IjzYo8k1p0
Z3Fg0HhyuJ4+LgiyAzC6jgSuS2+RN29ChW3KPxG7v+yJY/01IgNLmsg1PHRxLXABOf8CLPhHH0Ow
mGbcEhNWUbXQHRjobz6rY3NQwMVbL04inXitiTmJY9z3eggrA771roWEVc6QkdUfH7FsOW2sibcC
oi9Mtd1fBO8gxu62sNQigOCz+cDGehgRM3sCpU2fTTwPG+c+jemZff9nHPR3+BhP0+inFJEejO8u
J17xQVK1hQYnPo5qsU7rchdK3peITCDmTkL5o2OwFbGe2qB+uMcWQ6ZbDWZ1VhIwXBFWyvqbBZAL
9HN/CeoZyce8bc1Nb/QspG3xHujUv4qnJ1WAR1lJXELNz4BniqpoGE0fV85EJhbJY14YFljccmLu
eIieXdEFyYNknYcvwZSneiY4ZxqXMgZ44utSI+ErZBoH2cFGsJ2V3OYfsl6Syfvy3ESCUN+74sgt
KC53ND8ap34+gN2tevGgAh9/D5T9fMk4oahSq+73pwD/9ibnUWMBG5LGjUqb4N1AlZgFd+jj1guu
0NgnXNzRqD91ynndxEXUQQl1YI5ApovXQaI0XoG/KBzzjiYCa3ByvYXuWL5/7X7sZ3WPspTTWTTc
Wb7VqYPDFO3E8lU+YbfH3X4K2bNEQ80Fk+1qiP7897mnCBhDpdmxW/lOvOXMNqdw3eYHwGQ8vsKd
AEEQ59b8CmOjzRhUx9tt2CpkRqpg2bpNVPso2GXNrm5I4wlnLayZhnF++TbU7mcyDDz8nFxH9y+g
HacCYtAaER9kcBpW9rVVAJZjdgbXTdJ8mpjmDbXX8xKWYauzbl37NFPb9/UV6Yh8Dl5i1tssP1s8
G99Rmfx3SBpRXCiHcCNxFSLB/Vy/j26DN6AanPRPwUH5aAvD0sGkYHAGTCcoPGyyzkAHIiHtOkzM
E5TB2aK+Ce/l70sY6v3n9W75ukBuI6snn6Zj4RD9Ocil8VDOiPcAPlqi0Oa41PpoF77s3pzH229E
+Axij4P7iHKToJTPrTB295EWdASvT3kuHE8sr1rH6Oxpz+TMU7IAcifLwlmwBrwiFJvYWx+4QkE5
XdqbA5bSLiB68VCgDotqVYun66ZsHo89Vs7OcA9sqnY16yIfxjFZxBWheJwo1tXGAb7q8kGSns6h
i2rlSF7QGuGERS6QfNfcWuNRVv9oi831btO8iMngjn5UlCT40M+iDHFJGIgJkgCYednp2UzfDyUi
H9hZ6if4dkCa8osxl9XvxzSzaN/n9lSgGuO/btgyS2EEEs+6+cRpoQ/FTRfM9P6vPDX+nEe/zAZV
mNZvlYj/tGlll1EAo4Wojlk8adW0lWVryxEk+xHz3jB0di8DWSh+cVS8auebMuxMpU17nHmWOcsQ
yH5hj9pv0yF6awNJ70KE3XzAXd76y+wcEK/odHBOdgP2CMIaXvInDQs/4Ur6P2xGNX3lxoZLGi+J
TTu0tlb3LAdDFwXZ992o+Wx8Qx5BLs37IO/gnFeMyaL2Zfr8oej827fMYlTzshS3UZ0RJigd80K2
PTiXOLMJE+I5A0kdMnUDorLIq114b0/3+ODdce2X3/Wa14TR//kiMYaW4+aE5G4YJur6CuLx2EIm
eKSrxLnkwm6Pvxqn0pnSr/j+6rpb1NiVsFITYHAtliLFZgEA8//QQabS0WFH3yBxlu4C5o2vv1Up
3O5Uu4qPjwZtpeL2+35aZAr1oY4fm4xJwpmk2V7rHgZa+URGH36IfzOjbbP9rFzXiyirjU5oV+QC
i35wU46adXt56NQ8T5BtprLRMD8R1cAp+38//yE9PX4oOqdKTj1cDbRG53062Z1DHhWxvAmeBk9F
nMZasK46CbhZI51lB3kI/Fjdod5kcC/nFVRfnml4y+zoKcM+cibOQC/xz9f74H6de91hMzKAaTZw
V34t3EbV3povPsoxCrMxPHZ/by5M8s/yM5FCWaW9I0TqlGkhe1aIEYMxMW5oWNyJtzptQR2DvdCi
xuC/VduCMTRxvU+Q+BBXwAKhibLVzNXHjb6R7hbIY3qvvWwse4uid+H/UnsktAgYHTzjDnvPwKNt
WJegJG1i5eNBOn6UhME1mVGffHc1Aj8yp3wQMG5GjdbcT6ORq/a7seqEpQHY2PP2A3wZyhHO9ttX
vjPiNPAKKG3jEzWJzBs/nKjOQj9JDbj669cffISXmZXhFoZJjbaE8DmS+MfH7BkNphqXmHq7MiyJ
Bp6womxc9PRsPSfs/+pyZNmkxKcrhXmywZjDLMMmOPM0lXMlRbIMGT1WL5nnVbVeT7rNPnRDrJBg
fL+abbS/PMhn0W6PXCKWiz+kwVTbECoLw5u354jr2+jMbB5NeIUeV9qHKOX4BLm6cCeb5YeB+HGq
bmOEExO9YU8aZNwoHUJo4Wjecdma6eVBvfKoKJiRc5FIVMc37al3D3xl7yepixqlIX2Tyyb9fvja
Pkr5MoFwtpP0aM2DWk6diR5tu1oORKhU7beQUkjXBC6d7OqKHYJC5IKA/X/KgQpGmuRngGBZEzwO
vJeqG0jNdHeIkzduoGJPZt37mHYPgJcYA+HWCZ4f/yC4AfU7NGKJLzs7gSXtqtLgKEHTcSF4KKeU
CuKTf8p3j9UpYbT7BfEr74X8XsCZ6gP9U7YEKKPfQhQOE3h8OkTXt5zIjSAQmX8f2Dm30dux/5IG
tqV2ZMTrDvswJznUMWpkAiWZFDi83SXBinbYWvXAvWqHydxKsUujE687yr8r1U8I+J+SdEi2j+dM
elEsXKJdA1LWqDD6DnMXBHP8wZahM/9C7wUTZK9SY/BHzv/rLJ++BWUu12fa1vW9erU3PED9T+bm
h4Dj9TkqTsOQcVOkJII0uso3aWCqKzSlcWMGGE8FHX9TY5v0pGRiN7jlbHdvCoSy95zhRGk4c378
1pXK/0wTwhJ2PQ0RqiXnF/58gumONHmChVYk86D84tDIkgL5SfD1m2edqTw7RFTPQ/kkJZOoAoNF
DGesu6rQ+dzfCOMX1aVZjBl7RLT2Hl61Zz78CAukh4LAsmgKES2rBdf4AnBFNZ+BT/N1VCdXmoYH
oyf4nMuWTRKWsM3LZgw6O3njLYjR0e5J2l2Ul/qYbeO/EZc+NauIzd6zw0obyCusS9N0abphAcbE
rBkkoXNm1rdneMvuIqHybPpcyy+E3lwTgDFuD9F3nHn+z7nmjdscnm18KWCDhNcJ+qYBAoWe2v6E
+rOD5oK9jU7IuBG5/BJUjHmXC/oXDZflBzQ2uwANbpVDBudwYH/spJVUoDYfdK9z9da1W4ZZstuD
gOV7HuTz8vzbR70zqS1lGy5jLlJRxMAxlcSJKqXo8KcGn8KeKOsO4gm0IZcGdABqz9olZdRSzOVn
rc+a68N31tTYnu4uSxy1QjfNHULS5Po1y2GlS0vOhn/II7m4OVzMJ7v02fgU+rmH5wGKd74Xu4Xk
LVM76CD60/5UdQfjg0d90dM9eyQvL26wC7XSP3638f89CiqR1fq3cAYmhV0ZD9ZgqB6bFExwhwhM
1AFlOSITvNn3mhDpXkShqON1YRI9nMx4OPWdVVzzrtJt7xze79vGsU1syphY28XkeWdAj0kXXvWN
0/g1EuNJdMkAOIrFcwNhqkORUrnce/oHTnRur7ekbfHR3CKFMTEdFStQp7wjXxbAUMlAa85vmlpN
x6ddJ9Ffn59OkPUma4SE7aVhevggkyfcWlgLXzZhIKORtp5cROOL6U22Pt9obOSeX476xtQ+m5YX
Oihz2isBcB3qVLo5MoyBxlXfQD+TDJ65fXYMSU0okKGJdl0YbHO40uWcas4WAplDs/WU57fjr1Zb
VFMgX34/qckSutMdz8//w2ja7BV5Jzh2oxtQ5Byzz8E6Go1YtYPFOT4P7l+EC5ZEslZ814X1wj9h
KdPjNepyB82wA78/z0/T1vrPUkNKY2IAwemc9pFhtjsh1Uly8LYAhZgsORezi1WFE3gfUELQ3Akd
tDSrPf7Zl1XoiHKJhK5aYmvv6GSyVh25MtratVmQ8VkofouMkW6aNDmIy8I4vYTzMBXg0mzjJmO8
QsSkrS9c0XgZmt+eegISTVo+pl1y0Np1Z66V2YMAGiF+OD+FzbIFjG6vMQQtDkfHN0kXhaXOjb4i
srRflgOwlf0Bk3/cAKfiXWQ/GsKCWuUUK+neDQvuDt75HeA1i5KEEJmGdyem0kAwS/byn9AQcuGe
ij7/af0B+fsnh0xa8ZpeR0CfAEpx+Gb/M4f0tDdBfhzWE3fYzScdDGuTYPstpXKr+pJ8iPnYMHn+
voI+BLAhUDCzztPQB7DA26LI4qYdwrdtNzWtaSnwMGBrj7SufpsR0ptQxxzGsyU/8+T07U0dxOiH
lznFHW24oE+nEOh6jvqLlmZWkSUARCU9D0F87l8RGfrtXaijbCRUVRs7iGnm+qijkA8q74IbcFRu
U5OfN4QbtmAIDaBSWiWJNaqr1UvkwWj2HXImN1TJtppLU6Hk0dbX9/zxelFoqgBFBVXsDllfy9Fw
GOz+4bjcXR2TJyo+wSrxeCtPLOOaivkW2Jw3H6J+TuFdLLKr8jNZjU+qHgJdnS2vPYkvWT/0oGp9
ghsV/3Pn0FC0obwv7Ku7oYT/42suxekrQM1nZV+HXqhTLHwWVFQiRL6Q6gWKtsyzBPp38ZLiatbs
j8spdtxBUuLx5N/RaYiWikitCWsgQXYpAxOpS6ONVMIVO1/ebzfT3dP7YJC2Za/aUS7xrHgajGnd
og/M+r9SYkJRFHM+xm8CFmxkG4jh4+r//MiC9aDHwN75V+HHsiFQCGLtynFChPgj9yFnnvNhNvRO
EOHLuntZT0xDRpheIZO6tVGWq2tm8q+VBKwKM0ks3WX1ZkP/DgIVIxpfwTnSQiS9shOxP1r0Cr52
tlbeb9RQKHEyiJGCX4oMM1CdH8fXTnXskJOmZlcr4aa6eqBs+mt7/KxZXnOIDCdKoFsPIcoHHk3M
O65eZ43gmjihFpq9bzR3aGcL6GkCl/WDIRKkYakiAvAw1LezGQbMF8iZ1oaCmPCfuIncyiA2dFSI
956+xRxyGGcSAmniB8ZuP7eafbt5Veakl9rqXnI+x1m3QcIMfmvbLgqIb7AhsBVpgAEoxKMye8Ci
+uJYwOSo+2nxYkQQYXCMz57tQzvhfQR+HjekVh3kMhUunUF4vjQ/0hHcxUdalafgrkrlzQU21mfm
eA0FGj05U6DKDNpP2TlkgDwDNI0pmZ43Ilw9JXwPi9D3cLfkSeJiYrlr7lByhzKy0T2H6dYdsT1A
oraOFbhoj9nGoBNqJTQPlKRIKvErxUtr3mk7CC13/605UufAYP8BSNlify/VfuNdkLcBzyAuoL6X
y2L74d+KjoBkO0U3Od+724ZCPcYQNzlwokl0sbjBrd+OKySb7X/G3ETpwD6aUcLAtSP072AYNq3j
LWBeFVKItdKZul7corRb3+Oxu24k161Q52c6m3ldq3XmHhVpGREsefdP9Cqn769veFIg+C+TLdOk
JggGNKaAa0g4jWjPzzY9Ylp+eL0dpt/APFMZ6Iu6lGPKhBo3sQYBmI1hbJDx2ywPaGRPt/6qxCeO
QarK1fkSmurGsuSvCCvsRv5krHVkA70oNmoXgDLmsg5RGMjHNzaGcLFmyinAfPsikc7HDo8baJi1
BUIln0Jb4/emluoMz/v47rQmz770215sQ3YKXpAbuTBsPt3+WLkFS51d+u5uMdFhlynjVQ/eISl9
8ZkOUVSk+e6Ece9EqLjQFPcS6pQkBbB5FiLwSAK+VXGUDI3Fbx/13hFxzvPsN5i+yiPlBt/fo1DJ
+yik6VL6ehOxPJYu4eaew9aa9FnBq83RHeI+Af2KxUPNlp8TQfnneLrZZHxbrhlclyAEOhcivzvO
NMCRIrQJkZ1VPMAo4AxUn5kkcfrRfZDUc7utbzGM3qu1A5koiY0wlwacJH+TKaVq9nWoBgpkEQ/P
L3/41vDM46KdvIGOnzewZzW/8ECP9MjGCbLrZgN195T++i7cYbdsGbWij7lRX4CweSiNB5OwVHTD
FsRNVVBuvwgZ6FsVFsLMgM+1NxxYf6habw1CWUWJphnLh19IaLDJKCcxo5kv1WiiYiumeobbhOeQ
c5+hnxypOOD8vwPPGz7m5CIN4kPZfiUvIsE2abHlDP4CXMmf25DJQRReTW4qEAzS5V8qXXRRclY6
mxmXwQShjXbvVx04tve8ZiOZtX7wkfPFypT03cxjLJEknF5OIEaYFYge7OoTxyVdWGkRPH3Ek99y
YS1AMChPVqzOHzDmecSbBFDGX7vi41Y13ihMBe4U2LO5iCjgTR6Rfq7HqH87rEcYHx2JFANDuXin
ZAa2CP/is2GODkS0lmi7L+02yOpejUF6OruCNo+tkW+yWaUMhvmodv7C3mhtXDREh+x+ZDZNQiKC
7QBRvQ5zJJOIA9ZizNJ8HGkxNNa4BEFmFAEfDFDznNTZMxW64OTTDxnIwSH12RqnohKzpFDQ7k5g
avyW8xc7Exw5/3aG5BaJxRHHRM5u4E31d80PH+6PSA+qVQ9rjAfKMpiJgl7AohjzgNKNUvA5NOOW
h/XKF8TB/UKJ0mzMy2gOhxl2auni5Z7Z6t7kU+0nf18JnJaUoN+3RAm7YIsFAPwnwrGXya4EHx6t
UnGzZTAvFGtqPMb/z4JjV2VAJVGDCT/fn+RsREF2rZ3u6CRNFU9ibxjbmOQ9+Hu/v/hbjOOLiBNB
Pnc/e8AnJLo1KYKp0v9LrHdiJROqHcYeMWQXjksbCFzd8upK49Hmfff0cHXeYLkgPrACaiCUlWC1
21FYqXs9Ye0GK9ovEDSP2NfcKkYQW8gnyzXpMRfBtZTVqYWZrgIcqRZRYKY3xWLleEDZ+mibEgta
ZY34+sHCmRqVzpzXtQOBRW7Bbdk11VCi3uJlcq/DM54njB61ogFAStOk7RqDqNKj9ucsA9o60HvR
VktfYSWs5Jko2MEecBF+DG1n9WTXEC51qcrvb6QaB6/XHG2oiS7h/34tYll0QJjYGinZ9mR+JdPT
VnhlJIb8wcB6T2wiUwczJPx1KD+UZj5S46iibmKQPoXezPzVeZdxC6DJp+nGuXrQt6gQrhbnp3GI
X3QmpNtIwhnXFWM8SeHG/OPhUv/m4lDImTvj+QcAckEk/DdMfI4/yNjLXnTK3IaCkuZly25wWiAL
7I1mvKcnVwAvoP+XRe6s0NGOe6gR7+x8vXc7q6pgFEpBfKA0AX6Pg/xsmofKmNd9e66lxYrz7R6h
KLstgN4+jQn4IS4yyxmgitYRDVTvFMqc7T4B0vsO77NpLGfYGvQGRsZWerMJRz3L7/dAtXU03smr
Zntle6L0HRElrBYUGqF+bk/IUogbss+eqMdRn4tWPFqzKMcgXBFZ1IE5Jwlcmdx23f4nkDsEdhCt
uJYKYgaaQdl/FI1s/qpaDJlxU+BfQSjpNdL92xKRMWKh8pZt4uxnU9iYnb43RET611R4jODH+LKf
CY0waBQxs0uQZnaNqgUFgvorCuXWi9A2dAzA9fqVYhwSV9pI72uSMLXfXFHjvVGB5oLlRc3VPbIw
z1E/HKius93iNaLWdlHjArN1rUsgHwwKKwiXOShPkbF2en2xv8q3luG4OaVKLfeNQUyX+LgiKeEd
3TRg8zKWr+VFH2Qe3tDlbNiuwg5MX5S+euykWcGTfb/wKGS3rU0nesuz7DzgmeuAk/1eVIcgh4ex
uGa4N2JrmfpEZHRtakl0rPOQyPW/1PJTkw3KgXMe6hdrUANDkMYbibzlatsu5VaiHVX5PVB68suQ
2WbvEG68NCfP1iR3Fm72t9HdyceAnRltgXg1nM/8GU3MjfAQFc2N16AriZc5iL2L0SgZn8vQ1rkQ
XbXY/qYcJ0Nz1kyEWf4u8AK3pl0Xgs8vRbX6vwhEREeAFm+r0B+Ip1lOrRY5KU5IjOCbh150tY68
tx9tBu7lDvaQ2s0WEVdhbplXzX/QudxdOpzWHd2c9wObNCKNpJ39d0den4oa4Ei/zk0aEcbWu7gg
DRIFm1KZD2NVIC7u5B8P4svBGu0T5jUcTWNvQimvsI7arSuBYnpMxOStX17b/ov6om2LK1gd3gCZ
G3X9r30uhMyk91brQY3DM3pUQ7hKKBFxUCznfDYajL+VzNDBFtGhz+KAG3FWZ9PeKwRP7+h6NCUj
s+IDI3vCfwf5/ejAPGv9+KDRF4FpQSNQOKpaQ/PnjcZ7B5k+McY90gn2uAXWKnO7bVghSiv3gDbM
t9oBT9vbEhtqCP2wQBf9fUCHzF4zRvKKzUL7a82/oIhvjDn8UDQ2n9jou2GR723C68x7CdR6C70Z
PUMVqpfTUi1WUpUIC4gNE9eb0M/EugDHBN3IYG0YwCMda+I9ELvtyXrD4OKlJawMINOiHZahILkx
HQa4kr8ZIfts9vcvZtx49mBqOrTZ1IiJrIx0sywgrKxl0N63lK4Va6Vn6s3QmEOBuGH3Zc+/h/Uf
G1Q7rpZwAnMhkR9okmp5Bb7EePZCHeL8ENKyLSoNvYq8JuZNqQqS6RQPIk7HLGHmvqbuqAH32krX
aF+5briHBaqPwYyC4Nx/aMpegPQJllbpYxC6ziQNb+V8QEjySPChOo6xkQUoyrmmvDYspF3q5H1+
QZ+gdevOK0jDJLpitTn7HF5YoGjBc8VcTm02N3hQbKEmdxJSDh266vBIDCqx3AEDKrKrQuuxPCbY
X4fTg61wmBfUZFTOf11mt4ViJDa0rvtfFNn2pbK7XxggwxLR29HIQWOW69IMVs9dnNs5NTO7M0Kv
pWYiRDR7nyrcppUuqwDpUXP/PjKo61kjRemBKxijcux+qjX5igDfz0rw/wMK7cnuG9U+6loXdsyR
yrOOShLjo4MFpGPTwT1TB9RlqAhS5bPv0FbsFcJk5qGWUmNYS+34H4HnNpSzP0ixoMcBbBZLS0cW
6OOpWbCeE0rZ1ik4nxqp+EK+zmBf98abHjOH08UjzixNYN7lRsO3JJR/0+QfmG8RDTRmHIz1kH6x
1IByB4k7gJI1ARGm4O96Spt6Cn+gh63An8yTvvRppluhd6ryxivadpPpaSmjf53OBTuR5L8swT9c
BJVK30tJmQFjV5GI5Nw92bkpf7swlMlmXgIrXmstrKyrRiWZTp1vApuS/pJP/+ZV9c7S1UO8LU2j
Xq/EoMwDVdBP/UQXIixUmlP/qtFdlmQ6DSPnM7uU2S6kMvRdGPnamBobe2yiDOqwNKXeCKTXSZY8
liyuiewDQoWCCc40NWI0qPD2W6GRIPTkjNSov5x9qy4W7Cp/hK2Oa1zXJWkO45X8LK/pjFouLU/1
UtUtWi8+Y6zYekGL0NVYcrlz/28EEwau903ZyyjdtIViDju9c5nJ7fFcFYjU+LwzrSwoPgrFESc7
R6wHDFDAJgW/8+odZFcyWINPOcuumiL4NBDmBm36stw/6Fo4rp8U9/R0teVbpWwHCZX5I6jnxlY/
Xcb1zyMxaeE4W4nPr9gsNrzK0tpPYDVJjSNQMwwYuqUT2Dz5fTrC9YXoMSYm6OMMtooQSm7H8R3A
C5raTXza9N5UD5Gnw9+031Ty6beX2kQZKbp9XfPnikGTzhscr3gzVl1j4Pw+83iu/yoj6V4Y/67P
zVpu9s1wAFwC+TAmsKIYrRXc8eGx86r0jrIOoPAqUfv2ZrviPvAdx8gT20vt9Hpu4P5WLsato2nd
+/W8ir8KBw6ZutxLAy4ohzsP8wyAXdjuThqlmSRkpzNU5lsj029KAE9O08BrJO/z7eMQkuiKF7VY
o+Y2SrOQVRDTcVqzDG9ds22R8YAg4OkHjTw+nESDL9CpSZjUGhbh5u0/1AfTMPUllroHxaj4KPrR
k8ANDYLHUJ+a7mVyTk9pZFoBkq4jMN2g+7joiQuGrYPXKniG3LoVM25NcAw5QVykMdy5tyXpqRFB
eQ+DxmjMRvpwZmBy/Eak0GgZg+9Aouspcbq4tiqmvt9ZEfPSfpWjUShcKFOT2skpdc9xOHlcRRqG
6UaY9+fMz8r3iT0zkrfyKDhQSKbyOmQEGKp8kfusobpZSvWqk3ZvDadHeN4tA6oeJLT/dw4y3sAV
vt5IylMWqed48ZIIN+4wPzoxhNGm1J6N/t7d8XHnjBJtT+33Ot7uQIt9leYw/6aLHh9dAhZio+iR
Pm7o7dHYHOmsNbNCIjHawmcA/j38avOa1tgPpO1gMMRRaFz5O1WnadeqTuLQ1kJh3iueiSgkV4qS
gY8nKq01NYdaeK97NRjQbcaXDG/AXGDCbyPMcDHgqsQuICVHKEA2qQeeQt87Odyk4VnPkVkobJAe
yqD81lwDvMP/v5YW1Q+WY8ZDS4femn3QKIn270zucMlLxdNJUCNvSpFQS2X1WnNRY8OuQGu2pwJp
hqvm5WLFMwu9LYIEggVQA5QpEyxeWx320eQkftjNhIrbY8wscLTs8NM3DD9Ja+2V9tvllcqp2A8/
Zor2XyrmVWk/2ye2LQ4yTMKEFqC9pYXCI+j72eaaChCT7K+2sBJciAoYm/hNcOo70danMfABQOoL
+Fu5yVm88/b39CJ/FCQiKvYr6lf+AEdqBNaztjfieXWtvk1tXNjWQCUR774fyLn/Bc55KE4vjPcE
Jwpa6LLbE+28vnvlJGsm/Rg1kKJb2pK/GgdKJPO3mYCKkBzMQgNG4ZvSgwjPcoEMNNYVtLsQ1Tbz
P+7COzM4axdcK+64pGqFNlw0xnBZJivcoKTeCXrRJuvbOiCKZjqKmBH8WGkxDQ0WsRW8o3lEoFGt
uE2YOSxh37PAig7VrYm3kpc/GZnIPss5UqSTWIRCumKj3xJIzt19cDQsVz5KjbtXpsF02iucauJa
KVHZ6krQwdrYlw1zCJxMJMcrb5/8fGBCPU/USmYXpH5zB8tL/dOZ6BmNktY2aotnC3ZBx0fM97hj
lzBG1GOKq8KJKnE4tWSnU/oyrGXMmwAijmHrtcNV9ypMpCHKO9OA+t3P2NyV0LE+6D4XPnUduGP1
l2os4ecJgNjtK39A6Wb6vtSL9YZdb4hXquWFt8AYktqxcp5F6ZQSciZMrpWKvtEqSgW34j8G0NQV
BH5GSLr/vFws9l2j6aIWclUxDC5U2mJPXIbIn6ZDarIdb6n8oXHlK4UpPLjOMU7odtUn0uKYYjEi
IhMI6eY9htGLtYmPbWNK82+LLVdH4ngblgr8U/ztKxy5+eUCOfVBA4dJIRoJ6beR/9QRK7FMC6Dw
mtMH0p+CGXAQfNMO15nRCZLu/hJAHu+k7ie6l8pfEoBRN4p3ChzvxU18EubDHcbs8FHXW3cdXfXB
8TPDfuDUJKOzy9hVozVPES1dYgXMfnXuw6Xb/ju4DNBjubO4Grl2N++8kbhb3b9sAMRjV1F3Mote
1ACjLuYPdY5rVNmBLVsH/xgDV8ICyIXm56PrmgiiaRyaEKUhmKP28zgzSRUHqRxDBing5nQPgxIB
jiMKjEmaaK7T6NBbRNHwGy4ntS6GkuoCpso8XFBtxdq9JiUgtzEaA+GNUefWlVpiJDORCNbNObi6
Vts1AspOBok8bSvX/Ik82DKMwSf12SPJLYKksbdIqFwabuSw84jZO9j0cJJuq0Znu+CYR74onLFC
SFvM5KWukpvr2END1r/ZwWwcn13603GHvwpQU5bmNmlKvBvxLvVo7bab74I4UGSlMUrWDjdsc9mp
t+auGCc2NEZ+avTyKYnPSfNSRhGquRExiWkorY3nia0mq36zoW2+Sf1Z3kSwbKdkx7ZFoHpiadKy
Kwt0lYqKXiW+mgyF85FGJ7ivyDkv90W8EE4DOuJDPnPeVNPFx/5H8SVNt4aPnQrjDHBpVKySIob2
HhI18UVxXR8ham5wYYs4buHf/fZ6yBkn8Gnj1ZFADOZc8qR/q3Jcob04zO/5rzd7zuw6YeSsEZpc
8IQ7mWuxPc7tujC2ujmGBgNu6TWkbbGOf4wx7/fHpkzb7ZEbOH6pBJrBGVvT5v0SlMVsJGloUCjf
Dw5uYuVTk9/R8A3kXRkx2XrOODk8sNODkwFJ63XzbuYZDJOFIA9QO6FwUYfEIEtEEx00I7MOr86o
JDjUZdCKian9vqpPmPLw8LNFeYTrg5F+6Fikn9077Xf309aq+jx2gZ7fA0ytgtXXuZyDL5G7MBkl
lwpoIOHbaSDMNSWYvuo+sHs3m1w7PNmcjaCqktRlFZ0bMmlxxYvXCStP8AuSEVMJPFoGZOZ4tc+q
yr0KuMlUwT/2aFHHvuMW19oJAbFJ/Hu8CwzYIEOb736pKzHavdD+a+LhCPRkrqdNLHI07FMJ/9R2
7LKubOUu8KdkPpY8mlqdfZucLxzbHJu7nJuLLglauFIBSFuoUREvPKwoDItWOxORdU6h6ow22ZkV
P0hGwAbw+ot3wlGTnBYGCFktMJ8iigqYEGsO9ffqSHRnN6I71D7fSR0/RFU9qq9+VIs7G0xaEguq
C/2FadNaiAQSos2k4uJLoNKjmKPfAYZaTkdqf1sS8LbZwdm4qkVbVcoGmPiSL52RR4T4+rt1GoKM
6gbkx8mThtaCS5SfOA+WoBPOH20weZHywWCTJVTndx5TYjNu74QmpIy2wfZHxAgL9flbqfJ5x3WY
vmJkoIwGRTQ0jRqZ/tP6rA42lOVws4KMutI8er6BmiA1434UIKvuKJqmszGtD31ByBLxnPzLbPRX
+EQIL6KypQdcENaUqlCrS8g1M92Gr98RxlCobXJ1x/2EEyEFMA4GNTIhmc4t2r597TBr2Wwpmyyn
RxwW895DxW4+GifeVJDprbkZi3vucdzqPTco0bIwnu0n4C3uZOnohNa8RH0sbqLJpclatrNCovni
GSW8QVU2/07QYbtNQ3tersGkSeIgnVQPzuM7BoGk2nEEW9AwzmHfEkHzxK1DTR6Bjvk44ZZNvf95
5jeBvvVo8Qzf/QKRyMk12pSKjujJWZZvtzTIbLnB8WTc3fSWU1JbzmtnU+gNmecIS4jZmudsl63z
GwbwnjYNIU5o5hhLfTAZrgNWaK5WAYrP8NaKELLlNJasLsaL3OuEL27lm5oEyI6JFhRvTg5UfM07
cvEbJbwCngA583dz2ODacNnR6Owp/S8MqTJip+NjbgjAq60wy5G5M99gy1e3vgadUSx++8RUpszU
5jfR0lzEy6tyAegiJnHcLDCLk5FkW84qzOENqhmSznjtnvEX9AfNkUXi0F8gIskq214cfc8FFxJ1
Q3gg9Lip7KVU7BwNzt2HbeqJ+pgbTsPdtmTp3t0EipUy6KNXmoQQlwpJFGSbcQqCPFJP/BtmhEQD
/SzcAKMScXbWO3RwJKd9VEoPsBo9jAuoIl+lHteGp1L7mrCH+s+r7WWXBODbxCzJ9qm/Nw3C4rLk
Nyjohi1TmvgqCIY5lZ7UlhWWVYLNv7qKe9W+IhDb0zabkP8ERsgqqVHqjykxf888/zKWSL9uL0p9
1Ik/j9MpP3EvAILs0SU3r5uUpiJJuwOStCTFDJqaKWIYC0cJX0N6uLYX2LK2bh98axdTLYqIb66p
o3q1rSGw44ZKEH2/5OCddm8yiHC0nhiNx63SeG5d7QGKM+cUvlfM1mXnsGvjMkb2n/E6KblL+gp1
5zPFFIh6yGaWEcEOYyHC9pACPtHxPvOhnOnfoMEegk31kDFtnR5I47owhL82el/ddRFSd1eXbyNJ
dVhIXbGfytbphh3Hg9hKAKAjizPYClNGU1+ykyEUC/lYVS7j2As1YG+G5hvvJuBpkGgbIbVFyl8W
VLc9IRySANaIhP11uebDeGTHSoV3aRn7cerM/2drK9B/3+Sh8z0zqysLiL5Ur2szCBZG9j1fvbv/
QlSeVsuq9lXUU0cP4XXQj9jz8813F38Z5f/Q4Z5FiYHl/H+/KcK28JBHufhH8q65YEAaAfj424vl
6LC4yP3ucBLK9EVPvF+SEH4mABtV711Vah7stOGycCWszu3RJzNwF40Iwfhy1viZ4p8l6jggGJ3J
iMw302g4yFxhDrFCuhW1GxBqL/TxCVFDPAnUekzGxfug83/gPq2PVdzJQeCH+znm4kDrXS9gnOOl
oc2Fgn9wrDZ8+Sah0Uy+GvtvxELiEihVjagnC77Dyitow+EY79CbPCoObRwc1BT9qaT9xvGy97+u
L1J0Av9SSGXg4ZDLyeTnocTY8P5vLm5vIj8k4Z4yFM/qVR/J8tfs9eNz3IuyoDPWwZGjiRrTKPRf
INjXDrsNO9Qr/xCzNbGuquYuQW9o3JzZDcETG3ZMzAkNnT+7E+Lz/FAnn7bzPuDW3ELFzMvi95nF
pKJsbtdjTkGVnqa4wm8ZxktF5D8cLTn0S5nJybFuC3I5IKDeN/V5ZHYw1Ew1c6BgVjZRDPproHAI
QVInEH0mbrekkeesIniiX27Z2JWqjIYCycVCeqKatCE6bXZ286dyhgaTA+fc40gw+giwgLrdg7QQ
uTf4NTbxiv/e/B5C6OTlVT2PREefWnIjRVSfsni8128s9xy1pe1u4LGrwGwIEVhxCLowZBHtBBeC
ZTl5BCZ7wUuEHPsHSx35LJfbwuQOAtxIObIKXTLtkynyJw4w5UPmP0s4uPWbMmtsW20EP07eZrVq
U4KJ4GQgqoj5Je1f20rO96JxeLkOOdrye0t8/bSfuyzwfoMlX87Nh2YRu7rfLSxWfU0pzEuDcHGn
TycPMpt22kjE84YMmM8u5PzydO9BEPfYYkef3FMlF/drtwUKMQSaDDsERj9+b4IdVTYGnRtOATlK
VOBO23aZ0suJNbQQXne+glb4N903r4hYDfdQVqAq5j5zOjGgJSd4xnnITpFWGN+3AznvwtUNh/sY
8MIvA3gx70QVNtVHmm2Shq2ozS3GzQK8wjj0jvVYqyI4uEuoBwJaQ/Szz6b9pYl8fEItNIr6RWaB
elahSgoCtQVQYgg5rGwofP1YzAK9FueepCWNoEXaKMHCrYAMt87i3iNxD37R0BF+S5i+WTM0lkNg
Uhd7cR+zf99jiJ2l0CAp/gyoZbq+4fnNjc6MWpivwIncVZcaZ19Goec4NL+dAXVi8XQxOb7O+aUx
c/WdYPFnpZratGtoUifVNnO7Mt7rdfQ3JLpa75QZYL3C23DsIfNGZT78tL0CVZ+iDyaJMzFeJ66M
f/izqRTDTOS5XGCT32d4nV5Q4x1ClOPfV1+ItLEVFyNd5yCwBHegcghZjEeersLuKDJq4mBRHngn
ilTGTBAtAT20aLirKYeSnR82T2jkl026ZSbjAeeRDHFpzT0aJFjaME2oZDRHsYLXq6zLz+TyWVn2
Xa3FjF+8LlqVJLpCr7Ewvl+7RQXFf69WJXdv2uoeqdzwqeGqK5QdbbPXaRqCSa0h5vW85VFFK8qT
9H5+LMcsBP3ZiDS693C1BPS9pptQDT1CM9USCdUyb7GHaH2NlZWz6QSAlad4wiQAzxqwzKsX1Tsg
LvpUa7bZnc6IQxYhUHZUEUJVC9ClqTIKmLiW2g+FviYNDQnaV+vV9qfbCAR9IhHF/ckEp9feG/rF
wMKrwOCPmCzpIfV5XddCCt3pKqG3IAWCfYHtTrK3j79z0cV57QtpezRLW47E+GF12vsHlIvp17oY
nsJ6n1TRf9hy7CXqVg0b3R1XMPTqrAa3j4PKMFPd/ePnz7FLKwSjmQ7qAYl1feP8Z/GgewWzlXAL
VQvXGWJ1fW6ewUQI3MrFK8SnKfdztil0rzlj4UeiO04iNskJNm9nUT4KPMZKUAZkxwEpGxP6KVO3
CCvUpkzF6s2CUxtqNTJb0BM043MoYn75Hb0ikUhjuEarnQG4nXF7FKMxQzSWwG4oc0dq7MZsPBs6
clREyuNArls6aNn592z3660XpYFscrdqIv7iGcIS357f5FByaSiO5xHoSKhWfobhZ+ewMfy/qW9k
9g5ott7TPEZRqos3lUguK6jGWSdd/kY0GId3J3lVgu9hXrgFJyfwLNDM9D1WQKBtY+QnTbcLBU3+
OZImNeb+irs/veSPkBXteVoiwCJXG/ywsf619B3piTH2kpNFHMDHM3CD3dPwVXlZ/d/mJTnOnlnA
ostA4jzBUNaHjNHr4aTcW8DaBxK8j6YS+a50bio/BzFPqWiAzCFPFPZdU+phJ8FpgsP6nZW2OC81
Sd/LUTPrKjlkct5I90Xo3WTtQSJ4zwemMBbnkINJm9/eYz3KupKXFQmX1Znc0CnkyQL5IsPPc95D
5Q0uF0X8kMtxitHQF5dxCl4GsXSgSuSGsuxEP9+Hl2KfnzsxqNKhEGDbkJlXk19QraKgZGNEf3rJ
OgiRNmCXk0MxOy0y7zF92k6Qb/no1TnG40DLrmKFnJ1ugtA6iOEzdP+wMRKxcDsvNzNByqh1wXY+
sZ2pe+SGyvP2OLdJkwL6DN4LLRKDUhJQqnxSEGnJo2jHL1rVlcG7IznH8+A9/Uy6AsSjOaY+HmhJ
KV78zg7rt4yDSPwdVz12mNSoAa175n8t2iElYtL4jPLSG9WXeg5LTpNeVwQLHd1MLz3nqLx95kLz
k1P53fGmBw1K/r3AzFfgCCf+fq5Q25XfxTYeh9kSZxFDs3qCD6PxQf0wi080zhuBx1mSiHTEl5cE
YAA8rbUvWe34Nnh9OAFPehJTU3fZidyEAP7QOl4Hued4KMaw70fG9K4gM7jc3dmPMEhiWvjsJHfo
p+7YvtIw673yaknwk4yq3nHdcpdjbJXJ971zROk3JMPnpT+6pYXqZJCALg7qHKl5doG/ZFzTVCmp
VJd0wu4YKW07/jwHBtRoM5AVqy51a8NHmppKx+51nOSpQ3pRHyHquWv+hUhfv4gcH4VEEq0ynVPG
0sbY4sNmtmeRs/zpi8coWwEDDqy7+xT6YUlvey4K+NQyYqZabnom6QAWT9LBgo9cRTxXiQ4p+uvX
20igvHphiYhJja01sUqnQvR6S8kxPfw07ghsOo7bo/CaUZkflUKaCCRqSPVMf6+bfGzMCidvptBD
Mxw0pt2LcMpJZ5ZLsutV7UmI4gyBNHJGW3CCojoVNlkM81WkGxJhFyirsSFvOzDZg6fGMXaPuXid
WOevWkT58aFDhmZyo6CM70yvF51R5U5RRqxasQpocjuBtMBreN7u0mXNIK6lMmubw3T2RwG2Ht9d
GYguC/mTqj586nuWMLurSi0nWPh7DX351bZ82ZEyUsMRJ6RvUMMKJ68b6VJVbtySIupju9mocCxt
BzoDlZIXo4GwwwnQ+OoSNJ6I5MP7p4rUsWcQvLSdnEdNAc3bWQjBYZEG5qqpb1lP3N9uqYjA9FL6
KHBwHwQ2QK95jqWSfBJbalCNI9HEbdWNjo5VRrhgkL+1gyDZdgKRdn/rsXJDFnXMjx++oEkwEUr+
ysC6yngifSGYcyzvhesrDeTxmINQys1b+gtytuYXDVyTio96ohKu0SoK+tsf83P98aTakvAX0nOu
2D28Yk372SA2e73zwPgKV0eihiDO9DUIU6OefKIXIAV7fpFs54mpkOfhUEQ/p8MWqAJ1ri3++r37
v1rtGwHjakY6T0g11x4DtX5Jc/3BSIYpYZ6aObhBXCP0EhZ04H/gbm8TK+bU28W6FGS7pn6YcnIt
f+wuLNzxw0pX8AfGAkL/PgyGK1/4HZFRtEtahqxN4lZHAnQdO/PMloq8AFZQfzmtYQJHqXrGtE6A
6rLM3e5dh2ed0AGUumlWLwMtVnWQ6M5hXd5eZAlN3BiLJ3kh27wvoZLnVKrobcxpsHkQQaqpiyJJ
Wh8Y5bGBYb4o0uu2kfRPwz83cy2Q+uPCGkjsAliPg6wHiq74cT5pbUqWN7ODikR3Ld79XdX/r8B2
5oJwFvc0pGYm2IRgVYDfG0vllnPaDB3LJ0fpZ9OvI66hUVBWua2b/GAyN21V5YrW+IrIGvI/QS8F
ABKgVO0YB+iUKSZi1x27TwGY2OMv0J0ikm3d9R5bMSwqMYZzcd6ZZw9IBe+ugeQJpoSh2fxUqpsy
htGF376Af7RMWLw6TtU/ezDr5uB1o4VPQpyEaYEhZ+biu1yKWqZEEMwhfhW3m9Wq7czSnv8BJnW/
U/FjLQZ6cCU8sdnvPKVIkxY/ZM3xWGVjoXiwszaFPM/czeqUJPbay4gKiboE4H4NAv+fESBtLBA9
f1mJG5MXncbqDQvbXUDfjQJp4mTGrclZWNvf8iEKPoB8gLpE2Sso98yCyRSu5ILrgsr6+mSZbz+t
3dYp49XbuVSnaDkmvjt8EWpGQGOtY9sVKMzjs5aH6T46+4YG08n5omo3KC54shSr431qzlDrqAWI
2uOaMXCjYK7VYlJ4efkw6K8Y1rK/tK5zrnTghhdhwSTdLQzDWc9fvq4dTH+rmXgQIH/qmuk6RoMD
aK1+RD1aru4Ct4JfBL0haqWd9TjAAz2vYPi9DDcMeoRRRbG6DH0N/A4Xp14Qaf5xQIhO/7gDYUWn
TZfXd/RENhXdlu5iZGg2EJDEs8QhD89GJ6PDgefZurKh09HInzkZgq0Uz+H7MezTepE97fnaYLl8
f7Vyr9zomuO1VBRMQEsiWfUHUuGWZ4iQ5Vm2Xr3ecPA85inGbWuHKQA1alVJMkaSMiSbJaK5jqAR
wYO4jImnHvuREPxx+IC9C1Q5juhKdAAH9aa2RwxSF6NFDMVCwchypnp3llg2WZJeVO0vmdq0GXm4
E8P7zGlnhGZ8irFymriUiHy4orWXPo2aesPIXHx7keOMKLQLm9/JBWu93t7dZ22Uw/cfGYC51UlZ
a98bVPskqWtIitzeBpXMrGCoSCDGmAh/kpi/Aa1rmsQELvlYvTf7A3RrUG5KzzPzqCFmdHYcAjr4
BvzSMA3YcgLxOzIMm5bO6PxU0u1yh/FH987KZIpj7VU4I+FwQO9ixJt6QdpewGiZxdMYc20mEh5Z
Edy1EGo1IM/XDDInlQ+m+ltHDFNUSKHO2B3JH0h3zBiv/Sv3YQyb1XfZOhWB9guw5yzeQjUtG5IC
B9W5GrFA5lErLgswzNH7nnYV/4Wpx646yw4y+XMmMcVzvTqBbRKtDxO8tNGlfN3sJGRZ7s9KXCgS
GFT7qL273t/9NYlLTFvwObppyV3UeEQI5d+BQ57A4fVyvGe7mlqI/Md5bDsw1lxGPJ5439nSVdtJ
PWAxNFauQkJt9wy+c1NHhWVL8tnc4LkhT0wSgz/HFUfIYDUwf09Ep3u25w7bsMd+tyCjLgdCKmW0
Tm6puQPtk2P6zn3eogmGLqRfCvvn/jOTqZSaHasleMQJ55YUTBcTPi/CapF/fublDWET3Kiow0tp
VZXUsJOQgHuBDFOEAOfxx/td9WHDaHHeNdSunlgZLw3yMgV+baXKW7mK07wnmKk29zU6MyySewzG
pErE1emQIEhX1iT4URWyXMEskORJrXgJ33MFgPzVy2GdpHNWUdANondHC1DivTTYqU/iIUyEXiMb
66OnR/sLmrD0/8+UEXIr6ep1UTvNNRkoZ2WFlWpsBm4bGFOrtE56WF3WgswakxFdwz+SQzXAehBm
sWYJinhy5XO8RMcpe+6SiKRzxFSEWxZPI2Mpoq5ppCmZQ+lYKGo7/kpJ3nV+q/Yv9fb3DqASRFtR
BCXLNM4ad6tbzMuBuMxxwlEsj0PrnIsKwc1Odf8VBAYC7VYA6vwAG5DajRKSQl3n9mc6lFyDq2h9
esfsBTawZqOdOGRsLVfd703CSSnTnF+Qm8cxE4UQmaCU1H+PSEWaP2jWK9yNCiUGw/giJKqfUfbq
2t7dTobGWG8e3RPYlfOq2lwoGc1rIf/YfeFCKgRFRLUXrGXGx6Vjnz3tZoDkq+//iX39JipzUhk1
uBCz6Dy1r/YshKzARwYYMvFDMpGzvLZiILFhOACJFzzpZrrPkf8hoBKWPX2cmINiDR60f3DQMlAY
Uwt0j6dOp1R5d9JXBBMfMW9eIxIy0FwJqdKOsKWbB5Ax7uwi/HGovbzE5QLgz7j3flbuhjbiLR/x
K+g1NcN6v5muKsmYkoLsTELo24+Sa7+yRSi42LEpUGUEbNFk5Tl3Rh8+5sKqLIC61YrzMT06xyYt
auSKZ+KOKVf70rQwlR01PZyvonVzrg8nWoLGAXL3QVRCGE752Ptp8K7m9jxo2W5hjS5lbCXRx40H
cZ5FGHifxW2EwkvWK7ROMQttZzUxnKzGirBWuFeTGSToi+CfHnOAJuxahxu3cWogFBGLFibaauPs
MtW7/iMTKHnLBWT/NW/bOzdxPLzmXXpM/Cj6Axe1VBJoEWwG3abeVzIA9wYqdod8hmfbLMmZlP1X
Dwv48wVpNUxGcq535vnNIsxbUHDqKyyLday/FbqyMxiVU9GXsjtjhgseWoB1h+bwK6lf7eoVEzlx
YTnGZ3d3stiq5xcM4NrFDAGzK7LRPuKnYtiDPbjLTAGNQy3g8DgFr+/q0TpsOPUen1BFaTUkqfuh
OA8fOX0MekfDWLEMGuTbzQMqbiBkFVhsn6qfv97gBxf7P7DGRUKRI3Gr13EH6881apmEL+7guf/g
ydQ5mxsKHgAwFVhh8BsBgE+j0OID5yROM8W12R9mo6a02/KkFBCwGtpbxCVHOPVP32Ws/0Jn5PKu
4NUKz3vttUBxvsoaYjCMjqj4TRp1tXnbdFVib7GsbGmNVpAVOAyztzaDLmmLymm91EixvuF+MMdA
G3Iu2IZffYbC6DVDq9kZyK9yhRAweHfJExvt7POtoWniS+smQUyllsC04dJ1VrAisVW9PoeYfoaT
jjKRwD0/YRDtFCtrEMAor8SkK/5MQ8veowoSmNz2hPNUc0+BqtiyNaVpfxWufEKAZzaec1yRH3Hb
5kna+SL/dRvNiTImeT9vRhxZ6KCZZScOJUliuaapIIJbEtCWFTsBxWjf07xG+Hmh4lCjL4u+3C2k
4ajYMcQzVbJWncbfMFKPrEiIcxJlfK+4V+mAeqW4Iuj8YEhqcZsMRV9DYSxIYYqaKmCGzEEKNF1L
3Eos3LewGvmZhEJb+e7OmC1WkNslrps9FoKsnvaQyCreH0lZVoR3GLgIdjnRpq2k68h0bEUm6IOW
IFTvSvMtpJAM+n3+3r+PelZZEfGoqJYdybUUPGY241ACVYJHo+jJEqJlgiBczzcGagXfNYyzpJnz
jGXNp/UoWC+MeasI3h45UiZxj7wZwBtT9UQ/dj4lV8cgUrsOZIKb8SZEzd4j8QRSccs3ExGlRzFT
XUbmF4OmHKWqGFv97mhZBKh+3rUNTUfjSm24YYVJuHwfsTrGI2wjW5CnP4zQcXrxmCmV+1s+b6Mq
W/O1HW8cIv+G0PvRIZCtgpK6MEPUtNIJl+EriK+9Bk75htg8I734mTs8wqxHprCoYStSZLZakYu+
8dH97Z9YmDnNWQE/x0RR2wvx5P333g1EfIMwb+E9sBWMfriEdr0lGQBgIQJWr6SEmt27sMGsL9G+
rI4I7P8+/zxmcDoYSGRq/r1EnAiXqpE7WYyhrbs4ZrY9VJsG0hO4t9zgSyI7DSj29jGGwI/dOYmh
stwtRR8Ogtr8pq7PYmifvX0pT/jgu69/HCca3W6KbkzWi9WDdjx3I3yz2/5UhZKBRmPp5KoojV/D
vFsOBqw8eGjQe1m1ouOiKfnxXeRVJ0okR0jsfP27JiGs7qQX7auFD07CtuEPtEvBNdTx7wHia86Q
NJ70nG+Z1hb424N8254BlNJaDRINggogq8yxSzKNUPIUz5JPC6A3JM3TJxEHexGaNzaNZmg7SPD4
5Ksfsa2+qGworQaaEd42+o2oxAR5cJ6Lv1sZJuVpc30C0uqVawc+8m4yTS5MuKBfm84R1rt6v63c
N+S18e+uUqEZ7g3xOPUZHbeoUhIM4DP/ZiX1CvsXDdPby1mOFMzD1TMKHN0syu/p3bPrcgC7UJor
x2CHCHvGQ0Hgy897/65zSxXsvONiAI7sCwPQB0X7mUyGj80+oxJnRISmYZwUFLO9SdhYdPKzR+xn
Tfuy9AQFSmpB0uHAhcv7XRlEecKF6YUwKHmRyQBRSqNQaU3FOgAOGYyptxY44Wqo5WkTIe6bUyap
acF8Uiz9uKbw6MHjWH8xuKJ2Gas8flXnZkosTZD02nnR8Nz6YWkS0dQlNcbsqBc80Onr7uA2WEwS
AxijnQA4kmcVCIXqJxmYGqcl1Q9lAXkrDOs8Pi4AuWj2PwWlWF4WZoTXK6aUhh8yNTCrLQNgNZnp
lJFkYbKPKUvtOlhWKohUpGVXYTWYb2eNucufhQFrjpk6siwagZmC8FCD9a9my2aJS9l5XPrrqrUh
fc/CJwyGbxarEOpLtywuA2HpOFgyg9mnfmZ+mfSG14kkaTGjpfiMNDh+Rxgt+pCBbTRWA6//lCz+
eGRJvgUQd1jr8Djcs/5EOgH3f2UqBMIpHMFvAak9t48oPThVulMcQLfHYc7vqxZRNoPAHHXlfLzk
6kUCGEmPaHVu1wSYM+vfhOLA+lmQGCq/Tck7gzFdCKok64r8iKEP4zx1FTWtvI5+wiNxBJN+Pekg
DKDDwDHHesDT/fUFcOAo/A9SgEoona9FVMW4kgUiTrSUQLQO4Yc7DcqERofyiQr1DTAUPJRQp+oO
NzyUqXSXLUYTJcPlkss7jIhqGhIHXi9HejTIMCK/IyenCJ0EHEb3sgNZ2ZB0HjW48EXWIeAIu+Ng
PPRMnLRt8nSlkodPZ4KDKBgNlbZusszs4UnK3tW257d9a5LvmBo5EsXNuwDbUtDyz8C2qU+dBG98
Jr+OvbVPp5zLiE54oLtJN4Ji6NrlGlwzW7YKUu00bUw4hm9UAja2pD/aozr4rQo4pXZUtJnA8AvI
MzWS9Jvr7FJlLZQbaudr57Ig5wapoZNkUsIPc/c6anFxI4VS1lf22M+VSBH5KFcI9bs3CUKJUoLh
VvuoFxgbhpwbHYyesTf6nObTVtAIt3bei6I7xT996+RmRnY+o6MqdN5fA7/yPRqS6juNVE0oE7so
LNXkAsyyP7zB52zNyXenTQmjZcnAzcJfqSsbJVPTrNaf+bNXaEzMqoibyi950UKWSZpDnlKEMg9x
/YQfYR+2SdhnquXkylzL313rskkxIsGoe4zVEvLFyamqAc7hzmQ5WtHXehJPxcS/FmyyTodMLMIi
n1bo8cCKTIzMucJYJ7wrTc1uTXToyn0MECKtVAT3p6cfdrvC8QiOE3X92LzatMVPfP2HEddtrgCd
BUFKBYofGr1QcDCW0FWBY117wDf3IgC8JC2FWZEtmWslIQGI8W1QnZ2d9LQweJo6idtxMPtZEfZa
5b+7UGSSeNt6lJCsdnYzCkLeFEqL3iAvkhYgs1T6L7RYLCZYDI4fxFxKMo1hecpJKm6RoUntrFIB
s4OTOQlk/Aey2Xj31nNwnFmsO08WaddVRoVhf6d4SMjXh7uZKC+9gJFz8LfRZ3NoaroaIKx1j7b5
OmSRd5owjYmXQzsg3RtOiJ3WZdUHDdg5902niXrq1QJqhiSPeo0iYjw0Y8hyLbKlLC2g8d+/Ig3c
s1s0o+NQTTZKBOFVVSrI+enSorTWQwGPRwX2fTCa2u4hUtmXwYYIU4LLodiWJEWES2aF3Z/t4vb9
fl6LP8tbFrzuUjr5Dy4VHCMRh5gVlt91MUaEFxn9bq2qxJrg3wrGxeyhTVmVe5t0rtPrkVUJ1Z9g
sFP+An4RJktxpTz4N8hYeFUfe6u1VIPkoIHOuvTNqdJ0NwCuY5PV0AQ5MT3SjkhyUsMHz61TSbNd
iQ56p/RabvdOtxE5TT1iOCjtTOUNAG6C3SN1N4/k7dPhobk5IIAii5KEHp4G/D60FaL5deFH+SmC
lx68IquNetHmpzgzQh8ix3TxuAAcTSpwbTmOoDM/fnPjO8iGuuXZjbrvKoozCfZZHKJn43UCE7CY
J/kOiPuvC1hjlBC49vbvB9DrGvg7JWHAylYAiDZzydvWOfzRGdATIhEKIZOk7bC6Ht95iELF7zW0
ScAiG7CnsWOT5N1n5ORkiN34suWpGdLnaRga1RF32ECa/qrjYphim8jwVCgGLhamL9iruLVAGvFr
e0EdefVwDJEz8XI13RwE+1mCb7hlkIwOIpzBTSpEnqJSgCWRNact30RQKblzVC6vr76NK+mhXFK8
NOgjmvxfYiW9H+5ll2ICdS9LjmOmCZAEGCaEIRIUuUdnJRUALzq4AyQ8CBhgRjp5XugGyirDwxv/
qPWngIHgSlwxo1bM71ik4PYA8ltWzEP6fovLGv2StQFu6+uU/j8TukIpd5oVQjg9wmsHZy/WrUq5
6o9I2B2TaIZFH4s5m8BS3COszf2Iebe7BXQLZ0h+XIKH20eekJxJSf6eaIfrW0D/XsFJmbVIT22m
u5n8msWYg/0etvQH4+MduNbJFL1C3xXk89z2cYzZSWhCeBK7/y4bTqCp9oXqLha33k6exH9P9Ts2
qY9k5cvnY9ouvJ6pflQGgwhpxE1LRMP67Sr591hXzrRAPIb98yWHYaUwWCBnhsxWnb2wtufKkkFk
WNIZvDdJX2von60/g44V7p4ZZV8oqGho6mYCOeilvdw7hNqowsRP4LxMpKvjT4iT7Jh1sKjr/qG1
0sqZSaw1dH9cJ5VRHiUWcwZp0DF0lx3abs+k7C2qn9Xgiki71DtwPmRT5VgCruNP8H9uNYxVgM5I
q3QF1hufz4+g93zF+b3cDBVS1qXPNZuP63XqetH0TdH1I8xelBjhJHq1iCiJ6zNFk8kjtzS97jdL
gy+YXJ7pf6uVzgGT9aVBtWoJeKIz5h79grYh/fFSOZpi0L/hL6BIhOG4vOvN8DGPU9JTxYrsLJXC
vPDIQ44Omlm1wg43OdTHHpip0FtOm8ph19LhnrwCg3U4XEiCF820riiRRn6mo3kDdfyD0DN58nTC
+07k7x0sqE6E4w0JF7z2Z8zFX/6D74pu06MAv032771KP8RsIfuAJHdPVZOZIUwbE1YFfPp1cEal
nkbku1R13GTZtRGP+fulTgwvhGM5A5Ly2LiCDCZnLjpgdY/zcP4vjrYwnh5vpQfqBVAR8/DbEcws
EiDPptiDDjbjpqmJRwTzj1F4qQbT9LA9rB5LUG3FhPz85KeT4g9c/hEfEciPon01FEKRkdJM681/
csJEkOLxlvdAV6ndIIqCGy/NmCc0RP8oOl41p3+I2DJyxRPu0ZJr6OD54gldUQJpUrmGWP0cqORW
sied/TD/lIYIfK3sf+Iwk7dAjfAiSWdsLCzfYruVspH2PltzsNVJ5Em4+zQGVRF94XWT8lo32IfS
d4osYFpMgjRaWQdIMBc6lHJlmV4hhmjcuFcdO8lXnNCz6ihAmb6cJ8n/Uq3lICeY/XMGVJmcltaF
ybFSsuQDASGv3MRuykEJm34Wjv3Q9MBrc5lFYlpXQ0iyMs6Fa4LaB0Wc5FGhUGSODxdPeIIxNfQN
s4SixYCJYxIq5q1FUUPz8e6fR6ZZTxUw0cRGUN8fRwwUjecx1fzeDkzmwcZ/ks3w1TtRuVm2pVNj
kl4nZFA89aVqE8KsiVfYBXqXsXB2eXXqZNl2g80xPxHWZ3y1i9JKQn+QPbq5rAAsctmBdcHirHZ2
gd3cA0Isc9ofO7djh8K6OBcd7fFJMiJ4OL/TpXVpYWCmyw5I8mWvXACLuSqRjP2vgNMRCVXuqxSZ
IuS/ViOeFJd9y+PUE7IGNSSx2AODXad1Wj5uGin3cAtXgF3hbiNNzlP6gZNpMe/+JpKps7xcE3Dj
g8sOOBxtqt+DK1PEerA6/MTxlbImoLGU4HQgbYp7rh2Z9oe3cfJrWRFqAMAgQ/guRngRya4+p85s
GYGL0pVXK4vvJ+XaFP33v0jFjhC3n4UwcTpGrMi1hcok75jVW7OOx5xXmhC9oFxwVsxWPnmKUGIf
yTySeYCRxBOlenzeonwmAF7+rWu5IDpo2Z3uulnAQXFCl+KXZw6FaEft/+qZTvX9ZFURoLoPR+5X
bXyXu3hFEp/X8txyNR0ShLAr2+roqgzfSt+gxtXk58LNqnoAZDMfKAQg1+XA4BjdpeagAPzq5OnM
TivEaiMdlu5MSiAxiLajV1nXBn11CTsmkZHu76GY5OSrjSUWWGZKLd4EjVLq1nJ2JLKTsSbLGGFg
R3aGYdb3MPw6Z+ZsqAFY4V/zbdAA86cEYE1hFIB/70nYwIUKgLPbIXZyuYsxr5aZkcZLdYn2INQw
ZAOTFDsBDQrIflWZpdoHEQ1KIPQRelStcV/HEbjtP+nihRouGvZn95TVU6dq5P32SgmYhFFZ7cNq
9v4S9DtPlV9U7l4ZydQBdMtHaBcS9LS3LHKa1jCEvmqZvvxd+HAUYTxKn/LVGg1fw4rQs0mSMA4i
FdwijiFu3LucYYsFcQ9IWqnD8KmWoHQv8BZ+2l1JJPdlBL2P6rkiIa1XtjefC2URtzpsljRqhk9d
y8qGIDMdMkCZZXcydgXU4FI3cCKLw4k3awG8PBqRxrVIWCocPGPpifa5zw7Pw0LtOHHaOSjSNK5H
WSTbk4SD1tiyrABDQHEsApmmLX6nIxqiE2EDUbfsCP9ZDTDyaIeRKZitGEsa33wXvi04Np2Fw+U7
psAsyQEOJo7bmJrHIdHqdCYpY2Q4SxQ/Cqw1VyAyHog/eYbTWoJHnOxPViMWSgpDMoaq8FL66CAd
t/pMJRw1rKVEvDxgSiHgeriErWM7qoHR615fE7wZvQxMdM5qOtleudfcCPZ8pUCPB5ZARMQ1Fhc0
4sPJy/9n4WPQ74Pi83I9+QYVm5gCV4LWYdEQzi2wAELQo2L0dVtVRbne/AYUsOeHaS7keQ0Ycn6d
PtwZcXtO5UzJhGpw6jIW2QCzQUs0ZJfwaicaIeGyEnes4nUvkFbYmbyO5IAfLdhAL7L061zX9lAP
RB1SGKn9+kardVQFWADS6aUqV5L9LQx+YUHA6gMgEBPSVuRX76bPJLYEkFe/ZaVC/UKOpHHIpF/2
tN7jnlhKB02+JztGLbnle4imPnmHY6W5ccqKC5t5eV8ZzzSaoU25vcxBSkb7E9zqMTy2sY/F67TX
k64xYxX8BE2Ppd4+y5pPTLDxkZpRbO6VHbj90JNA/8/PdlS2IkuagUVR0eT4GZ4WHkXcVvy9Uu1f
1YF7hdTaPV1k+adXoy2M1gHzBnlNLk2Fzzt6TtK/Ee92Rx4v6IJHlsUapZn0XIdDaINSaD0WEQEm
bQDhT2IxpDtOilKa5FVG0EXmQ4jSuY1F5D+7TXSZayMODv7I0yCBZeBLdTRalKWfuD0dlQbXcLMe
pD1OuBbCM2XXrBJoF3rVQOqOiLZJaobzevjye3KvOmy9/Xvqw2TCYvRpuXYGjPF+ElqPkKABtjb7
2oEm14m3aUryEKLGbkDas9W7SOpDYLT8yOFvPvT6IB1SdQHZTgSKYvjDaky/ulJ0FKFvYstwKwMx
+Dzn2l/hhns0QzugUbhsJkuhMzeVoHIDTGZgYvpHu2MgkHQSCX1A04PpsTZwqC72nlaNP9p3WY2R
Ppo1kHChmoXLa4X5V2mHGG8hUxuMmdTNYMjmxVmGxzE7+XJeBaXU2GhXaTmlwwfoNGxDhvv6i5CS
ZSWqxSHjP3KwzO2fHYlULGorWZ4U1B5KN+1yIto5frwapwTf8HfhfpHEvgIBg93DkMHZ4xXOi6UY
w3+tNzLsyq9MiEjq2k7bHS5mJgKWl15BNNldR+8yvnRbqIFE/c08vI0Jb6k/F0HserjkNmAkquUL
PohD//sW3ALItQwSWQxChH4YhvyGGacyoUy9uJnP/Ru1WsMS02PBfPEKVPLm7odz93+ZpBIq9N6t
0kyDCO8OA4kKuVUb3zVS8jSfYCjEy99CaaooAoDqZePki1MSFdN6DlcRqx+oQU0OteUGVO+bRM7f
pAoL9LwtGdEMTCSNi2eKtwa3oxXCnCjnsQUjkBFxb5A8qoqwCdJqW71SotTkCx7d8dGLixTEIQBV
l45NsJ99wKQ6OqDwNLr9jjuBn84bTiLgdNcGNOFbtNN4bk3wsSgGbhgl5tra7O9YRKe0Vtn7M9fj
RVrJ4Nm7xvIOVGSnEbfmx+wdT+dwgBX0T2vNF5Ht0VKXsroztrTYrKnb2TmnUhmB8FLhy5/I23GK
YAHkKAgC4/4eHJG+qBosYrOktKNvaCDH06GyCKNCrFBf46Q2racvBSE0fnLwtw/4QDDRGwpECt0I
+Eh5bN8qjnyOwYHaNQgMJ0uzwgF8+Ny/VZwaMsJmDL8X46+hqj37+bWEzNyHrF8GACyfkK1pBsSD
e6Cc6jW3z9Ij0xtoInsJXM9ShGvtpaO4TZqlxjJQ0t3t8Mazar2A2OzQ3RloabknDK94chd4WhKU
BCU7CqzVwTMF0gNCUpWYVm/MlS3hm1tByT9W6dlvdEK+bdBg+CJzq0A9ilFrgEfdNaOgb1wASj5A
eseYqYr2gkVl4X2pgqyvapcouFohEArmLDAECi+0xtDPuYpdmk89vO5Kn1fzXHKJlmXDIYDn5Ygh
miStUqa2PFatRtyxCHcBCIodUqfozUOdBSV5jwNsLdIeOyeG1D4vEgtPFoXBIdQtaVplTf9VfxKJ
58qe7L4nbGG2qzdhHoTwgs8IfLv6hq2J63/O0YTN2QesN7ws7YXasCYBBnAjPc+BRcdJm/I7mM50
OLI7B0DOwvwnNi0jEDv2TTezxCrK8i3hjBH5etrg67CYRKem5cp6gCMVHNRlgXLw0VCRzM5y9AUM
JjEk/wOotrhH9CZcRdF5w7QWO40Oz72M3+fB5NAk0u+luDFrahvfC9Tm08mroPD2cPI/PKhH7f+W
xwqK3Gk7DASHpCpX2o76jrDrtSbWrrd7M/0Oh+rt36Mz6mjxRjHoCF+0C2U4cx6xDwOMyUbX8rXh
ZLk3pyqxFE7WvNPE2+oZY/iDEyvoFeI4uPVTkbDTKLXu51ZrSjn+9L0ixORqOkB/V5zKeqvxKyQY
Ceeo1rkCFFV0vtihUTikdnQqElDchNQhiDBD2/6CV/cA5kqSa1GFrBnkc8YlcZwQnZkJWMvZ29ez
W9rRGWs0krNjJrMHNmZK+RbQsPvmISIooepHmIwtsFI1zPf7XVwgAvtX1fS/JA7DyNiq3dpGxg8h
aS8XWe7QOHd9QxQAFWLTTBq3xlqI7M8ft70uTQMFuB0LcQym+fBsP8CXhSFdtp3l5HCegDjYyQ7V
TZ5COkrLApM7U0AUk8LQKrLEwyU15pU1M3UhuhwjuC8qvt3dntGDAKBhCaU/dRc9wOaHHRSs2pHh
Me5lvzs+6Lf+QhLQf3Ta1+zwgkcj5jlFxIwrpoxjQu31WDqTA3lCEckCDt+lywKfPzgvoUMt/h42
chLVfNsoPLAnsMAKEWRQJexxtUS/EvzM/6wrMgK82Zd7ipzdPUe9MUUF2RYXo+TbOYkh2BnHJxYX
qLE8i4OXGFbaCijJCIXTsSr21NUpXbsKM6EqmTM8sWycenc5XT2RT1+gjzNyTpmVOiDMQYd8o9XS
aXdzIyPL4JF2gt/IzwN8ndqR1p2sYQ8BLWQditpLZ7wrFtdwkdnl9xAlpcXu6ZLzijyFoaqCVSrL
LzmLCWFeTd+a7JZOpeLRDccH1h6gZ/xmTF8fJPHYROFEWusdQZLKBY+VV3TVTk/51vEWtCr7wvdj
uUqsI+c+TXzkV7n7Pwhe5gOwBjwRoRz63QvfeOtJl+22gv2vpY8ZOqCi+jmQ17ljqs15WeiCOgmu
9WXHa1goyXP8P046Dd3x4avrGLSysx9vjjgzRTlOPgJeiL0S0hMMKewryTyMH8T9Yule9qipTuqJ
8jcdRFXjBhZl1SLmav7LOGbRyzbHSpLZ1990YmIaJZzBab6fEEzz/IPjV7S2/bvY3Iw99e8D8FKw
6/I5PnmK/31xxGN2hh0FPAUJCY6xgj+vnTWBXYlGPFbkVjWGpCZZLT1Tld3RsaFfSdDf8o7oK/lN
b4XpksxiY/d+gUFO+sWOXVOAiHYM+HRyfk79AufUnvlvrQhCe4hHCAVW4vhexLohmvXxOSe969Tv
mooVBaw8pHB7bC58UI8annCBtjGNjr99ZkFKwI8gZk5vGo7s0dGDERQReTQy7FRaCnYjNs9cHL4c
qwROFzkry91dMYxTa/90aswA75+ZCPL7rrnrVxENAqbe/wH++VngZ5gLbY7d3FkEeYQYlow6NdK4
yYVK5UvH8moIa+r7CS8YCdaa8jJZ7h0f62Nmk+6zw2gAxExpUhSWq7DJ5SOorV0leB0iFdF5q5eq
xq6QbPiTGhYY6zeRhG/GZHC/KX2CpaJSl9jk2sertu23NE+l5Dj41poPHVgTRlI62Vs6HQPFXN/J
MhP0BCTCWgLCuIkC4MeuUOInMliKv/KPjnHtBH+cIyZ+JFqkC2MDHRWgWWQmKO9G6v2Zhzk4ZBDk
7AYlLEbQp9g93L9E4vqDv2yterlxG/ylJ5/2aRY6ycuafXY2pqFCkebMPY+pC4QleZ8O/JPVHZqf
BsKyQqOiq1xPCsMtAY1jB1kyzqYwKwcoXIxSumbKNtdDEX8regTq8xEtWT7gUuI7qEwmFjRN/BD0
3jiApm2vagmZKHCsHLX5YPX8kN3d/BawBBbiA3xk747fkGjjGBvUrtZ5Nm7+8sbXuAXj6SUH6Wcm
BgQiE+8aQ7AkUgOJwiCr1sZ9qLx9F0/uvkFhEMG4gwGyYcZ9UpEsXqSJmJjsbB5h0kKWGfRPqTMc
sDV3+7mKDWeaVLoXWSnpuscNreVpaZ/eYUEdvKnvbUg/WYOYbAtNG0QRlIVsYzRh/YpVpVjBAKK8
mmPEvicBTsvLh9nnGPufmV9W7aMnD72Oruat2GJxv316QZ0C7LfXsN4hxoWAWxA/YI8Bqp7XPi8I
EQ8z/41xNrKdSeVNhLum2lR4IYK8a9I7XEny34rnC3cl3KXlUa7DaBO4Qs+GV60fmHDQwQ3bT//L
gXGDg4G0uefZhROZ0p3G4qkwVmIezox42SM6fGQkQC46GNRscLg+90y7z+js2GI690vzfVe+VMLy
o1LiQzTd7zlvHTKBKvT9xx+7nRFv+6KcP8UX9KCX7+y/j/tmUMD4TrjGWtyTsuLOUbKEJM0H8vVH
Ye9h88Z906fLzgk4Mydi2mtB1PcdhWc5rmLvlOyB6nDD80Cc6nW6xnA9BU5qvSdpUCMYSSkjMsR6
yDWkm+EkVcl8/NsLdT+vpg9DQkxUnCf/BPFkfsJpTUvrKZ+WY9d2WECKwSRBNV27+6Vf6to+CqVO
QipIXeiqoQ1yKOqCpQlg19X7iFOo15/eISKAD21Jnw8Ttb4de48rgI6hDN25kGXne07P8v0UZbfF
DGyuDAdHvuCN4kjjM0O4yGLUqGRTquKGRhE5LYf/WJ3Ig+f9QpWte1rDC6OpdkkCD0DSs1leJFBl
SGESZeXfm6GXyV5bMS1oKSJOKzXcuIUS+75jGI/NSa01gKaB9QlXWaGYco8gZ6q516+oBfDuSJ9P
T5qgT3TjQsUJeet1shiJNw64eSY+NFCQhpXjkEkKXVdsEqM5fskKLccBry1sryvt4ybUIxhA/YiZ
ei3hCfsMxZdjqogFKyO51fd6bfR6vlWhxMr1RSIUB3hkGVzeTRXnhOj+Ui1IRkUKFCBLy92/R2s7
1uc1kkBFP/+ZyLRCNLoPuJVLpu7rgeIiGdHGRU/FcEQtiJYs87/2BTT+pMMfXwQ5fgJkLfh2k2bU
HwB+xXYgxS5aRnw3Hri9Tl+RCcx4xilekQwhnJXKz6jguDpDniz2Ic7EXby3QNf8HPFHZvg5bnjx
+gySmL4FkQuulOYaF14bWnd1pz2UJYeaIbiuULuCSb903mKAh+Wooh15jVDafnH/YuE2KsQUG0qo
UPEr8YmSPdKPkkxfRuvFd/RYV4iHXWLwHa4+t59JdRhV7uGMhf7tD8/+mTbco4H956Zm8UDezdmi
Wc7OVbMv2CReywzO1gHB24irFJR31eG6tGIQBcm5syQCqNQP9IadCXLWt3LjGxAt8HjFeKbV7FRP
AGeI2oalHGg7fjh+pJVIXXK66tHUC9QWGfokXtFm7c5Z1nA9EyXJ7DslXeUFDz1jM3EwnV9lBG9E
kMiXKijhKpQ0b37b39qIWkXMyTQn9clS8tVD+NEKBggnD6GPxUHDz2Lyfc5/umdXYiLKDl+d8M+z
ouglnoWzoqCBbgTMiVedl8RIEl1XPHVCqVNzLXe4ms9eijjn6A1z2NhZIcD2tlH65MALBpacdpRz
Yoa/sWTvbyY7TgLRwNAOAeCAJiz1jixVQGAw98ZAfVd0PciIqq4AKXdlvOrtbNcJFzJi32KYGL/q
wHUsupEz+fmqoqCIGPunKBiyWI3fEPPlaXnSnnPde7G5YQns3WnzA3PoUtbkYqbKpxLWIoQoQdz2
LF1NBd+SxRR4AIMpxPUNrT9ss7ym8n9EfBji4r8MpiM+yelW6C77Xn6oJnqyY5DvVA5434KPEmh1
6va9+0s1L8MgMf78hTjCjzP+zArTfBgCi5EGEFrIUH2Y3JwGvj5FJU3Ht14FWGcOYNneOWSeTm3U
bjMyjcV8SFa3kVC0kXmhcvnuYIhCyMOM2DwkzLS1D5xyq3nldnxuLE2Jhem6S7sm7xHObyyUHEmH
8DSjfaxeb/8bR/SVtYvgPd/r4WH1fQdXQMMdJawimmzZC4XcJ1Pfu3o3XYzLm+7yi4WnZLMUBvm6
yg08IHl+pXihGMBAvhuLwmf/0fmV6X96olXeNA/Z95G+Eu1sKFw6CDc/ETzeq4vc0pcQsS2qebV0
dHfse3kkBUYTa9ZruGhyE5BD3U+E1MEP6zEnD5WN4ZD2yvFeE36cpYwUgefYy1W7ORxAT97Anaog
1lrrsrSXEAngqBjBs7LXkVAVTSO15kPAYY7JWMRCKOTK7/JZjitRrhzzOyqvFwxJSp0JAt0+hIGK
y+nNUuRuaoCiSjFLXQWUbB2UsuGlAo9pGEnPnOshhsPFrHrsK6N4zqeSEBk1c9KSjZGjhlhQ+DR6
qG3LBd5MzqJGy+Lf447GyGRtACUdyne/2LjBqbKf3oLHYFRn50APF/XbrzSy8Gcd1sWMfKk4hruT
ONxPDFKbODxlpUdwl+Ru7E/bMTPFqialXoqfSWiwnlmcTnpU4f6JJnm90hCCIBRR4SoSDiccMq/8
jqTpt2bIvXGEDQwjcBaaT9dPROVocAonYnM8aV2BWQ3iWRsdqhyLOwdqcZQORS0u4S8MlTRhMlYQ
6WEMLy7kYLBrqQGwpdakDYCE9YfD1U+awE5G6d7EX+dbftBxi1U4zJwzy8UjLMiBUE7KXgzlx1bp
0hHqYBFrgIo1LzA992HHxabEb//adBraeECR4Q4gnnYdsddqofwAOHKSopmyuiZrva8Ya+5Qullx
ij3aca8HpTVN3mg2klqaSWoikVtnlmuojWF/uZ+VcD4rvEZ7GeBpsqnyAifi5cNf4ub+LRmwbCmb
bjOAshCYL7g0XVmA5vr4icvyjW0S3+hfiF86jmI6rZpAC/ExqeH8SUjz75jpgHTYWSv0rzoM3jxD
peHqzvtcr06g1HkwVl3p8FTnwklUX4cQ3w7LRTb/AFYdp3ql6ex2PQ6frldHjsFkkyfqpuJG7KIN
uY6/unToMAPvQ01F2zpX75vVKjz7CZ3tY6bBjmFHUgMAIsYjAc3MAYZvDjPhFxbdtSPi8ZKlw7oK
rxYFibt6ECTq078HYnmfdM+Tfg7qBKKDCkJ/Ibtwt1wOD51RG79DcZ5UcMBiZFhyVWAQBuWncvL8
hr4EC6d62eObrXNfgs/uh/IFwSwtX2weObpaZpwe9JtAZqhWuhZngRV+v9wZtpI1fWEuEIX9ytdz
d2U1FyZpMmsKFUIprUR7fZsNmddQ14C1fy3WKnS7pAjfslQC9Jj1MOXZ42luS6M3vdeh2MC33lqG
0lIA8iM+eFkZCpegiKBSZ7ekyrzPdhFvXif7s+Th/RWtAB9VFOr1d8LgL6oTIjH10B1Gxy5onnO2
uuOMJ1Hwd6zoWFwwJhFyZPH/EpvxOXMSetB19eJbxMgODarqIEsbenmmSaKmGc/OA6WXI0g2qMoj
BPy01vJWJTGyBOx1V1h/ZICz8Cc42uUboYOcKC0HYpFM5wi6KRyshHup0Ug1auL5hBqJZYTgZ6l4
hS28Mw775GfPs9eg86iaA3JNWOcLjYBDfmsUED6agWeONg3dKO8FeZjk+paJBgrSmocNjQsnnkGe
8FiJM38Vhb+NRx3H794YtqSOu7YlwzLBqUDy9y9bOmrjciOy4uTnKWuMnM39jdWtk/FbHlj4OBBl
OI316FAPRHQxzAS4ZW4cdyZMC/10EP4YOF2793e/8qRe4O47ru7idjVc261/6UrneEvk8NySVNiv
5If8CoOrHbohyyvdlmvl4/fN8i5OoM1n2BJ743LGKhPAcSuODe4lLULHSYAGFS3j/zakrZ/7s61d
0G151ZKzDWO7vfzoDVy8rrr1Rfz97XXVUw9axo0qpBQiu18Hhe1AM4bYoSW16A6xdJ8PX5SYcBzt
jjTnd7qK/8crhWzpXIQRwh82eoZoEsQLX9DJdf1pxfc5lvWpt3kDcu473SXJsVT064o3BrU8RuZz
LCM2tL3dyr8tXQnUZWAMQmTPJI3y7Y6ZPf36r0OgnCOlkIIMgofTL6oFbBeRp0I4Jn4Rs1sWmgtl
oHxMBGcTdszhzdpYeh0UNUtwXDqzdlpwkZykJOIiYhEYvrowZWF09qD3h4NDInkeaTc2kanri0Px
4cym5mWagjWzSnskV5Nv6jb02Hw1/GRK4p7m0KH8BuhTsUDXv8nWHjyYkRIDLozTPGvDuNEENAfu
uwVBgvUS9wvA2otxOJeSxIeUiaHiXVCgda3M5E2S3gyz7rDlPaJdP3JeqcKkWfwg5pyVSCVzT7Qs
rF1/6Om7xFRoOqZtMcxkrIq7DBLTuYCgSN38JxBipA073LILkCJ2xuHxttDriMtjd12otzwhStXu
Zd+iJGgSDVyaTr2tw12tcEefqTaUinVNu2xSJ/EXx2sn7huQ5XkaRy1IF1hWtb2fyUbsXM7iiSpS
O8tvp0zFC6lLRAzVW0I1HBmlTkacP8mvqqOsRcyXFdQg5VFxhznf+vjxK/cCzFW2Q8clIJcpWZvN
almXyTAMKDbhLwB8gJSeA6vX6bK087xLomJKZsLmnDZhEcK3DA0LCI/ykPG1B5A3wScRxnHTZtXd
Z5PoJCLMuYvkh7t3qHrVMGUG8GhrRAP+Z1w/tMEibtXf2v5A7DJAbhTtUEHoY3lxQP8bZ0BLRs4n
gyNhIVY7dB5Ym81bkTYnMygAfBo6JqoMKyD0CVgHKZlo7nAQbbggA8Q8O4+8jVeh5K6LYrXyNE/j
Pp2nQunqu+F37OzXr/Qprpy9uWapGFEX0axqVPIs1u0tT9qRG7VgGjk+pMJZo/AccxU3xae2uNiR
dTraiKmofpymuLHOfnb/5xg32bEztLNwaAMhHcEgiS4Mnjp/lCgkMxdL4rEWV51VDuA6lEQ7pC+u
eMxaJBNOkLvh2AzyIimOJCUwwp1Q5aAJu87xJELWr6sjG60src/KZv8H4C9avzpVkInhDQKoOOKv
8EDYXrGZlzr+Xut6qciBGifXVP/ESKzNDdLXvuBoUq+eUzMP7Zo/GxK4GCu697oGBNCWk5AcUxaH
fxgbT4Z26l2rVoYw2P4mytxow56GQ/o+XWH3n0q3NHMDBwDzJ2n0XQCb839hwpLd/5jqNlk7TWlQ
ceYTZTy1fmxVeNPssBDGa4NyLEPSHojX2KRpfTGR4N+CgqqieLC6/6U+89OqQ8u/GsVmdlpda5QM
VZ/mc+ajeIN4Msn4d69b4M3ingyuewbISnCxtcgHXm4PPOiPbvIvmaa1XSRqWABTEWy2EZwKzWEi
+xUsjwpCxCOMw51COZOak+MBLGtb/Xn6x2SjfVkj6pwSghGymue0k2oqb26vvb3UMWF0NTtHtbQl
NDgiqaM8/clqK900Oe14yoLj07sfMtNQVtEzVm0hrE9kZ6KCDh9jkHBt8bYJ0Wf9Ot6kkYPdTSiY
2qDDHptfSC2NrjKOQLFrzhQsHdOk0r9cG3kgOZDuPLYf5SOvori5FgMz67JNFvD6bEmLWR+72//b
HstbnbHF6Wj1MUn5iVVIPFpg1sGtda8SEIxKO+NDVuZHH3BM4soWFiZAX/JbuXD6Ie23hWq9B/M4
fD+oezIkitaDoFHu3R70KvJFBF+r3TKpFWGJ7vfi6Ol1a0KMwbooPyGAfTj46WTmZPKLumgQUwUu
B7c88bs6Qt7sv9CGHlxVLkUcVTuBuEyVitORF4+lMOrD2AMjggwtVMEhCFQ+AJqc99Np2OIroS6L
nccFoC8tfIQKG1dxgjVTOFeNa9letxyjV9p1vJLqI5k//U2niN834EMul474Xq3R1848kZ74qYun
as0EiHXoxolzWtovAn77llBOlB0rR74TnNMpQ/qfOOFUqW43rfz55/lp3UGpuj0Fnn69wrz0pYF7
kywxa9pgNYk/Br8qH+4lmqxGKvJmc2kMxDx23wZG3FCnir6RO/oQF+YnyhF50KyJJTq+FEtEZsC+
Q0uUrDD1hjgK8lcIlRS1PIJVUEnzfh/V5IdSDeCQ+JhDN2SdLsBfIbgimhxeKbkKNZMIeipzGbok
QeasxqQP3fp6ST4E+RXAf2GDeevzNrLYQefovbxkcq0s3YrbCaOfcHY55kZCy1SdaLbxUdzsNZGi
b5mLAbqJIwttHb3Ray+n8iTtJ4XJ50YhwpgUH/vAi7R60wB/bRiAEF+XKM5lPoraSwp69jxE3GLI
Kh45A1Yai2Wec/VP/BMzuqe15hvufhkRO8BGNN6hMZRXZF9nWReV9l42TD3LGAWVlRSHJI/GuSLq
cmXNEl90Rg+D1KATEIsQQCjiXRr3v3UShXqhqqht/HKEI+8PFhkwCv4Km1VLPJX2O3tjlLqJvdZ4
aIw1/gFT8Ntd54rF116nco+3M1wmkQHj9+/laDR0uoliKMJYz//RZhd3LD0eEsdqg/7/NwS0QyR3
YRgqoeUYiZYFGinjDoN5EdKZ9bqfvVhNZxkLYYyl4ScMEQ9+NnzcTLH4Z+XIwFUxHPmYXB8nbjyS
CkAjRTo8USs7Pb/TWaORcYZJbmYXelNmoLdQfQaW6N9QyoVdUw9P6RfZ72oTowN3r9L0VOKPCTlt
PXXM3v2QJi0E/OhPioSy5y+OUWagAkGSGQH4P+JFXNfwyIVyOvnpzvaMK/pfptApZzS0NAPRmABb
lqUUT+7eQLas9xpZI3rgpvytL+Vc08eCe55vJwva98+oeNLXqpbu3vdSRSSVVgkbiQ0T8+oBtySk
fjF0ThTdVrrD6iOnBc8/PHwcVBjqStpvQ36pst4TwwGrD7bTV9ZnSgdvLh3s7uqRH+CyuUW/mFLa
8HV5apSO0jDSlCC6TLOue6nW4sIxL8dttfExAymNt+fYbOx9OIigZjgGshR/ui1obN0dsZrgtWwb
bR8htPWS9F43u4SAmq4G5RDBuA0HUl3WqDrEQzOK9jwTpmVDM7BrLRUescnVt4mGM4NKL9LENISV
Q+7uycOYSSMH6V9iW4iYrOys7pjIT9Ke9z0qMmdGtSTfxilMmQfN03ARFOsG5Oegwn/mOr0luBX5
g9T9SOVZhfQEOMunh0gKVegY72tfx3aJmz+YnLrK9GYvMF4b3oTLAI7QkzeXCPbNUpvYexNfBBz6
vPvdoj5mbaqZPxPtWGkHWWc5vTL44NlGhBtYaVLAVSkyzA4nNSPX04WHwYz55pyZC7Ke62T3tsW5
IhEjCk8pR58ve/h31MFSoPnHAsYj4qV0rjQn2qxsO5qt3Fu+G9dqWKmKaG5NBmrAr6OueP+04gYG
oVHB1j8Zu9B7QdU2rXGjbKqeJflDnxqy9V4rFjTf0LWqQIpHvhKXmfxK1zxwOa+MQyEYGvi8zEm2
n2xjKXs64WDa1xnt0GP6E4snjrZ0VnjvS/4UN75v9cxRwzDgAKXZZ1ivuz6EoWLThDEGZYBJ/u6+
8CWQa7N1dmuZgEuYSbm6uhxBcKgZd6NCVING5fTGzvPGN4vq+GklMOAdg/+zzBien0seRAJ4A6i0
RyMIqdc/b/YK5NuqEcw/LMM/2TLxQZ64ei62UWeuIpruCZj7KHSy/ZOa7wUHeGgYM2fAqwfHRHKx
+GDjhvn54xZKTQ96AusDzv2Q1ZeEy02tnmc7O8WDsAv9YEuSRptfXbkwRepbpxugRDbMCDMdfyCF
w53DY23yaLywryIluducdnWgUVKyulT6TWrxWLUhOrafbMGLsE/R76S6/I+ZybKSGl3CNKrPY3K0
2rhfpsVXhzel2mT2gAc03jv84yApom7HeRCBXND/seVRmMtrlx0NUAz4RhiLwixnNfOe6LnCCuxb
9yjvLRuZE1mbDgX4EzESaSMI8Dpmd6GnfJ6inyXzOWkFPpz2Cl9YA+iIOD5qAJXrDYm7Bv3no52w
dpjERME7+D6ufB777zB0JboPNyXIfN1H1VMyp1AcHuX7mDH8cRYKU56uJ/ojaod2Vvy7vlDdp2q7
2MQm+NUqisR1Vw8edrjRsF5PcNqQLklOIn1lIAl9Q3jlwGjxORAO8TGebvYmkGenrAho0IPusoL1
2vBnKRM5Xkrpfp1a/dg1hpv0t9/1N46jKYWwtKgFXdXxBW/CJvmo9D7y+TMyXKyVO9lo8ytgLIdi
C5SVVMQyeklcVp7GcNwgqbl1JGZI5J8Y+Mwc4ZIPK6Qb1TxltvLBEYwiqBrgykpFqOfpJ+vLjXIv
7UhX7C39beyhyNZwIGlmD4v+k/HF6V6XFWzuoELJ5yuZ2q2JZRXc30VebOq2uLcQBLMljVRhyamL
KpNHTI/3akil3oASV3/RN1LeI2rWNamTkUJJyxx0qIEvYsQqk0U7tTaIBNb/sg/tDMzI2B/a1j4V
/7OLrjKTqcX6aFnp6TIRojlESl7DNl65zQEG7vEg8X7c3uZRIPpdNnRQvtPrc1hgi9ofMcx4AzKS
aLyiD+wIdfj9JRVvnJA1GpsQsV02M4UfWTsDot4R+viyM6Gx0pWsREDDWslANjbq/h3PrvpNIQVy
SpkLJSxHHT6a8mNmGf6vfZDUH7ZWvpsuOc8Un6gGaLHpd3BXr8yJshYw9j9NaDDzScye4t4R/8jp
Q63kTMsXX7Vua25rdA9/vYSa2REOJaUGHfeltZnhpS0OcHrWLhtRQwhRLzm+exf87bZeVGUbHFP7
Bm65R1WeEnyDpRCAUP2YJKbxw/AQh7yI8CN4isU0ifN6kBwUXOGH+TAsBIeu6an+nshiKrArxKfu
15ofWwDaoZPaO8NAP/dQDvKeb5PmXV1YiOxjbrnpr7jTx9MAg/+md/PW7xv1yOr2hgn/7v/qiaw7
MU/BdfqlfU6XyOY63FjkojWch+Vz/Kd0kK9CKW4gwtfSLFIdFMzX7fYTpcJc0MvDiFO3eu11hg0w
ShUh0nUp5oo8hpe3gEA9fJsu3gVYdMUJAcSrL+KtocWe/O39+R1TuS9+OxKFEi1XcjrKbPJh0ygC
gT2rJEBndw2ffCMbfh0CY1mSUQ5YaFemK8z8xYhSfxtws2h0RkzBedMyBTI3tnA8WcOo0l9Y9Tej
C2ZEl4EHK4DlK2fjFy0qHaTrXUqHTlFtg+9vvl3zKMJMq825YEPrJDMgJhizH7Y+evXwe8L3Gob/
usuqE+W6h3+UW4SirUwq841Ajn0Meu1YYvwUKEmkK/C+Lh/u0FXyvbhBPKcrQLif01/eWPbMaLbX
QO2tOuYNsU1N+JllyBgs2PqexRmE9sFBIFZdsnx46o3JcxGa8JL7W+qgMheckAQmA7zxSTF4sXF0
Tv0001dukt1ZCHLwgMDvK+1zPid0FQSwKfKmnG99NmFaPGgr1ErR4Y2FZNmZwq/9lh+gBBC4lXUr
jOReXUQoqkusnX0FFfMRpzzgmsDJkbjymcq7EECie7zDhJooaFUQAO/ny3L6aMHkFuMt+MUN+bPY
rZ7jHaqOPpiVvUA/eyw7F8qNKGanmi4zOW1Is/jkBWYTtt80j4+HZxRLPgK7H52Uu8QGKw0ehubo
rdibgxMTyH/gi01eh9rhYlA0i0Ew/8nQHNjlxetjJtu/+IKwok6KqEYG1CCmlyHFDj18QUvYAKfA
Kgp//WUgVN6BxnPBPdlIayBnFl4F6PBLU9DtYTay4zpd0ZODusfHZt7Jl850w9Imf2ryLx9cg+YM
CJoI9pr/kaoT86E2K+e5zqi/7cXoxoZubzTzY0ehy0Auhct1epbHY8q2Q11U8Q+33FLlTL4N4Rjh
/yBvjmNQ5rhdngJ9zofTdrYqp8z/e2P5sXr+sOmTfJZRoRdXSETGedzzbcKBoABzqoP5sEoyWgPy
DRu3Qmnnl/rGDyGPpEKCy+kKC+gOYJtOOdf7uZIfSP+W6aY6sxDn9mWLajQC3T8dQnbU9hF4wKAC
AY5QsaTUrna+H7B11MF4XNZ4YbF1DhDSKHWCvCRYbQbTd5+yRGNdjzBGj5sTgI38Vak/grr9weoT
nKTISDrl16PycwshHpejYTNWuNpX7fbMz7SWdG+GcGpdR39UsKkGpPYnJxJ5/as/fN+MlFqoAsrx
qN1tdgGAe9cL/xF9Cr9dyVxCHRyxnrsz5CdBKJ/EpgQhNMahPRGZCIK3xxj0sLID/3RkC8ncuujC
ZtO5SAf35sQWHPnC6KLISgVGaO3sWuOoQ+UXLknsM8laMdgYOdQVO2Dr8M66oHqDfd/7FhDa6iG+
7pk3c82s7zgBz/deXH0ahEFa47y6ELHonsKS2Te7fHYMi3ylyAiQLPKeZr5DFZnEfohOCyn5omb4
nhQSBL3KpMnlT83NQPtDaZk0WoyRBLF1XKXSAHJIPJtu9y14TEUh7I9X8grgk3Th//iPbsvYPG8L
H6sMmjynl+sQvbfWEBDAT5JRsMq4jWHNtcI2dkpYtw8hL4Hyhi/vyb7Hm7J4MwCglIxMyolCHJeq
7pLaRl3QGM/b65w6Enfwf3TULKskRlm8i8cJ3tiTMKyNjgm5D3u0r6Gn7Q0fRt8cuhsaklMO/UHO
sDApgM9n6WDrxGvwbIeCZNshhl80uhpxjECtg09LaZ+yKGxd4YrpEyg5H9UZFN87tWRNJJ2ilMCS
rSroR8yOxXXdLj/uhgNMcLgOUPJma9kqbg8J1LjgeCbhIQTgQCsJAnyJsWu2qe54A3Sdj2mTBgQO
FHevqYJxWXOSuO/c33vvPiV66If/SnxjEAkLpoXK33YNz/2HcbLlONfDEINsxQKzESBdGc0wpgY8
EeFfkwuK9oWY82zRvqWaryYslwwp0U4MgR4MTaCAWcs/N9j3T8yPw6Chzk/XbnP5am+GZxyGJA/S
WWEltMsTcyOe8uMlWLW7lyLVeCLA6D25S6uM14A2hL0WdVVWBC1Qb92zcOThdzifj8M9Z2IzOGbO
FsLLBAYV9bI1yfHktSd+wb5SA3bofKS5XOi1/yKoecmbA2uLIQkEP0T+Y2f1OCcg3SfpuZxqWM4L
HPznQgqJ6ZAepAOh21b4Qkx1wDTCsAgDDp7IA1LRX+w1r/OLbPaqunMHY9jzjfp0U8G7lGb1pe/0
/EuVIm76zB7J1thUE3ufSvGjwKY25cB+ckmN8crbY5p700nQx7DeBkIpycc8H1glp7sGCKAnpL++
ctEdJ734W2c1wJ/bwSKXVsyKdDwUcDV8HWGdiwO+WV3uqIuQ7uf8Ug8jIUqDE9LknDqHqE7Wa/oR
n0AOaa+vXtUVp2rpVrMlCqzGe2bWmpotCxy06KYkAStBTA1UeiQ+uleRWixacOIHJWZtkPflwjnE
jv69S/khXKajH9ZgVybGuqqkISslFcjrGZEWxp8f4VOJCPc8T7XfVD31NoODQtALh7twvL4ESlHg
VzgC9rXvXNSKZuVHHzx+xc2fTo3dpYIMGoj02yzcvKwuPXndzFRMcECOtaeV3kQNg7uYpJ/zhXmj
KcgjtZKo2qMCcgdvCto0FvhWr7bzqU9zPIKowVebq9arSoTELFbD7h5NkuDH+FSOn16AGutUmWMl
MMdEe1518XmGcnG6HGqr9mCEcfS3hiybNrLI/GVZf8zKfDPwR4Z03KbqdMvoeNgKop/TCOQ+/olO
N1lv6jZ7nV1riCiF2Sx/hpGU5+80PeE8NoHNPWu/bQP1e79wJBrR89nVUHjDW2kv67vNKyMdaDh9
YVeYRzf6irl0LC+ieEysNROggN18HiN4ljkDH6zWNcMaKx1OnhqnPOm43wprg/xOlIpttka5dB75
MuR7al/zEEB7nmiQIyP86+wGKiQi2NNDGX47zjIxXY5a/g/s8s6I6oOhMMvOVUIcgqzZfeNKQxDh
NA1mZHfzgkAFZj4BvYq7ojQAM/u5hgQDdpiP+B8ShTnB4IAvSLjWlnbEAt34IYsWhWZYXwc/X3Ie
v4+p4hhfVnyR9OOZSKTOz8YLUvVLa5wyP5pAgjephOZ9zsPLynJ1zHkOvDS++bZDfcW3xr+wPnKL
NHr3f4DI7PZdQfBHEZ/RvKRxD8+LtXBlStbXY2KlW0yj9kQTMT2sY2WEkioeXZcOI+a9oG/VPE0L
hPEH7S/kdWKBi7t+iZ5VNlTfInAy9KiVZ8yqeaQINyy/XhSlCCNwE4q20Jy/+eTXhrJv65UYWYUn
xJ6HGKNTf8sdOSe2apI9bY45oenHNzlLNcYSZkRuVJIxhhXICQ8RDIOOntCwiDpPNa50tKJO+1xu
dExzHGqUl+02N4IxqGDN5NWOxhLIu6EfCJRGYdXYI22pxJiyKLpNB8s0v76Inkldg1+4yUPCod9p
dkC1Hw7+crrO5ondLO0lhwPFKQ2AvhsbQ675g7GbEUfUHwshx0D6orFBItUAXEp4FlAsJM7ZWAFi
byDbb/D9zrUbkQrM9Ffj1dsr0YUydUb5nWH6iaNWzGGoVPGs0uYe08E8iujZClk7K0JeDGBMF2/+
HoGVjip8x2iC0Yiq6vczyXLIS0+cAXD5TwncU/FqNJTKuj5q/IxNNVgrHPix7KH2EPscnMeJa9/a
VuH1w8h6syR9ubgP4FREGGeb9wMEldhbCU/VpoLYy5VykHLpfiSJzpdX6hL55Qv5kHzehILAkRB6
ihb/LcyuZ6t0Gr+A3dU4HFUFCLc5mNAJ7b9xG2kszwwArerxLB/vWtB2VE9IfHLNfym5yIKj8iMT
KKEj72VMqI6hSjeGjbhs8akulBC4a+EsznU7HmofU5QeUyVt+lqubvShBBGNMKcs+dHpr8mAfdF1
JMp8yBDEMqqt5yCWS1KB3kSo17rtneSI16oEPoq7xk1ahVSm0E3wsxJh0sGDlGgeyF3XXew5M3TV
dScPxcuevYaJPrXvVOH4FD2/A9Bh1zNhK3CcFl4cPF2CIHHbQ49EsY6oZdHubzzp6+eAPI4VrYjR
O5+aV8h9UonHMBcJRQR+ISTQWR7bN77u6C32mmtawQtrNgVElEj81PsYGX5UMvTjF+wY9/HXoZty
sNnmrkAnLiMGdCbtKMg4C0eUY6yRQ+FEazZ+Dd9cMyANkT+qvWe+zge8elZPe9+3KHKEPJwLdsA6
4STlp4GJYtEdj2uwYjOquHxvXjiDtwR9a/yKhYROwEG9sDMrx3ApavyncybBg7X1zXBYkZmLUiMF
CQkJdrnuHc5jlMJJRtPM+WyerP2wybOe9KTUqp2X+6/hHCUKH959ch1bonJ4/xL9zWnZV+cGU4cE
wppD6AaEKD4RsCApzHuuDrW8yiDQEUUlX7dGVP33yxvKCBvX99JsL8VN51vJDN2EdTuIIQS77yAh
flW+hjL/UKYrmzdMNrxztqQ3i1UpnKwGZV3CueQ1FlIewwUscKnEhtqzWrAusN7VO7noA+o0MjF2
FcN2Uxt48YS7TvxVpNAvitBR1vjLs8OpMQJjZ9MwFJ57jdYIGjb245gSsmCmzgmmI7nurVbqbsYX
VYk8foVTH6qStGbWTjudD/Fy3DCDqrnYeLTjq68F/U7gjlOoppk2eIqiv/hyIDDZX3kB6gITGrw6
9Pjc/1yKTZofEMS3aMZeZsLJ0wKlMG/yX7Imouzw23/VzLTvxvpCZ50ezrLzUkkcen/noI2b3+tp
XHeKxUJzfIBVyguoqek0iyIHJZhrj/s3C+d8SPCXqnC3EMRnV26N0umsw0DXRxHkmv8j2Zrd6iKX
xgNOm+H/QpHkYtt80n57jQsNfodpouFeWYZnX3g2WabmOlRvo7JTW9xVqUPhDeTHEnEjAlnYnQox
kw8GE6tnjkP+LrKkCqHtBjEtO7Kokf1UcjD4yAlPYpZoXZxhcHoY5Jpm77us0p+KYbe6Ppd0yOoz
dAHYuJomgadO+/4HdlIHsAm28L4vnsGGCGTGfkr8NbxwSQz7JfbHKQTLJiK1EzSbFKxe4RNT3g4c
On1XcevmsTYuirwVXb5xwp8ENXhCzhP17WYugmQ8wPQTY1aHhULAuu5F1oeP5zGy/dyU9QwsgHuH
Lb2oAaabR3ImMKOTWixYJgbTp1GUG+nbtGIOLCuinKntF7sb4Fs9Me9kqjWSB0RR1nAZheyAimLQ
YLymo+yhf1CiYJh018mdLYlMj9N1kif8mZkWayqKGUKM3Gh3tx04kwcUu6uzKAiX1uACZ0ImUMPz
ccFXsnk843QJifuPpy31SgHtnff6AQOTz2nT4bdYLgkBYXXc4gzj8g2tb3RQLQUNN1eSnAe2GMT6
MuQekoHbL71JDK3zfPPoPqW7RRGhDZ+rIFSAkfyKERaV9zA+9VkLO3fLMnI8CVYafV6zLG84F82y
YneLDTTakt65JxBJ88Z+t5XZICCO8VKxEr3QiCoLoLkrZOPlo2Cg6VuW+SWa8Id+Rf0EamhDgHF3
aGZG6H+sFm6AQfSKmi20FOG2SJg0MCKEzi7UGLrihpl5JfSJyu5m0d8MLLpP9HL7ZZDX7MHIOMR/
MBvnxFWGndKtKEaouVSdrkbijegL4aAgKnhF1lMZKm5/Lk6LMt/bxQY29cSKwL9r8Aoc04Ef4Nda
B/ap95qghRI3oldJatoqlr7m0ycq81pBiRgBhIcTbcPwnJfBMRdIBHdTGqzShcHJbFmbsgvAxIQd
GBZJc//irNOsnFcOLY5/VNvxdXvTR3W4M5qeXthVpKtS3hgl2mthshsEKAc/f0okmIqpYuFuasml
SVRurUFgVLwayPTPT6laaedZ/iTsQrHcwTJP8bGsaYUj5dQorxekzKtywrtztTdTgoFTXQQ7D/Dj
SQNcq3vbF8pfpVkD37mMaX+UIOTmvfzjHaUwgbqE3cgOi/dObLBYPZxZVchPrAZ96bpLSVE2iwkX
O8Y4CFQ8+XsOfI9GTld3pGpLIeVtDz0OlH3VAiMZSM75g8b9AIErkuUMs1QEAJ1XPYNl6Ky+pma6
1fXTAgtcLfuCTDZbdkQFWd/SQTHAutL1xI4YmSUobhTo6rqiGdFfxJmNxbwIZazEZiDXR8nEbWRT
D82qp/94v+ICtIw3An73YD+T5jYSEWdQa/YN84yBqJGRJW0iAz5mQZNiqmCCaqHMyxMvXGAbTa2D
6uNERrvYvF4uDw+Mk0+Gopx2T3Jxv1YyVUIf3vtpA3+guMifnEaKlb304nJnKwE3QC6Wksg3+8x6
4oZ0AKgveN3o7Dqm2Ou9WujspL/vsL+kEONW+qzWmgQlBbDpHkgHOjASdkvWHSOmHxfJdF+8ljBn
2CiE+S4xAXFVM6kC4msAVe1olOrKu0HV9GITNhVbWhly2vsYe9N7B/w3OPoLlpgbHCTwiXeO7fdv
iFl4XNhdgp1d2Kwy95jxum4sqRNCWnoz0vG4upwHqQ0bF7F1rEQCz7+2no9uv0IddWIGapw1gegy
RRqqIHew8SvqimNR07U/wUH50HjHIB7+heP1R7HKiAz8/sZx/PvLbru0QONyS+ath2lUfdVfA4Oa
84mSM1Ig8nVfeaQ1bKta/UOApSEVrOLCnbEaXvVGpqusUeL3q6xLkEcoYxPbO4bY3Qs8W/bXxUfB
3WSunSOWPKMC8m5V0c/NwyzeNAmU53lFVzj02lTL7dZynmXPkfRd5hJorhNGuajkWN/eTsU+KzU/
gCRGJCivUcR9e05Ho5bixVhejOB2b/W7IHTq85hSYos80e25Ed2fmCQtlJ7T8kBGUbd8L4SwIDLj
VbVxZS4k3uwp7zy4Q6Ee+4wR180FdXKHUbP9CWHMQyy5cDHRjpkKojhqMoEGY+BZPXLJ5JGKMOAr
CtLCPKdI0WJYxV3w3LrZ/XFqO9qUawo7rWLQdEpp5JM9sSDxS0Ue9hzMGFgmlmDp5Rl3RtXgI0m/
luwrLz5DWG/Y04qG+ug1JSZIbSH9X1gP3+C00PUAZG+WU/1DZLBvvtNHYcsR4gVilQUiiAckqIXk
omer1unp38x34IdCW4gndfMJ01lnRWouyoC/rtcif6jWFl/Pn5iTkHmgzwj5MlwH9w7L9MldW985
je3hl64Bc+KQyuZfF1+RJPzOwglOEf5wXukdUsQvjRe3wwNpgTxKOo1eUVp5hB2iJiVqcNKjGvv1
ilPy+KcP7NfY/HcPji3dScqyLzN14Y75v9s1ST7oyxLXtgKcuMVTZf66XR+jd77khhwGn9elA9c/
NNEXnr4/X+VnjdL95F2ehUwcHUWiTyi4RxEu+KBKrKPtUVJUMQc4qkziTQeZH3WLvu+dj5QlMsPy
4xXfnFv18rWpCoAJdzNixNiX+ZGGxjTEPjdq7JfTaaU77A4+q9rwYUlreW4R3MuaQib9wu9toa5y
vQuZ0pCzVakGRNQhiOC7yGb1F69FQIk2KasV5qwnxL14YoPOb1E6/FiDlRF8ISLCZURBHoX5wJeH
gyBA0xsWfcYU7M89YwqqGrG620g2fjO0iBhs0OqidERBTk5oItX/kcr0MTNSPaGEshMrgzAofNVW
37Nx9/3CwleLI+esFCk6GOErbUTS6nuRbNYZEVG87H3z8JDj9LjsMuFit2Lr+HZRI8D0ceOP4Ec5
y4DWcNY/1CEZLFaNo7692bkifacyI/+VMbZDZGXFYKcU6oM3uRvTAXJB6rBKTmWbAuWE1q7IOHkK
aFRJ10qjcqqGKv7AxMFS2O5Cr3iYJ0/zmDrSPdJrbdOwgusc5S7zdr4m3msssRK853bcu8DMjunl
LWmNWCsbChRL23pTr7pYQIWQLY9JmzNYdPSKFaUhgLDnWh757pKtATSME5Y4EfKXHtH8ennmintG
YhoL3kslpao4vLiNETduu5k2RO+U2LFeEe7ww7fRSMMpBOKzzX71Uxfc1sVzwQvxqsR3Np70uH4S
vq7A1X+zUDf+fvBwzLutT2Jb9cVQ9xxoouT/TCrw/lBSVsZ/VpwJDofNcG24zMSl+OSuJ4OLELKr
Z2cCIjz7hQVA2wd4jWDWaZYz6tKU1vZTSMtZHaly8p4bypw4Zlc+ZSPNsdGne6ZZ45zeUTFLKx7l
3rQFTXBkVkpObhCxESueBDCawE0a8y4i2ermyPOs0hSY7MEAnx++hp2smJps/GEZy4LlY57zVMex
fW4tLEvSgF6IYUb2C/S5GSinwk1hVeefKdNrPT1lBi+7ZDjHStHQ+0LiC50mwn182e/cFJvN8SKW
uj9XEtl0FsSM4LpFC2K7+wD4Plo4IPndIiV0aiVGQaZCa7n7PXJIV+aBVJsoUL6lL028G3f61XVK
kzigF4Z8NrwktrxRy++1cBfQa8mi6QxMwmoOLrTvj8NoaW8S363BC0EwWm/mXt6reUySx8oyvZG3
iCS1KqahEr8lFsX4HhbqH+f0VXmZ6TlOzO1vGtB1PBSBhzihMAGnMV938oms0Xfsk8zKK2xf7k7f
IHDOwpk+RUr/PEYGqZ5c8LkNhAqD0LW7eojPdet1rmgLNdrKyANPMNNLDQbRkq96SdRW2uWcWHsy
d1PRAXG90celHNJ77DkL1NMz3/osScYu6BQjS6gQMSD1S1nGDuWF7L1uyH3ZWp9s6pYTwrtMq3Xo
ko5QbpXCxuxS2BvNh7mo512hhwB8BuIyGZaRfKqTe6FrPEo3xFLWNSdIZzvcJMHnMkQ0MjbYnmYN
VEkx4Els2dIxWnAe02bS41+vuaIzQ20zXoCeAW+zRGTrW9pRRcxZlNJJS/vqdDujt32Ya7r0+WwV
6cKlF00PCpbWNhcCffrfVi8rIE8gNjpzNbMlRj9g/bMQljXRqnX/I96mQFHsONGbSMZmw0PTxxSt
P00QfCgnxjPi6sPbMHQsgEGcgm81fc104GlPSG+yelDSjmSEIiGjhQ5092+Y/UVOZpvPy9xMHBwn
Fg3MeaeXHNX79uNUMRP8VdyhZrLzRx/xPnCVtBWaa1bmH+5xmcBHUyazZGQwZEwYERJ4+03MHdap
egOojPMFep7e2+UxiIoihFQpfLju4P4S2v/N0rLPsXPXGuUqvhLRjt2O3XXAa8CZR4HBM9TwghKm
V+3bbFRRbG3CcXCLO8SvKRw3WRVCjUMFc/3YMT+18gmKjmrJE4iZOHFqytbemXQ/UXIRLAbjeulH
EkWmXx/fODDxN8Fmfr886qm5/fI0WPoNVTjsjzTBRHNhl7u+46slG92ZmU7hRtCaDhoedfOv2tmF
7P/HBpc/ACre8B4FbaUlRuX42O/4o2OeJw6FVWK9CSpNvzXVkuBoHLeAx03BdlfDBC0NsU3hRq6Y
xA680SGSs/PO4CiGoFg7dJ/+BknuafkXyV7aFOsghyh1qWg69Bhv+dMESpxUo8U/pY9QwTYbKmT7
UPOLoGGAJ43oGfF0lsirxJZiFczG9zQ3xxqXxIomBTpXx3t1BV9nucM9rTTMF2NxuBuC1oxqO6jY
7iwQUZxgOrHci/zXDx6e7EMzn7Is5+pQeYh+tY+iT1nBhludhFbOak+W88ESNR9Fmz5hVT54hfry
+og/wuU2Gc+k10Cjg8RhTp1xn9mSRwClmJp3vCvYEy3sFQ6DjlSACZe3JmGhuqOW3xLP6rP5jdW/
DD8/9n7tBLZpZ9+L3AHu3C1Eu2uOU70GlnCZv7XiJxdJ612FmZrxONQdMvZUGSYRSzbgQ+kUB+ee
iDZlyjMXbTVaXMsn/6WNykfKTR86SLdGnDfWF3IiJYC6vgjjgJ6ij/fOt5Q7DQtncrmXsxVP8Th0
xGh4+gKi9Za2N7zu31J0J6SbVmtLTucsWRjUXSemN9YIh/Sf2w5M/6Dg3lwky7T+5zzEmATcXrUx
0WTGgAC0SdJPpA+mmi8A2YrPtVrB/2wY9yVfocSrou7SLy2MXeLfngarn6OQCSb5TCQIAxjBYPZJ
j+Mv1d86oujbhJ7gZn7WLF1yv1ycGR9lefekpM2aWM/DiApRAgWWLmC0zRc2a9QsxGO10wwR0kD7
9ZiPv6mrHrSNIFcPq2oYO1M/+dvHT4/qlKXbJ6PQwr/WPoS6F3jxn5in09dqdiqwFGCzfgmvZuzM
Uh+d5c2mP8bicGvcgSt19Tz+Ex8CGh/++mE8mrYQeanhtXJbWtQ3ONOKFBgt3nIO1gRxY7oFd9CB
yriMYqQGhyTCHx0qqgEa09G7iG5H4Q6X/1NGQaOk3FPMAgZ7bYGbIAwmvlkIFnjCCvt7z85Wg8at
zUCQbZKW9UpVA6mWsrmOboYaIEfS9EAsW3jj0ZCWNppcgcMRkQYq5BiIfN4L6NgiPcl9pn7+aj29
yyzYkbjPJiIO3fEuAQ+8X8tHKlJUzF/j6nMHicpcl9iohWJgA99wjr7uJok9azD9mCbpofEUeGw3
L1kTOpxvLy/4AaIhg0FGmU71kLSdaPbCyVY5LSf/35C3br+UnBvaftRHNzvuKyOwRQS2PyVbVC74
OXCm6q+GbpeK3kntza2dHyq5HtLgfql8V8eHaAPhphYoRpK9kP9p+7ybHClPIOGaLuCmeTY3c4Qo
LJHUlYrZBw+sRHxOe1qwnfT5QnpsIEvbvHUMXirihRcamWOpfgAWiU8+n04inGu3FX1EMf7idfIz
bb40TOOC4cg1JTi6FCGkzbr4NbS3gne1ITnA+3yF9gVE9zPUsOOu6iCK85G2gkd1Ct2zYK7AhoRq
AU0fW3zjSAZMpoiuAZiIxMQ3Qp28ReLGsvBY5xQf3ZIHKQAgmD6iLq1fnlLGLRuVxCur+Y7Ck4f7
2dxZ06xhT0f4+uq2Pb2NmuQFI0MZ187xgK6rLKFRkGBCrjkhk9dyu+3TzkDFLAd+riwwW8uINBKp
5MlSzicawGYwsjJpNn8cZ6rd/9Kni+oYp+01m/ETBaCo8iCKMAIzig7+JODVkRtHG23CiFn5kkFL
8gqt80IapJToRe8YvFmr9rf0R56gU8YNbWor3uCHassBbl8JtnMkODohOXueZUKspmBoJg7/6MxG
ajkOr2A9jL7aJPZTla+rG9QKx9lX4zlCYU8gTJpjUfXeHRizQx1Eal00+KpJEWK8wTXbIV3EJIzS
3VCtqNt9iXmcdjwD3B71hmk4efXt1ns8JhUrEKue1W8CP56Jf/qEwPZmcciBbeEQ0sjzY4nXk0Sk
LJDCKLM5mpCFL5ae/sEXYSSWdFsCZNNLP6cnneU1/NAEYSUqYQeMYQXTd8oG5l+Gv+1WBs9Az6ks
ntdW3M6T7zNSOrh+Dvs+vKnPbb9lm7Fpt4NK8ul0PYzSbzHK1343h/T7VMBYDiMLnDid16ynyRlB
3aTyNWlKFFc4yinBwALQ+xc/DpKVjgVxh83PZwRRtgYtMwBs4rmJl9kxWUQ9pAYd95SupgOvmMMS
eQDC8piW1Regd/Eizg7lY6/bO2qAPxpahHCXu7xxe6acSTAy88AV9Z6suGl9viCDkHaNssnlkMn+
uq2MbBXt21TuMzmssJe4cqg61r1w4KgZie+UYn2JAyD6U9O99AX0FRkxtfx4E23glB658yatzwZ2
E/JAgUau1+D1u3KZiHZ/zi07LAnpyRZF6lLgl/g71feGzNSz5RvnRuW3V+UI53InuxJun+PX3Ei/
eEKqthf5rRRJHDhXumLLtrI3b7H7f6yW0pMe3shcF5A37xZm429abcvj59J3j1l4ObxlbeI1sfmp
lmMwobUbl2dfpXnEdDWRxECV2nuZjFmECR3xLYYJmjfGmClY7Rlfi0YgX+md1aoWOByduuYKtVQ0
BUHiIOuDNjuLlwG72UJDPCKjHQmPEDYqXHOF82R61OSVR7ucfoFEA0/PnQWs1jf20APOyGjC2y/8
cLw5aJ8GuwOdFG8X1L2UBqIuzO+jYcv2zcxspr7RriPJ73ZhbJegCAtf6Ru4UTKABQokDfDvefQq
cfr2D25sEtOgzOB+/2wmkD3OhGf5vKN3i53n0jnnDTx6plNhF36a48L6NVYjpOuQ0awIzs95HT37
8dE5qkQgftHDdaC6RGqwRUmgYBld5SLagz5HI7tuvU6K7vq8HcEd60onrArDUAIYhHe3MQKBVdSq
5PS3D2vUnX5PTwSUtlQrO/cqNNMldPaZsBxSLXCtZ1zYckWVYgJaplNKZdEczG0q9H5vvkV4NoUe
m5fVjVJdyPTQRY/ds/Xl7Bp+dyHJvcoV7O7d4nYgy2QV4EgQBWEMXnR9w8vL1sSpGoquEzU2qkQx
oHAuIUofVn+GWseuyz1swWIaOPMd92PtO0HnPmKW47uFzatKSsLboul7ltrOv1rryr2EVQOG3Aqr
5Y/yckvIOg6JeZ0nrRRBjdWrgY16BdsGK08NKladDZK2qinYZg+kZcEB9fibsIq98oRgMhN/6zJS
phN1W5vyguBMbCcxm0dl4Q/vKHfijPWvfEI9DpOZ3pRpHWCZA8XBuT0nc81RRJ88sovV4L71udty
i5Smb9PE1ehLt8biWzeU031QqAIR5EFT0BSn5Xi/LcaltvkB2bVVCA6Go2NYhjO9RrRoAMo8+Ats
eC/+tYoMXIz86Lj7/+e7Nji35R6tRDR5s8jhZ0akkTBkn9edKRQlkWcqcZGMfSt/QGx3cDXbFnVb
Z0CoDc9e0Xp3KAcM10UOuQULp7rAA7BxIIJFx97E8t0zL2mJIneKyNQaskoSE/55Kjjie5v1WMwE
0W4VdvnICdSdXPL0uWmY50Kjb5Ps1WKcE0YoagbZi+strkkiXYsJZI8m/+rCkD4y8aH52/UnHDlv
Li7EDucpo6kpveq8PaS9v7oVzNpsznf9dbj11cVPJHyHyIxBVjI0kFNcx96XFlsmw1EXu2tEqW6b
VUIPFvHVfENjgVYirgwYr4fbfF6NlsL5M+X/Q2o+7nCAfWqIFOJ3ZfbVGhWp230YWPAkG5M45IJF
wwAS7SfM8Tpzuc4jIuYxuTiO8UVZbf++8Uah1mAl2bndwXtNnTUlmuN7nIx9nu6bM7nJ9GBe1M0w
y1B2MFE3arRVwFi4QqFurKzQlv0Blchrrn6Qfv8EVypxE97sO3UxRBXdHRgYuGKFE7HzLa8aMo5e
2pq3WSr5ei6iuHdD0P2lKE18w7ZmkhjonlV8JgP8u9jdu8ta0a088tcfTPsLphc+l+nsFLEuQuB3
Q3VrPpmr2xgvYH/ujYgoaEV7hz6B7DQLn69Dtq9WCrgtP3PBiKsvZKilx8CXQlZasxJPG6RS7t8Z
kFj15Pzix/XKOsNIRPvFKNOCX0Htlmd/L0xRUP9rddXDXtRfJPwtHojZnaI+ylm0b/iFoH+7N0oi
MRf2n96S7ROKYrCKQjwHlQnsvQAYZqw1iZtzMxDO0HJiPEYfkFB3WOhMDinC3NVjb7KIOgDSC4vj
UWIet8MyJC0ZNn3WG3lMRbeF9gP7EJS5o92cx23/2XVpU42svctRDKiJBx5YwZRnv6wIaNS6ttub
b7ErrDCUvM/vUtbgqhl++/1y5Wku6ebg1BFluevoLSjGr66RVZIJY2+r2mHkmNUTkb1WHQWj7RB/
Z7siPLdqiXvRBtvo1e5Vo/bEmoemy0ndb20xo5vRhNtt86OkTflgMscgIPOZSJuj93ppJLxzbRw9
l62XriePzsda9CMND5+g5tV9Li07AxFoi6tRkDNTbPfmGR+m3OBmwdHMZ/f0vu+b/fDbNMVXMRyo
LjvszehVrOfjOews4bpcAI5kCIOGeitAdBtQJEKUQzgibSp4HJfvHPAQZLOm84fYa/8on+uFRtxJ
aDLGPED0vMgF80MQNI+thbAGStHxdh/Z+qVza/OgHYr8YjtYkwk/iBWWsoQKCFz5itI1QerLEMus
2lL18R83KuS+ufQDgjENcSaGsg1BnO6VJcVen/R3iSMF30tZXsfaiULnEdWOcUcIVmlUeEbwlDuk
qgT6Sg2ng3f5Qb9C9/6brfcOJHSsoa7U363QDdIckV84SRFFKjtG2gKgItqp+A7++mnk1SB1CF7Z
EW9oAj3QEAksQYX2l7OAJQYKLD7Gwdbj7Mohsi1kaCMb6vuYUoI7u3YtvFNa0eiqe5YeEZc+7glL
/TMEZhldYIY48Lwh9DfICR442OkU3POSLGqrYg045hcZUiqk7Hv5wqhzMpKIb19PJat87D9KtAxD
wz0NrVd9N5pgZYKoasGbQkFBMx23UUM8jKrS5xqCpgydEoVtNbaD5Voeg64y9n041clhfjlBWo1F
3fDpy1oKA56FtFIQ+t2cYf6FtCqaJwnEdgJAs3ZKRB/UhqLST/arIzArwaErbkk7kX4jj7gxwNT2
qrBrTkEvTq6oITwPl56Sn7Ri/pgYRRnaU2tsprMWQBxiTxYlTw4wKtkOKOptW6GYdVqPPbaOIuOy
+MNaV0kXsm5JCMyf1o6VvhdoIHWIyBDhSDIwPKXtS5hM/dP1gAOU5WlH0ZdXEJqRw0JOSPhkuT+v
Ce3nR77AW3aEAqTg8jMGKo59HdGhdZkVTGulcd+Jt/Fj2HeGv3WoJJzE7tG5w/fxTf+nYhrrUs0+
32vELNe0RWRBYARoCM5ixDZtwgTFjr/sG0vGILWtREKuEh3MEX3PAlQAYrfCULyVApuwx7jBnkhB
r+pKL0E9q2EYA80Wqq/HprYx1KiCnKNjQU4A3iPeBJFkexojkA0ZttIVCD94JX+6LjEKZNSDNtVX
uk5IEVyV/dM0Xn8ZC3Aj3Jeik1wLdq2puBlI98rJUGlIci9uCmVWtE1GSSRwUgfrtxaG+EyoliJt
js5DNT7NxYP5qe1leY79zD/9VZDO2p8+txo68FMZAYXL1BWZzFICZPdjdoA8hRwGYnOE9lC/sawz
SWP/Gw+WHOZeVm9xUK3LHj0sI6fLaFNtOPBk/3OcBGVrKIvYnOdtYuJFmJPyBf4/UesUkxpNQ1fJ
vpHF5n8RLwAw6lqcRnl2pUfZ0e5pJxMNyLSrwmObRuw727hbsJQ+eBguPzVN+lhqPCWDX/kIk3Zg
9ocZZNVqbAVUY1rXv3umCKHQrNfXX+o++t9S2iWqjIScZysHjKGZix5lWgmnW2f4hdp2/7sZJlRo
VuQxCyW+GyBm0yc59idUAfO1jRwNyrj5aZcfB+wY1vgMpiFAWhyUiotnOksRD77ggNuhJ1pofM7T
Z/dawtJGuBijzkVPPfWTa9vlU851g9+7Caehz2cKmMSdWHdvaQSWbF2k09ULI28Z6Yako92tPvdn
l/3XqAh5TQ2dZp0bfnenExeyXhVdM06zW+EnNw3uXIHWaphPwpMkZ1SZHsNJuEliQ2d0KSGA0AqD
jWDZtX5Cgpjg/16eZ53feKNi4fS5m6eff2WF3cOaVNJm7PskrkSZkH4Tdmg8d+PEjEO81hOl9m5e
LYiA+77XQ501QCwrEu75/SAmX/VN/nPb7ytPvwOQc/r0b3NbmXK0ir1th7Uc6u8+KnqBTJLlG3I8
ZvgIu4THBBMcSodR7JDT9BarStnHMbiNCnHRYhyqBs6uhaueIgo8zev9o+xhg0zhUUbWzur58wgM
oE2wj+gXk9YDlWCbF/JpRozWR8ullb0jHLPP88GcHCpAgLFZvyPwp02cpoQQlMPjIUWMosklV0be
mWkadmCuCeEMqYXsovc2SfrXyrjoTrYwGEVGI9TS8wv2RzDF+4dxlvr1jboDDAujk3lAcCMqujC9
tRri2m89PH/GczDnc1S93fTEPttkpTODcq//nQyCNSQUSXZ43t+DoP2FDg1xG/N6hz/hvqzvqGnJ
79AG8kyOgHd+qrT83p4r78O/R8x7CSDP6oskAJxzirgLVJdsym2LhTA1nt+GW7SlSHS6zhrMLLRd
IriK9IJnLHU+NrCThI+o7D+xThWP0+0u/gp5aaDRl8YgCCP0cv+uNkCOc/jQTNLjzj5hnlurwo51
aOmSKBHIehFIqX+C649BicjJRybipSNvR/eAuPev9txtn4UqyWCGuVRQq5465CDN4np/ukT5LYsz
saaPH5gPcA+7eCrRFYMoKoB204mUsA7Lfl3JllEDNqmKrXqwybsGKo0iG1m07YANgzGPhiyQvpfN
4LvkNM6gJDGIlwDIQc53LPFR3Fl2F4lCueWJUJRj1tE1ybSV48Ti2R7IqgP9FmjU1NCi1didOZB7
iPfZbRdOirYlYjudoZjxOz22cFCykqFDCih2bfvPV9vg0oAGyDb2Z/lRdysB7z3gzYfc2Sp389Lb
WPxOhfFqzgOUc/cV9x08S6qbVpQsUcTI0fpTvSFoyXw7E1WiDRabNyNFuSQA1f439U+9mtuCPSRp
jpvuKjil9R4zOWy0N6cndyWxpMNMrx2Mlp+y1lzs9br15DX285hhUf3fF3bmBqT2bqBgx81fVQQP
Z1zcfpV+wbRZUY7HjZM13RptYELZOFR1rCkf63/U0Jk/WhcF/2YoKRCxNKon2sD3wSltgVsDHdHw
1DFI25wAUzHMJzxkx7uYD7L2HC/gsyz1iAYWzh5SNIA5cPla72M4YtfSAL29wlymYRTXo8PJwUwL
GD12oMlwEZm4vf42ZqxuaCIFrWBbzLRMBrpWszUgct88IF5qPEwa5gPiWLV1Arrzhv/dqsump9Qs
o+E8/ZfoJ/8q7r1rumWdm9bznKNgdSukK685NX0Wdeuwz5JNZZ+DMYs/SJncad+AuBssoRj3StNb
uq5cDSaf39kXr0hVaclxEtl+wkKAQsdxS6yJiXYlaugyR5dfSMujyX/M7Q7qYTMKBl3cYpxUQvyw
UB1SnVV2dvTC1eUPHZOtz7Jb2zQiemtXhzIANXwOJQ07wWJ+/u8AMGB23eXGbPneezk2bvZbvuG0
5G5v48WfWqC+oAeNBY/PfVl39YpKYIFjq+naxJI+CBhTKFxUwOGIbt3bE8w9hdLVorkK+HoQS+L/
vZo/sil6+gVhpJ0uRfD3GMdwxCGxtsn/a3kxn8iPeDWPGkbryqMQT/LZ0apxi8VM2r06m7eC+LZ0
i090MsDroWsOwA2EhwgkDi/snZEeZvGmKs0/BF9HMi/oCBXN1YpfMbBtDQsJHQ0HgShFsULSOhtO
W9E/4mhNQYHxtKPpK7LyhR4Wk2tCL6d/heIIPjg1RExoaIvawjTCXqF/t0qIDYcV438CEUuGaP1x
Ig7uKFnUtL1Qe9QyIOpqVWfW7cJyJW/qMjI8y+MKmyPIfbQ9cawAGLcfFJsoAbWJYtMKdU2RXqKP
xEOZT5uEOd4eeF6BMhNOCS8l2yqSQ8ra/ppEcBgXNOh37nBt9AzOxYr9rhdpQcGb/Q4qB5CUUJFi
Hf2c+bWikMWV0JsTJyGYu4IOvoXxWwQGdZ4xEOY8S/cZxdhvdYR0ZFfKActQdx37Z0IR99u/Ohgi
R3o8sKndVMlftAOfsu71oX/Jz/Lcl1hL7cMcLUKKjiRkE+vAUhPQkWLVUkyStIgIL5c1Rr50TOxU
gHcQTyNm9LuQuQ3U/LY/9SYALQVi83obgkdRRfamBLBNDvhtomN+8vgJJnV1vCPgNO/e0qRf23w+
JSsHo0xxlrkP9MG3fQwN3lbCwEuiJKcnrSMvQMk10az4VefCHTApJu3OdsYQNW7HeA134wCzIyUV
ENBJ7plFQOj8UhIooFNAojdnchmnkoeZYRQNqxpriFAK9mgw78blPW1GZBvqnasytz2HJtqXzOkZ
gpVtFKuK8HaiHqnA68AUShfJVEOT53VgfaR2Vuk8KJi7oe4B/EXY5MtLCaYEddH1T15YmrNTQKiA
57uTCAWAl6dhiGiHUsnXCEI3q3i2kxQU3AsDbYoHBNAmtHHF5Clg5YyDCm6bH80/BVe8NIVgyXo1
t/Y1/5QXyDKsgRdO+HhihD6KVBkb4OLr4XUgd48TNHHz1bR/Alm/rKrSOaj9rxZl1eCjj8VogGe/
hL2FZfw4xbm2bGugt1irNCELLInoSDrtpR5IYj6jfWonOQyI56dgA9fglbErvZ3pONRUWYsgWcy8
oIiRnt47w60nzq3fYD22kDOHsKRdy9w8WIG24QMBqRg+Eka2iHmT4M33cJkkn2u7auRTDYKEKFqQ
wdpuHCyRX5DOcVm1YKXlJltoe7tFxVFkbIupX4BKUc2vWCaTbbWON+VHSjpIeX55r2+2JxZqjYk2
5BxJn49xYysYDbyJiCDLMYHYWQpS3aF+eaqKXNdTRiXCsP1J0BgMcZJZFGOlpmXxLMhyhjltUXnR
Lxu0KGq8D8b/+rFj2QP8dQf+jzeEbfXqeanAeVVbpIblJbdawr/8fYlt5jHfhgeXt9/AMTjqYPan
JcWb9nHKVONeU/YiGLvmGRBuaTASYKFCrOJfkRVDLNjmDmBtxFTg81gfrD7KBa/h+IOxywcfii/k
+Oe+AuWVuUCHmKLNfUoiJLt4Qa2D9vrXgVTJ7kf7k7YacCNvPhD4SUs4r9Z18Orm9xJuy5WHzCt7
XoyS2zt1O+SMgElygkmHcLJammA4FysfopFpt7cfqG0p60eM7dLLXMKMk4bQJZzzwGs3up3m6Ci3
gdXVvfFWyn3q171zjnhzTgZhGhRZpCpoiyk0hZ0kb3cVX60ZMQAGqK5AlorQ8HyCxKWf2fUlyY/R
CGSp7HjWfeo/gGo2QdCUpM7JkuH4ffYN+1UjmJKu92HYgZvRFrzNrEXi9oDMiljiLDyedhNBDFSx
yJWbnjf+xnXXZ/tZx8FWuwIDhtBFMAEO3N6YIuDm0wKubedId0ggQEPD30CcrPX57recKL3R8a7O
ZY4lDOpREzKja7yL+ne217/Mi2x/G2k8J1liPalt8D8NVI4bPQyx/zp6Fa9IrUzYkxseQw/Meal0
eXOrOE1Upf26cZGUkxDvH7Smv/rVnApecR3SutsQaEgxJGr08CQLxG8tHh56nhNMi/AFfMbGa8i8
J4SFPEAEA/m8QBNi7Sh5KOWBshARW2fuSnKbHhd8q0XJIe6cEsnuC1KRf/x9hPvLDMkdL9aWUdTO
CocZJwFkplIr+Q7055Xqrzrn/Ps0jxXbybfMMDcR3DV+SrV8qs1EY65Q82J/hj5/zRR02Lof2gAU
lk+otFQOAncu6byri0Sdu+KOvQs9Gego5+tVmQOqvr/WVFf/sTxHHuiYTyB4wLMnTlzNOg+/1W7z
oir2UBOljHAXZV9AmjZ46+MB8e1tLmxZv+IprOSc7NForJc1iTiKZOEnBqU9rqyix87V8Gj3hIt/
7nxwraQQc7liMEeF/py8iomPXDtQ2S+gqTLBOnTUg4AdLVUoDa7llvB1gpPuFs+x9hBtnUIlym8w
QWeIng3fZTPFO2RLXb9bHJm4tzIoveUfhf48fVaNSXBR2tyjkpQTOiasiF1bLiKeHE0+jHj6npWr
tMEdI+dbr7wJlUkyWK/6wG57fnT8F6m+XfLGGKehr6MeFGa9KvroumqoSsjESi5SF7wUWIRw02+x
UrzRAxTJEhEVE6bgDM+mVDI24WLt2cpnijeGbsrJfj5517t5oS0g8j6LkFpUKrrng1C1olqlQX+t
m+a4MqOFLDou2twkafuBjyg37hFPnNGMDiw2dILfk54TyeBZErr4jlcbuhAt9A6AUg6mjWEBiCsu
kCAs+gsptDMAqOJHhlsA26MQd/QYPuXC0xafBBWIDip6K5gZXZb8ydm+lCnpFrPFJQKOXDOjHkO8
SZv3tSsTO4IoWZQOxqfUcbXRi1wuiA65h5A+8+12EKKCFJhUmRSrDU4GHUCt9jw2s4+lu6xEVfJi
I85upGiNaguG/UmfV7Y8Y8miVsodCKDOZeXZ3loQL82mwXShqRUczZxn6ClV2lwyTUKc5z2c/A//
ZKyf00h2sMmrxjiDN/MA+Fv10p6gofQPobnEqVwBDhE5kizPvb6vxfrN5Z1yYnB3+gfuLOlpGSNE
Xz8GCfA4KT4lH+B2Q048FNQDWcQbrETPG/Ess4AY3K0d/7Dg8kJiHhwd+xs4fvaQNIuyuLVw9hRN
2shBi3XhNROaqgkvinQOkzbB67Cjk4Wk0N9iNJJJ3ORKBcjeJqBZk8BGZT7S8uTGx5U2niaea5pV
MNcUNR4VM2OR3oWTE93eB+/X0uXZB8aPp0GGVXQBXIwosvQCZL7ISS4LT610ignITahfbm/emNpU
cuofu2LK6sNr9J6+zvX40/vpBSXqeHXH+eiwuSZwjgSGFuO1EnHHFKmA8opd5cqIi1530yPapBgl
xXk/pRM5PYbCqvkzow4ao5npl1sI1HngsNN+nRmSPArs3D4FA0zrOQdU2RyuaU7ONYn7u93U+o6n
Rx+1qMkexU79WuUQOc0SPvgRUXHglaPb9UGka+z/74ESXP/9kYHWMYnqciN5tgYpU/yzPxjzHPZe
jnzAY7JfkerDzQUyb/T3jZBpFeXQqaiJQOSrwVWbnOoCEx47ZZGv09M2W8QaxbvhY21VBXcAbRsg
CRXQBX6NOflHSu5dH75EzmnIPJUN48uh3KCa9HNiCh8XDHsst4MMMhrhfZy5TBN3qT9QzKiENlbx
z/MnIuZd9k5I5rmJGHtcu6PoZreJicuos6QuIVim5xShWuvAv/yQuPgL/P5VqlPSIOiU5rkIgr8W
mwci724dhSy1RKTLKufK64RakpAVMXgSFGNrOYlNUM3fCvvkGwWvsvcLFKDN/EDxGJzSrB08oZOb
GiHanG0vvf+CxqLIdf62ebYmxprPAAAyOIvKvfmRwE2GU3ymi/HtfDCcNnWi1hfW/rBkuRurEYU1
4e1HL2hfk8J0z7XANHsSJOi61m5Xhholio44ktbg9Wg6oTT7Vk5GcdYGpuIDXzoNQLfIxpQgUXUO
fhmr3sLvqW//3FilTWIWUtPVEsYplA81z3mJc/KhgATaIRo6KFijeYeuh50HHqTMp6aZ4no2+TdB
DuONc8oyXwSPYd23BVk2InHT+56RwEPdQGZWA4ANUVZrRE4zbZ0TJi29YAIK5TS5GnLqKADByrHJ
D5X5NBDi0/i7ZLJi3ikUUvrehuiHj3e4KH4A0NrH56HNms19tlNssP1vlnZWfuTbXTiJ2pCutKZr
bigLPWTODSXSvIKjXS+oMzwewv5aGtaD/DTjErL3X8lFkRiLpQdpWYyEu/q+IvKaJGqizJms664s
az+Zy55f0HpuxkyR1jeFWeHv5vORFJs/vlHw/3ACQphcXU04TfVPbIbitkU3w/9UKG+YOp+M40QJ
4F3LrdLIhMgxcxEFpvhYd8Z1K3oyLs8h7KcoIDltu3BiWLfOU4HLpcfUWMyO/IMlloFnxKXXaeMa
01BING9RL3vG9oAbMArxYX4tEZjxHqBGNArgwNDy5Bi5uPsblYdJM6F9XrARWbQJ22BEQneUuPfy
5QeXqj4JRDMOAjYSWQCdi/lvwS/IOZGbKiyIDF8Ce4ZToZXXD7qSMYR9GgCymdTac/+tR6V5LqTm
cP/vJKW9tuhxi6aoZGQKhQEOrW+MjX3WnJNL2CqutH+PZpTmrLglK1sawfbVd83LyRwZH1yNN/ic
TgNxbfulQ/j9ye5GN+Uu0AxD1RNItihpmYqUwzMVUtdtmBjpKto8lyx1uWBuvda5q+GKrWGyy07p
1EZfG0bF5BMc1dOWEUAkLK4ozSj0cphezOgX1ADoP1ufTvzV7CO/EMCCP0paT+ayvhR5cZlFwvdC
Uu27EUWzRY4GaExgR1rKwAL+qR/LH/T3fqQ9nEczW6y8+eWSXCXrWzaycEH07IduFgN8zDiSZlZ+
1/fZYaSgsOqULeCgXQIVW7SzIlPfANTHqD3Kz31djDJ5O6P2S8tCLKF8tkO8A97Z/BzzJtYfLY7j
5s5WRxHFsXMfJY1UVES7D6ILXUakqRNQdRZ0MzV7n3TirLuM+ZczKwspNw6FcFMtxmAJwgi/2ArV
On8U0+GbExVaKjdN7k0yjwR6izoKJIgtlFYmjY4jOPOFtYqc0gOHsp9qVSjO04oWP12XHg/ttu0c
/Jsz7mmceUvcB0n155n0rOCMqZqzQuHArDMSL0tEVDDqpo4jTEM8wd9sRbwKshQ9JhIjnYpRKb/C
9QikIBTj52+LFzcKq0dnfnOavHAZsONfXjYxaJSXQ/NddjbJa4sZwnKQ9FvMMp1TpKB7XLwIGGwx
Tun8etRjVQQW4UlxZhmkED6eNyz3l1XILHummTROHWpz7Gsn1OJ0475msFtbMJddcyIWQsRgoKAl
HoA8eW1QBDxIQ42z4JwhzI1h5LJIgjSEa2ixMcr51h6Ppe4fX/vLgiyOyS4L/cY+DzBVdQ6QPKoU
wza3vtZt98UGPFzAr3tjM6Qg5xI108wcYe/69ool5vOwUwEoYmvBMqmRRrb8k2i24LllR0BA/wK9
EtAM84A3/77EghboSrM1LqcbSW44fvKb0fCbcuPknwIzlbBV/sWjEvJYToafya/h3Ch94ZoncGjl
g+vk+/gZSpQ6gIhUsZz8Uv/76S+cXxZebjk4rlsuWjy5w93qOStI6gBXTx0Bvn3hdw/F8QCNxOST
XMyavk/naDH4Kqj3TL2q3UFhp28PH15XGyy7blIdh85Ragpgh8kH9YdpWGPbjcht7O62eQjMcul6
V0ht1/gTOJRRBSGyAxu75+4xZTi/C3Bs/7amuoWcOFz0gBhMyX3+2pBlYEBLCwTvrvlkaxAToNXQ
Ux3ySiQP3zHI2zmNejGCKN6U2TZy9R1isFMZUxJeB5Wl4ra6g0uxe9jeT4aOQLAR21LURD+zzK3G
ozYuJkTiwSP0LF4B7/3TbeD7I/pHBdreHf7OlRa4vh1i7tRig/FUXovvCMayPJMbduhPdoONr80I
PtEMd3qo6H1RYy7d+4bdCz8EVnu8u1lZ3+xozFblRuVF+X8x8/KgqS7i32G0krSK8NCWPIkjnvFB
snBf1YTeGEfYjGI0suxcri0obKhdOI6r3T+Vtoi++jttH050Et1+SluJPUfctdRkMUfN0yUlITfT
59ukeMYnjta+br48NTWixFnhWrkcuJYn9owxpn4q0vGV16aLP7V8jvmKQUB0T9fnSMzYjyzLxoUY
7SXBqlOYsNi2eoK7JhdnV0hmRMGETWUM4wa5IxclnAS/Lq+slsam0r8W4G55WsGMTbD/V0vS+jUR
M34MGimsitNuuR8jPDQAbc5t/dhVOHRYkyK0UnlbVMg4t0vHPAmlKJbw2bBaV+jee5dx8La970fj
bqkZcq++CtnAHvA7fT9IM3dZ1wV+ADkSF43MaOVLzD9jh5FfNLEXXeEHiJB3JFy9s6TATLFruAYc
ShhsohX/a1cpXlLxy2aA7qr6lUvuW0Dc1BVTWIwPRWUaMMZGg9bHLYQs1tPN+J9jqXKNiZQCd0XB
mkz6o5cikYtdxbckQfN4v4JBAzF3833ifddIeywTps179mst6GV8L3Z+e//rahGBbePCqoIT5crW
/N3D5yOeHTB7mVowzX3JNx1ZWqVqR+pe42tPqCqQBDsqalLZApniQPkl87vCGYnSv2apVA6iLe4a
YSwFq3IvxDQ+Pf+lXqdVg9jRPiYLbXkZdklDz6ca8RO6nP1z+CmTVaU3LhAsNonQtBfAmOBZVTii
JyeMxhSjB2F1Ch3NFkaqHMCvo6RZCyV49srJhn9RpJtR9EOmsPrnFSSf3EnuBe4n6svCRkd5IjV+
GX9HCqQIYsRh2+9FPTS6SioQG+IezeNYThoGoI0D+JkG7HLm/X3yKeTo+Gz+ZrLFTNMc8Pa9B5SB
1i9/LVd9WQKcpPStvZWv7otMUGADHnpLATM5Wf6h+6VLbpdX1oydj2Kk+034/idqwnWh1G3Za2KQ
HuCUblmsxJblXwWqDI3T6Lm8pil264RSArfsiI2ESGOM1SzHVoQwUKk+xS1N7i5Q2YXWarVGloXF
dJkb/Qtc8MkiNHHdarRhH/xDnjaEixJ063stETUcu1wf0ujiYLTgu7bIVVyxJvvkCOLeuM6o/2UT
v69dY2187zCy2Di4I9ysiXsk0KiKDMc/A/LkVe1jYQDwounq0fNC+DPUBAsuBZcyQtlYBq/x6lJw
jNc4H8XRiml+IJRLQK8bVS11vrOJaQGbH/vsVVfqYtIVlSf9EAiF3Hx/F9RVbVzgibNfRMGPVI6H
PQQKczmmIEPzP/JJWh8OnYPsX37mwVUWXl03+2wADww3vusrkxSNHtiyTgXOYqYfAwHEmTrGHA/O
X7yvVwnLdgYnpyLaIlQwqa82dZLuUbvV1hKOOmxcd8etsCUKzc8lVnKH6Pg+EuG9uGFFTyFtxuAF
bYZTWK/CKQzW7l80XocT/pP8HpY5M/wcboWoBHa6t36QXcoG3YNmy6TzcNjqjDPzHcv9Nr+CdtZI
EBdOYoxJILl2E2FlF6IBtxl6mqx2g7GcEGpLRfCEK2/9ej7L3alGA9F7CJV3ITZDk0XwIOWqi0hX
WgtKjiRULqqRtFxEOV31JqBt/yPXOHq/hvMoS7Keg/NhuF9K2F3wZ+621g+8y4M/ZXwiWzZEqGVA
VsiLIWDSW7JBWCkWgVdOPjKyjvP7agbw1aT5C+h8dcDG22966ceWZKKnP7l4ZOOh7EZgo+nuZBFh
sdn2HC0kzLzHI7zFbnj8qjZ0oIIHTrHxzLTMqWXQ6ixZXyxu1kSwhmijEH5TBHJ8iIlWBM+nXoG6
T/d53xz9tKZihjm5OQ7gZjSZwX9JFrQlbK6EbMyqdEicnf4e366biUFbp8BsTJFD1e15Z8Plkl8/
siRTp8JsA9v2J6St9/x8aOFnARvCG5mdKOGfEo8gYqMRL4vQbVlEGQChS5PLxN1HH5jBxMtNz1Kp
9FPI2noJT4M+iHqBO7i4sDBtiCuKAM49rHdaeMmfdu+Z+607uI9aZKPWYC5RWu+KdmXJpFLVIKN6
P1yu3vThfkbndcO7Z0mrHriL0YgKGQm6Xw/z72ZiHR40foAYD+Jwlc63jSu+E8KDEuPDdQxSibBl
uTLQj9i2PGDbelPQixz0+RYcnZuyHNHnYHkaCNRYfEYI3JflHRuwCZieP4+3Pt/D7uwA4MoCt2Xg
KOLA+JzcKv03eOUmvwQ43NGEsD8785mLKTcLyc+WsHxgSVLxnLxucHFnC9Zz/Ar9630Rta9VA6xX
59e5RD5zC4ULeqp1uSVlGC9Z+bN1MWCmxhy5361EJLItrMegtd7yq5iBR5fDMxVPFfRv43iSBCMA
20R2YvKtvLEkWvsUFIXMR1zcSsZAtN0e90Yec+D8CKOJjzaYCbofe/DCuQPgSbhXDK+UOBuZ+sE9
tiPbTm6eGXvsIOcnWOGc3bJfzId22JejxSrn3Br8mObqwOZkELz0X1F43+XaAJgZyc3hoCjXzOYQ
yhg97mkdAn03BGx8xT/U1gkqZKd04IY34pCMcLpHbiIprkJVZ32cLNXbudtPMtnzjnZMi0H70sem
IbsZCM8Du2EL11iMSQZe5bppbAJZxLZfxFqp82ME7c15xhpoIczj7xgQ5NnuJskg8yxmzdTV6sHx
/nSHltZFagawuwL2Krev8dJ1l+UL785YHakq6LxnKdIyA+72bA7VHVhdHBT9BboxslYXH5NI34Wm
3hr10LJZQdQKY3j5oeXRrBP5DTLZLxDYa2sgQwnRhNFu3QIdbf+WnqkWHIHHkz3pT3pKDpBU97bj
zYfB3YBU5n9p/DYZ2bCXi5UBauqr+dm1gWLd8n8cQRD31/dq46kYkx+xV9GsisVWRtP+Au44CiVX
GUe26jMtYLIbUQe37V+zKm0TGerX02zu1av/kJozwyEfNduAGdk4IEWrSog8p4C6RPAeTgp+1ZSp
xjZGoeTlwTkqa54O5ogse/GL45Eu8ir7V7cr11QAd0Ey4XJcU59gb7SIqGWF84zYEfs4X+exlHWx
+WIb4TAy8O4WLwQwHhga49ywUOryZKEI+UpDHg/oPILzbnrME+o84zdDFdsIbX2Pd0JtBamnpWBM
Lkj2nUVyxOt84ULIL14gci88yvooAPYAhUPbPe3gAPRhtYcyaCZKu9VVE+JccUzehWVz3WcBFRDK
p+atnAQdUMT2dEGlXokHqh+4a80uUk/2OHk+31+SfXGD4UjQ43rgV7Xqsp98i44MSb++FGkcSQGa
q1OMCmlJDG0ZyJrvTP4kjau1As48Ix799XR6zyfkt1LRqXxfhSQI5UFL3yF9ShvBFXGUku2Gw4tD
iyZr7C0UYQwIAsSXxc04bBaBNAc9rPXgJcip15bC2vXfh9BC/2ydZbcLSspzJSVaXFQsJ1C4bWSu
nxqA2noAeSIu29DqPoMWEf5n5arVnd2uWppklhauYBidCkeN1WjpfNNtpHpplyxLQFDN7GokZpoW
XLKg0Y8YLuma2Gj2ZTYl6g7v1MgbzOjZhnmY9U1xNCIL4cAGAvdYLTRof8rSafBJNbmfosgSQI6U
08tTWYVYtngxDqnkSsxtwc2BCsrse7lUX631rWBw+EKNtKLb2jMgwjPNQra9MUt6HsKRBgQWcUWx
w7CxErORHX+V5behQYttS2/+pysVZ9l7m8DSc/EpFRPkXTBzO4JusgpjN/9UcOBPKZ7TfAd8GGWG
tDD3Tbb1KR8sN3NnX65SAXfC3D2rMJHM7DzZ71U4q2N2CSiDZIoObcIfTvvhY+sJXMuMgT2mAbkg
HHpL+544gaaGUpka147KNeDVlofRcNsbxZngueX/bk1eKS1hZQNY5IEgNWgjT0nZS0HvqpQ/sVb2
pCuTy/R0lfZhqzcE8ZhoU5tuJk/QH2/954RyM8Y2gE/yr7tC4Yx6JTGkwKR9dG+sBEg/EzjAt/n2
Sur+kyK+BzHfN9dfnU2D4dImx3zP5X5Lp51Z9Uw2E5samPdhNtZh9bxb3aKONloN6YHcDKAFL+Xk
/LR/y6J3Kupeh/Dm/3usJJHNiYqok0oGTkbvXsRc4XpLgQAkA0/5OfmB4lQggKeLH5g7tg7ZjlAL
Z7LDOCbili9QqD5MrP9T7IuQMebw7JzGcY/i/AsrnH6cmX32U1HgCtdgXYKTK2POekEG45vIAJHY
HMC8AOvXorZ3hqCYwxlmHQ+JXkslIADR0P1IoHhH51L6QZjN1JEzdkUgFsQO7WwFkbgjN7bfFxTG
OsbMOmbwIzpQk61Z2IEeeI136XqZk/laVC5Zj/wt0HoeiySkSvarDd0JFzBqfLFkCOCue80D1K6O
pkX+QmjYvee/bEma8nTCVU7Q7W09IPkt2MXL6kuHg55QlZTa6OkTOmmlww+LgXuGx4inwbJR0l56
sNbO5PDYRv3NseJ+BleH60n02qUOAkikMnvZ5lJF9jRfwiBCwj7Up1TzHRuCFy5cdK40OmfPB98N
hkI70T0AjNYuDSH8FBa6GWhKdnugPyLeXzBUqNM1d8bAVreGbDaJIAlKPID+HzsT8KMXxtP8UbZZ
LL/gfpkbSzvjCTX23/R8sC+LPQlXCuaKBJZXeHG5NV9Mn2/gmntKMQgib1tRoqBSW50sAqBv6/4L
yrPzMFx41uzv5nEX7xPGvESRdM8bCSASnxc88wSIRcNei8jGhdyPG0/u2k/IwSp2l5TOYIOUINh2
l3U+u7jKSPzuBGhu4Bm6fCN8SH5jMS1VLYLrl3Va/YaH0n6bf30tpMTv9ZQv1YMXMFlElGKGS5jB
scLIt4wHvX4qX4/qBiulCVW6aRxL4XvRdYR+/tasolOznet7iYcbYyNBYWzAWl2dBC2Ze/8Uaq1V
kpDwPPTFqYjLShfHBrxk5vq1YbXK/lcSy50KS73M7hA7S/DW+aAB0inxSXireq8XPi6tUK/LmI7B
xNm9In4vzP9wq2m7Iuh0Fmfnv+UyfWvhiIKJIHcEDRsUc3ITjtN7ApkMbbifhrDsa6HYqixK3GFQ
PHYGIY1xXLydCWoP8EF8BkdZYsMXynVAtCGUELKAItiXG32cXFOkRH8G2/47wtYgpYs+SKCaaHI/
cT+jSgKkXIkFX7Fq0U09nv+eD3EAughngV1CZlnmF0uGOpA1/d41Fw+MbvN78Uw51Jdd1EP4QL1q
pnX+GtRR5vlqlzxbRDplAOBhX2k92X0OjG9a64y6IPRzjpNxOL4aDtrjQYCFaq8HEG9Cu7xUjKyk
lgZlwjFoLd9j6gS3D2QTwD2j4+VdKsH5Txk9gsGkHBUZGYmyY66+r2+fDNgKPYMphCk4qr67USk4
2vpDoSqo8AHVClecdvssrUdg8AxSPUdBogr9/Rrx/zqdekk01eBMhhDJ8dOVqLdZmR/2pAUoxPgT
uSXdf6Cm3n5ICdWAkg5PV/jxj3Xs7O0SOXRaKNHZDAnwsumWL04qSxa3HMiPQ/Tv6G4H8eQwolwf
18EEG+xHfvwIcY21ggQynFDGZe3HyibFfNB0oHCTAkYK25Nop0ieYAugk4r4eRr0eU5pkf3Gl2Ig
6GWcnJUTQt+EGyc/n97Okcp/3wmHJkFsqSRl+hLoVrqEYM3QMn6fMG2+39MHoy8fVzcLSQDtSA+5
cQPtGNmyXzxowm2ZNSSe/t5hfAm81rAPvAu83BqYsNwTpZUBDOefwEEKWb+3YIuiTd/zykGBIUJE
TOMD73blDsmwPt0L6G8ulxe9iQgJDA4lUWMFTQVScLH1LYy5sakpTGOYVTWRlkFzw04TynB2fXaQ
e9EZ0SiPengq2WGFuMTgSyaIH6L5tCtk8viOIevqOVt2Hwt4oo6b8kbLnRY+U+/a+rkKxXvHdhq2
W9ctjVZx4sP5EwFRG6f0nc0bD10f2NAsGpYUfVMs86IO++q0+3a8wvmfXqA/dRWUv3k0rv29SHqr
smytubfc5l8TLi5rhhZQxEbVBkPq4uopHw5f+jTFUaARGFX15kucUnwwtzKjPf2UggdxyTJXlCuR
cGpWonuzHVVT7B4W4p/TY3AJcraNURKdnfqpFVSE9iRlgfupkH9W2fs5mC8qsNl0z0XbWFZsishs
dFi0aLdvLUsIbm3IK23NDPtmJerh2WxT8kfvV9AlrI6F9jnXzjDfwXTCLjjoKFS5jKckKaaNqUvV
UVOyLRoypdWjFqNOlEjs1NrTAu8/myoGQnMGT/Sd8Se29MIH81HeAXUqpYBXYYmdARh9FFd2hdVE
O4V1hzmOWzX+qdBIBopOo/rq7Q6WF15sXEIoOhcmRaS94N0kxspCy4NsDruVTVeAd2zoTLSxnVVd
4ffMfXH8psyGgoebc/V/0l0PZjf+QebkFCTSH65wiLPfeBbtIcsYgvANxNEFtQzQWAM2Seoc1eZK
KnJLAZSRqDLDiU7P7K+T0BMpuSycS4QTAz6shW913V5YMpfRwKj9n5olv7Q4RMua7Eq4ZUTfgotd
xTHApeNBo2C/9xMbt26ZapjueOjwADdA9Y5QeKVDgegrZHm8tScwVu3iBo4Z2iHSE8Qq+ZrmADIb
1QxZMoIcGiunxL/A5FwIYpprUpR/fd5oXs/bPRMETBvi1tWR4eF78N0Xhl7R/U5Ie+s4BKqyTy5q
s8yqWZSR4UFhq7qrHvvt8CpIG0wF/OJmCBGlFBMJ7aPb0B58OQD5deJvSUZx5EBvigLMIqnc+ikf
GEaSzQ8+VAUHrRqVMVqUg/0lSVsuGUeB7DEc8xDdLt5bZGSf3W+Bhpylki5/9QW0XUc2eJn6y+FY
lM32VfXh6vY6rAaqoUdFzYU68miv4/BUQHbOFYktqZyUjI3zh4+/yKxLnXTRPAlC6saK6vKMfJTq
XwbF4tM3btpm3QoEXv19AMvhlQNIXPQ1TQTdmRzdzJGrmtp+qsU5bQhOFORIFWcdQztDjdzol8Dp
EUhabUtkQdEzSt1IVXTAZSdiDu4YgqoP74LeTCsv3suhiXCzHSkBFGh61OYvqDjlOUsTjwJZxKNH
PFugsUTWFsoTJX+XS7LnKHMOl1VqSk/3C64KX2LkSXCw+idYP5Lcelo/nkaMwtRn6/6/MitNlJBe
q0pvgAa9Kuts7dIF9U76VaeKFVCfUsY8DIV0jmaDJObe7iKywuWzF0tVK0hcvyyyPpwqk6NH/X0h
p6MoCGZ7p+GH0QLogvNdNVzyoGvRA/DzJGQRVH7+UGtQ1b9DvFH2CoJLPAoJnv6fEhcqku4tpFJZ
xrDAzIg9w48E8G+0cTxoVz4EdQaUjGgbC7vBnP5GmSyRs+XwV0g6uOh0VQZidYvCd996QHNOTQvc
nyk8l4oSK36YIUaIxEN6IRKdc2rtnlJI4yQ+iCYt3D7bW1+a4gtf7GZyKMCE5WrbVmXlnn3rtve1
SQ+GQP0ZP+TPThBR3MEMU4boTeeg5Ap1V6pLJCcXO2mYr4H/ihkYJUNWClikGZy6T/NeCYGj5Eyd
CnXp53HjofSAIqYSl7g2IUen5boapgfyqlwpogNoiKJVafKZSmDnpq125z4qH+OJ5xUUcn2FO7kw
GZMYzrTgAqZOkPDO09B1HQRfZHoPXaF50WWmSIwo21sZtzViAaaubafOqMEv0wKG00IF7d669cZd
wdJoXL9y9r29gSYXjkEhX+5FBCHGwOvFtXNpyCatqaSKNlVr0cqxlv1E7xAsfHmg463LWFV171fw
o0iqsDXfK6+CqKDhZEp1jJ6Ues9sVh7xBeJaoJpcr4JiJTSnoWLrNVus1DBImhOoLJcSnBjDPmGn
BXgFMQqIVbiqkvGQpOUZRFfEs4JfuJCKRc5SVz8nim5ejuG1ZkHG78GEjmG+7cwTJExFXHD4MrOQ
w8Hll7NuCAkfDkoF64JsSoMBaUwMAMi8lK4kuq8tH1Pd16XDW2d/KCdXxVS8Q38iyJ3T+J2SxTzS
1z7JNf4B1XRylqVl8oBjHxfwcHyDPF2+1hT4avhlVF6FEmOOWKZDyyFFMwcbI4CH6q2WvlPQEm/M
mU6OQroTw2w6Z6sq/dLLGuRLhmDjZz4ysrI0c7Q9YAyfJk3DufB8wOvKHUzsn9TD/ne/flucH9R5
6C8LO09uwpLktJwAALIZN51EpXxs9ATPU0nG5D/AN5WoUZ4ttUkEN6k3PtwdR75hQUtS4038h9Wy
vSGkK2R7biVRVj+N7hlN/FSYw0msxWUE2WcUo98JdcvntekvSqmLyice3wMnH9unKYOnVtUNfx06
8o3mK8c5v9qBFwLoJnhY/SRIwBG+zIKjMW3Lwa3lBvQwUmZeCIVzISMU/KUbFb0ZS6MMPSPUudGC
d6PxiArzJISMcgklm7V5Kt3iA+QP6OSB8cefkCbLL865DwK/REeCPDcCUL9/j44I27kcKZaqgMVw
Ds1vrbz6MjXhmAiMVP89xN6z6SD+yrzgS0DFejD1PI9SccgmYRJLwzU8tfGbjbYQCqZfm9sXtAvT
vRz+CBW8NcFSg4+AdRIgxk3k0vY4HREO8uBjC961NIE5WxuLXE6pe91I8vGQQBd356ayR/6Gfq25
GgNQER/pdaqiWW/RVwEO5VZ0SfPYImqbtvq9dX2TOzOKd1IEBhZktGkUfTlpBm/uIzNMr2zcex7d
DYZnihM4FnmpPF6cW6l5MknpMKlzfjgpf9WvLER2v8dczBlvD6TcWrX46rYLZgTDRpvQJnrF0PwT
eEJtx63EFW3rchNz22fTmTAgEyul9BL5tygsdPiwu6gz8AeZYicn6SepImcIh8846c999x6IG6As
qstK3wA69hlgi+1q2Cg3ahuQ9dxmhYkeGjDvhK9XegpdUFJfyhrw19b3cvbpTJR5hrwIDFqNr47c
gOZiIQh8y85/u9CKOPizQKuyOTiarNOS/AWgZLTM7RJLWbDMnDoi6s4djXfBZEWvD4CUw1rYmJyo
Q2EbvcTo4IiMAz2tD475rRNRsJUUHMjHe++2oAGsrxKbqDWUfr6aE13yBKgn4m5jVBqkxO3/eG+T
6C5EU5leVkLYJ+pZBXfNAbSU1XqhCyxwsghatLkermV+hu7c3WHsKuEApL1vqmo2jQxJuaqzBMu5
8RofTUj2m4La6Ab5VSx4/fO/owZC9baD+mezbHkECJa4yiV3sUOR2wvmieyt61Np7ASnLBsDfT2p
OVJQE2NXz6UAtxiOsY0vrNwSuHcnS4LTx24asRBtrU8DgihJnKS6c2+gic3Bu7HR70/ry92Jyrpu
pG6E7mhgfrJSJ6zBltDBTZuzvwgpvzs+zGgt17sHiOe25Bje/bZXs5vZpFEo3/xC7K/ulx083TYG
zp+S42eY/OjbuiZTw9sIHKdHsscfgoIfth31agE6kXu0tetQvXjFpWt88TdvGW0m35iTOowRYKTZ
OqzZw1kiN7TZBW5EnwepCjNqLVxfH80IiPA8O78PVi4NCFf3gWs+utVV7j7X6MvAz+9+NeM3j02j
JBw7TU3fDXoP6MQdUkdDBUtMRyPsuxIOWUoVe+iArZHbQBuXq+V1ut6DvZmrGquiNUM3QrjGeh7A
hxubGppSGXpPsZxOfm17lCjlDssknxORQyOd0gTpBm48JvXaJjOS1tYqmhEgiTz7QFPKYALWgNL3
3DwHdyziNgXFbMhITvh6fvVCeL1SMglbM4TlP2eCzXM2gxUSaunodKRv+RgPJ7IHIhRRnIUKqw0q
6MibK1c+IKMo4Y0LYaZT8CCHK4v3oDpwOS9BU1+zr36OzOJF0e9b1Is+C66AaBNnVr2+qD7Wig3a
NcJOP3qbx1lORk/D59nvdYOkIF347aL5i+2ANmQ3Ccp37lVa+TeJ5ly69sfKxN7T5GAhodeO2xvA
+ck9e2Hr5SdfQc4PGH4vROZmht2pGH3GKChbr0KUXLLTXRDrAPEbQRGGExRQNG59fbBIOdZ8ekvj
vjf/Snd2bd6a1LHtzTbUkJGD15LGD3nDzbT19DWezOYtw4EUEJR69Td9nYvKsARmQJbgAnkUTFYH
Bj5fgQ8qMpW7H7T2uxkmiG5wyqf1Gx5X6XDvb1yBzv85LAtJ2jvgqhgaKnuCbereBCFAlFT0B2Jz
Jc9ZACU384w7JVQvHFMWlPYDSg8KOGV5XKP9kgDrVDzhZziizN9NVACDmBw/rrY4qAWYXfjB0VX/
gfNxZ0NNvE3I37BORzQ/DlylU3giQ6mid+5nU9ABNaxixISg86DbHGqitUZoQbbtAZ3uyVzrlS5g
BQs8u8ZdGhCY94ARmPW0plYOvQBbI2ncXqMDzhyv8SYX/+shgCpmwlIpuUE+NX4rHd4h580bmavC
O734TtnQVkb6TtnclSjS77klMw9uKXeFsXMgWnlCqiKrKU1czv96xIGjbltZySl8G7Y8su+7fdLu
RnpczgfcLepVloH0t7WyY88RX57BQa9vAud3Y6TuA24yYBKeP/VhR9vRBUiR+9VFHREDge5LUAMX
dczxXo3vwBJt/cMOTb38DkZYLHw0F3nmXuQGZac4wyl2MfGMBiXM25OkAApRM3dPdzNj7ZQIkIht
MMkl9guxeSxZ7VVYlWVy/wCCCWZ55mcz+tWCt+ppgF4e9L5VjzFkwzDQAlxmHujD0UR/iFNDR2gO
I2I5epSbNwQPX7JhNVwhgyXWgXvtlYMnUWOl7aB8AH0dd2OQiig79pCpx/X17q65iGj2UL9R4b7H
V8ILOkbZE0kAbup3xfM3oOQEFMYlGCCfoCBytZXamtGU3gbLm0+0hwJr7mqGfDqLjTlqj++KvLCX
kjbqUmIoo8xV0U/x2087JWJUSAwlD16iw15kDRA9KCf1PT12XtjyK0p+ZxwkVqHvCakQZ06EWYuU
K/Qi6vc8gJA5oxN1Jsv6D45+iQ7VEnxDwOwgdIrOzP71D74UQijxJxmBLufXrxny3nRb4HRCkZNz
DakIBuEeb8k4DQUDPD8IkN5MhzSYomBR7nyGlAi4KXX767RTBJyjrLuSzdtLSJl8GwNw0yee/wtn
Py2EC/5YRncUVNrjQlDtmpEAEsgBBix279u3PTtw8qybFikzaHEYKFqqFngOPCWNsD5fbNbl6xIo
ooW5JSvdK9gBWiDNEsHeh0QBXPHEXyiMuVgaFtMH7Hm5Efn4adVTGTMn+EkyL/rjJWIE9NufIhkL
m85+bsmfbYgMA3KWGH/Y0cE0L4IJ2JtnlEgEGhULM2dV+11fyt3dpLFmJ/POgldHBE9zaZ7jRP5c
6Sr3duDk7F00udMNEiTmc9F77f9Z1iPlExbk0NMch/0gPXVbl5uKzWsLfWbPxqt924KuX1lagwp/
h7GRaCWlzcWCP5gW4KQU/C0IO6eiHecUQBM8mFEyabEXrLCdWxfRHeau0MhpOqvSllPNyUVPfOHK
mB0iP2uYY31qrUS9T0MOrvNqr28MmKs6PcfqNRFQHJ80DoRLJ+oi/6CKKRTs98FJi/sZhB4xZxh7
VXlXfNWHCoDCBwYfUb1bZfEvv7T5UQcn0IaHCeTLmEzdRO/EX4KSzDHWZDik95E6SFnVCPQo9g34
SFjfljVgEBXLQyYdsYmKMyGYNbFgqczxtIFNkDMX576sxuNaldWRImYOsYjJquNlBordbKVvJwME
PdPdf75lfFwKQL5Ci/ih9EOIOjTZk+eR3e0ZDvgGkxCXyYHUJv/oBxNdcM0RExehE9fAPpahgEfx
ZCK4XMsh6obWqVxgkepwDnIuxiT2kKnbG+fUim1trk/eLQ4cZkyp47GeBvvKUbtif8rOJHuZEeCl
rnMmCFpszUlQ5jN2AiTA6YankWh4CEa7F6uTXOMM/i2NXL4GL4naEcrufvWwwJZzGcyc8zjkVgJr
XeMNmRq2P507Mt6JmW0W/7lo3XO8zBp6xcb+h0zJlJ6wQPFtiJIJcvduwOyUg5XdG/7UPDm07tnM
a3Rtu3BqQOO7GeumT6zzQQsSDM5WnIQ3nMS5q5xsom8Dmxl4Z7ICwTFED5fWfvLwkOD+maDHSEKD
bVOoEj2PBlnf+7Y6eVc30BPEklkRzD9SX3m3Gc2Pu8yDrv65A7qP+l9D9Uz0riOx0TDrnO/R/niQ
rZbI9lsq9kByU8U12DhOaVqHlmrbi11r9mqpTEUod2BjJ8QLglh4ReFfvoUUNgA0gHofpL9nAJaY
3aVmld96Th3vNFaDqkeqSWyXrgVenbJqBDtaTmbG2fXBD4UW+QbJ1fBorlN53FMDaY+9W53+kYKb
ISn9slgbd3LEm6mnw3ZmeUd1wLT+AJQmvxcDDzCkwPs2D3qPcnJN2Q9PLRUdCfyXnaOpUlG6v0rY
7acmtOdQr9reFEHk4OyLVBvbjzzUxabNqpcJRVzvbKm+p8wroHaJukFl4PFx3r5HWknEogcOTsUc
CGL14W6OJlS1jDsjmstCkiJu30l+EKVNmj65EftO3QtrkzaM2QjvJX1CDTINg6afg871iuFfldPq
Gneog0wUh0he2PnYyMZlQE+GkkFLCLiQgg+Whdk7xVzZGttbzd8G4pNRFXWIBdsnyTU9ewAVJZ5y
89GlwPYTExL5V3nsY9Vl7C0WT/nZDkdmblxvN48vn/VFSOpjrfNEEW7CHbrAdMzRWQj0+I2Af6eT
yueT+CxKOFzXIrQJC/4ojrbW9xpc2/2LuclYgccBMNJwfA8+RkeRalGsMfmPmLPO7+aj5hwy3+G5
OpteX6cXse2tnM9UeYn+ptlLijQJx7QeBNnM43V9nh13h+emR+RBDNieLorS9aJTqpNzv5FkZbrW
vM87pEpQqrIO54gX8dlia8wnu/SbrZvo/1Qw3C0j85Ia47W71THBA1Kaj9V+PHFiFiIOxK671W+C
40bxZKBWY2eN9AOTDYFG75Gby4HN+Yn4lJx3mUgGiAVeQWj4ACBXLpvBWekA+6u8Fm6fupGf1see
9I8XjUEBBkE4NEHimAnGQoDKeH8wYwaRALtLpdHfDJTbFmjwZrNEV1LF8XJWjQtnus3h+DRQ4n2N
bbh+xIPPSENelVBNsf8zpQGOcSzlUO6wks1X/qdrHPBjljNEgAV1kfg7KOH1W5tI/yzwixzEcVUG
rNVNci7GKDf1I4vpth5RrF+D8Ci5HsPv5J5e2biTdV5bVOL8CNBZq4R/qj/cKOu5U6ztuKwPijzr
jNiXlEukzfH+cKSSR0fftWKcpNXq204WVc02WW/X7gazChIZuvoLhJzQdChCTZL3Am8c4lh1zprV
/P4YOMMLrNGTDOu3v+CDkQjCUQyXARPXEz3As0kdT1qCOhnRaKCvFPeDHH4JRt5IGZCTHpieySyB
YBSUKGYX6n6iIAhQi/biD6iwVBoffgGuCHVbBrJHYWQc8/NnKFDAbTGAAEtDXRa7xAJltUVXg1IC
E7ITKmra9JPllcmZVUwLDcOyLkXUQmCThuO4LXxajaJRPwhyHzyd0g43SB7ubTyc3wbALOtMby3Y
kqMvUc4VER2u2gMNljO8KFTj18bF476tbWnYRmTT5jRuWOtkTaKqKon+Yc+ikamTbDfDOkmNaQjx
wjjKjFMCdz/4eHkuneq5OPd8UHrNBFc5zQA7FM7o/OOnNbxUOMXUyCvhUAymVdN7V6Wu7YRlIQ7v
I71NXhg8tXw2nfkAN1x1eU4tLO/inJ8GjVzIJX6w8Ozi4GsJtachh5XFStOL5ZqE7DKwaws3RWDY
+lr2Y3y4fiwc2Lco8VVv33LlLnTe8G5tEu2ffFOJbZX8yPeYjWJSKjkS0kJd0xE1MAhs/eNCmxAo
pKYXqNqPZy/MEKrx2hlu0Mn592Siv3l9XadfvfqovAFE6wcmLh4vrOW+3Ns/KWL3yLOFE6hgQOjn
I07sq9Hk8eBaHrUwSwO7z+kGCANmNh81IIRGFefF5+lWMFaQz/0sX6lt0BQKbaGSjlnYfRW++Bof
1Nfeogw4rHxgZrdsAxOl5EBl3z6ub6QWs1Xw4AJDnBRGyEbhIbX+el46VTYoof2V2riFRBHWcnGr
ML3LWbSFoxSfMozhHGj/kqJ/9dXQS1WFbwpcOesvw49kCvqqGj6di7fbcP21027xms6Kse5bJRPV
nFU0iJktbOmv047wl75ogRyE6bUd57lqR+uwjSJFPnVygJjW0SR2uEgIvgx+2Euuq86H95SLdxTq
dLMHcd6kzlvgPjFxez3Gq5s/sPfg40hmTlH9ry8h+ReBmTSkCB5tFlK5L88yzd296raGj93TvR+2
AeafkD3eKRJ75N29a2S6e8mFg37/CIJgvPSvkljuQVFNQLuXSgG0pwutSt8k0UeCSOxjToW/SyAw
vAawLpXihTM+pcgfDlsh68/pbyj5LApSqdajDDl61Uu7eg/sY5Sj68lawsYkYbYiw/p36HnIgQn2
23rvtwuaxuXRWaqqZM+npGh9xgS1S6FItUUHtB0DdjyysWBn2nhO/XMnwu4zFWi2Eai5t14PqvDa
6z3dcXpH3Ljam4Tw9zpFM/M4+geOngawIWj9xB7BpebtZQMASwqQnZB2zg6bxppX2c1Qo2wvvH4K
hR3uAZkWTNy9iPF9Ck9v0QsdL9SZCg+MhPg1oM8R4ArStwBHkZV/pRgZGMRqi4GwkkVBIog82KVd
OJwlMcsbmmqFTUl/nCcdO8ePj8QYjAfYEK0Pkrjx7eWDw0wa58X7OeYNJJcGiw3JkO/E+yJkpHVT
XtLASJoNmR2SCoj9cigz4m5Mh1dzTZMCL3ZXSNoukY4wCpKbuWcV4BqAGYpIcisSG4qi8qmovDCP
hytdi2eM9X2oSJz+/MUaE1+v+uNZTR3lFQDvuF/ooQrfNFxlQYMbrW3SmE2zPAujKOTZ/biHDbie
0oySpFzznsvl5HlPXnRPaRE7zDg9RCxKNnD7ggggy0xjHI2zn14HVZKya5Ioa2dQmOwGWz2u7p+2
kKOCO6WTDHohWw615JOSitqUTxjyztc15QdbGCEW+BD9gK1KlslTJM1aH6dJFVINizwR9NWPDUYe
CqhcfaV+T2oK8AWKG0OIGd+JHdy1NNKI24jvRidAGSMxO/T4YzU8uxVWXx4UUJZYnYVIlaSmiDoI
bLJ+95CtAgmSpG3VYqQqvJqaAMtD84ps/gDLw3PhLU5+I5auGsk26/EVh/JSnxZI3MyveMv5yl3R
/LZnzXTh5xxssPOvcs+a3L21EpF4gm4tbZiaHin43g1ZmZSCqGXhnyDyMx05qgW6J9r6vuOz/7/0
xl0yIxmNZEKyYEXBON8KKvJgHys/GosQbvVdyi52g/3N5yDgFi1xx15StjYMZafO694oGLleHCPw
UC7wMaOCQ6io6YuQkRfeMTVxQsZCWdtKG8l3/KxPtpm7IdzxAeDAV2r3mkwggqrjdPrskJ5qcWE3
IxNAHar1cekIcY2jzfWPBRwEEizApRmRuesU+Uo2YB6uI1veRmIBd4nikLpQQ+Ia8b0n7prdUItg
aHcbwxwbgP5o6AMKmqS2uGN7YUOi3lVGL7rcxLugHZ6nytwcLqkrPiw6+T59PaeLCl2A7QPLFx0r
so2T0Wo4kGT8OOh3SHUgeeYxzFW7eTBRk7mABEG5Eb9OnCBrBDqnrth6Lrc827lWEAVP6pqw8fng
c2gKipoZ9p+ngFnprand+73nBE9kKR83ggEf8pG8X+3+Z4XxjO+C62JxfBPq4dDYTwWeTgf0m1e6
WuixP9Thyt5BO4J+fs0KsQnp5rXOx0DLJlpYGTYCQBxWzJ/00h25ctX1lybRsCPn1/HBEdjX54K/
9Y/Z2lP0b3l07+PyelAyUVFyCI5s+WiLFiUplx46aBW1AfVerwlScxc7remXEDDAdOhVcRjs3Fke
UNR1q4ULpu57pOWa6/tx+S4bN2dPCC18/icw9lhtuBT7ZOU+qt5n8ObTgcoGU2NxxCMioDVwDZCV
EP0lO6/C7O4Coa6tWmLEhH9bc1zQ64MFf3B6chIRAhfnZNj22d2dyoTM1JzqFGInbuRhMCkjdndR
O9ZxpL0AOcrc39+e5uxBIfNTzsj8OA49uOS9ZsEMayjmJbjGQOAagtwNlS/A0gGGjv1KsNr7TTxO
0TVSPUNq95ueWMyReqvfVmHH65DzypckdYVwWoUVlRNVicYkU5BckaOmhwK8vPd6z7/lXZBir3kk
nxtzmvbfUubOc6Yk7Qds12OBBgKI1avBRmZpeKbZ+3G4NwviOhVAn0Bk2eZgkJi31xImDSBpz0cN
gGROzBIcAJObXkMv1Xoroeqb/oAVJAcPHqF49MHjWN5joO7F3qRKwq0VSAid3NLL43M8R3pxbrZb
XauAj8Kx/H49AqfwD3Iy6T2iy/8WTK93gpw78SLD4bul656WIMSKDkQhZOXDi434GB4+QkB7JNRQ
R4lPqmKInqqjs9JO6X1y6Qk0hW44m7RVyf6XxLZvXr4Wp0sXb97wAlz+ou42XiNgqig+/i9NN/K7
ndQlsSLFOMEmmJRle9xC6BsxlLw+Mk6skOA/opOhkuGJekQT3HI30D0dJZwYKZs5e4USmIxwJS8a
VVPZ/6TFql/YuyhcwNV/QeRNIq4RAiaWEjz6Zio4z2SBKbYQ5fpBMutQbDtMBHF4z4RIUXkpqoXD
s3ibCPBsd+xaxV5vb6Yj4BYoiI7bWBVPAr59dr11AO/+dkQ7EZjgtj4Lfu0CRv1vBV3fd6hUTcUM
i0k+zjh/G2Uxuj3saKtA4eqM9Xk/pTxEyfBBnET2wMt6h5lHyO4JIZoUoY1H9z1db/qtSnDV+x27
4eQFnim0BH+4JggX1fhInow1fk9y6GkLNELhKAXb93MSgMSyY5gAIOXfszn6ibDQltFRXJgur96H
9H6ooo/DL1qOjArUtF54yiR6+WGhxk8H8Ba2bMnibwt3LC6YDH42PDKg5iwKAPPmkmORgK5I/+6p
m8kWJEmQVR365eV/TfEQOly3tVZ5xnehdFN/kihJys9GqNCFUnFnIf1GH4U7T4smJAyiTFvDxx8V
S9mErLyEqQBuor/yqkLZ7PPDZCnlXwOnLAnRBb9/g52wPNI4ie6DEzlFvt1gxB37PK/SVJJeZ+B3
qoQEVsRj4i1Fy6l//ASblISRm4nirg3RwDUzz5h1rk6BTwwVBs/VESg4Ct7W4zyPEOmqf0k9w/Ds
tsWq622wNySjh0DNk5XRpFlwTD23ybmhXpggi02RD4bf1HNw+yk7nkaprks6br/LiWGJvBbazUX5
hp8NdLcHYWdL/yhLZgjd1rChSGVa42nJzT5i9dgdG8vzlB4Cob1piv4evzWJqeaUmJ69etq8uMvv
0Y356DM36bsXCmqNOzwIC4Bqpajf2xFazAivZGYhj/jD5k379mKdmfTdCQUfbIRDWzaZcLYFiIHz
mzvwEUb/gEM+mQE3mqREABTPSrz1XqfrfwtxCzvnVzwxgEJP8fSxBRUmvdeqZTkj7QHGnZngbOvv
Ysqv/0EMcNNKIXJvf/dFvOwYYqIEJxMvVcCMJJc7wHEwYrNxvXJFrx4sN4mXHCLzHftOBPD9brec
6vq3WLRvKl6Qmh+ZbJVZwH53hpPydvejWWAtLPROCTkRWEJPSh+sYhItx1pwSr2ao8tL9rQ8C/9T
7WPhc5kCSr8RFnlUvCkuPbjfJn+RnA6/Tsa4jJnxmXLKOYSKfyiZg9PV6ATGaMYgPFR2QPaCzk7X
gONx3km3GlbqOPnlxjwqIMlsRzBhlD9B0oOrLYn3xAzfu+UM9jJhW6Ef6lfPyluZIMM4e+52t8pm
4p29EAhWZM/z8mH5YgRrQEgGre4nUG65oz4AB8BXqsCCVb8rBotYA4JZpo/UWwNNuMnaSpO6s8NS
sIBp5Q42QK+cBoIeXdg3dGbNbXZbwj1CUMshrVuI+/VhfxFXC34p9FeE66mBKosuzJDlnJkL12A7
NjbElzHh43G6+CV4bJ70CVCtwiajJGMmwCBLUL+ut5n/sX+Mpzh4H1IVbliqpiIHBBVMbIzXKsEU
a4k+1u8wx79o7LuiPciuUrEFP0KParVDAgtOdGsNSYqsRO6PE8OE7TxqR/jP1qrFONU080NR8olw
66xcc6AfVjQB5+uiT8wNrUwtwMjTUfMYQkk6NVksZ5w9VaoN6GycHpguqv2ed8levrlsIbE8mrud
9w1CAL/Ynu9kvo70lndaBrjAMrkUPtzKprBBbO8YG8I6D2Skz2iCINZE1XX7hkxI4j/XNu884qOY
P/hsEazlc2RJ7yuosmeXFXOD16EDxCT1KJsf+Zv6Ld712kM8/DsTsJa6kpagWYUu7N11yMK4IzjY
sfqN6UW/u3hhgWPU5CoFhNb2eoqr18N3ssvHVLMde8PfLZ6ZDeanG/kWWzJ3zMjgtwIcYZaWkIta
EV2bGgEmO2oK1uCO487C5au31ww3FnqkCpZBncENKdCgksbzuZcTJmmJWV/BP4CoD085DSq6ZdnU
fyuLXJS/OiO+yreGHhcdDkKgF0j1br0sZJtWm3DNZpUY6NqWknb7bEsQeGgnQ6bGxCvxD8LbuEOB
Oxhmy8BMlPoldno7QWTW0xWC2vwY5bI2beebjtgVKqBCjFgnJWIQGZzT+b/BjfJXdQid0yW4v+zb
sEM4htIlxuuxlOKKLAm95nnw4tidHztE87GXhBOrmMW3CuXvPafeqTwhk1q275qJNNuVdiG40s88
Ffa/bFC/zXp7ZWUijMsbMPk1bw5n+OO/+oueLaBB60WRFzWqB16G1+yYQiRzx8lUzQwlm12srAkB
oIpZFNK2zhlsEkGMVSnUOX9XfmfUAXLmy75SEz+v6fXfwIrEK0NM1zWcNzabxe1RjjdJOn19JvbO
32DBRIjFlgnfLuwMuTFZBqNO3BR9bIeqB8zy89SqKOW+pRZIlt09WC/Y3LUZpfY1FVgJDXCIfn/v
ImhpIS9DNhRl/ZZDakY7x3Rr75SjctQxBJS/4sBv/89R+DmyzFvQkZ+X3ICONtmajy3w4ld9ITwX
ibr/KzA1p2Snm7eLKg22bQcJHsDhshVljrUcu2oPYmvIGxhtokrV/LSE4rTGfz6R/LgRauF1CJo3
pgsA+VI3DJ3y17yDuNtUo3OSb501Jgn/kG6wr5Rk9tWdx9iKguEcc4zfli9FDL8buR4esyh4mjLu
LcCDZW/CWtKCmO1keb9fQl3UJcl9v9tNs7fjEVYw6N3fApeJarmIh7QQ3vcjNySRwyzto/49HjZm
h18GvqUyBTE1xDoktBKKihObc2KcIfJlcL6OIk1kLZFEatErAjiYueN0n0dMkKgkMp9VhPhwmtbZ
RtMVcg2jD0NDrG3tyC8cWtG/eUDbpZZEgxV8ukRIVLxQFpWoSANl6KxvgoU/jFRnB+UjG61Egnc/
OdEIM3QKhxjJ295pz2TNQeA8HYcd1OMmJaDUjeAS8KR5IW08uLexpST93ytxrCkHHyeGJDEsrtTu
3m7STlS7MZmBa3W2BFKnPK3+5nhZbmVNLuh2FDh/X+k8O+Ds38YlghAnNONKwwBDhDhhS+EuWUS/
NIYwif866Od7tHrDoMoQzxpWyvlMQyiQIWhuN15ePUxPaiZ3438RU1K0ZaJWpSaJYwNJE4LD7PBb
Ic6RrBbca8nMJv67ss2rU+QKRBdMfOVCLxazUafluvLsXN2oCpvQX7/TVe2P3EZlkzKThVUcYBDU
IF1RUXZGugQhTetKctnqIAMzOsS5wROrMOZxSyK+jWGUQtBXxR2JdgilSYR0EpDYwF9FuN9sPzDQ
B2Mnwkot2zqqtVWa6tKqyly4nIXHzeIOglZ8R6S/GpENG0KXzor29aqWtNwGCbysFq0vT0g+Bqje
Scbw7cZQ+8h3ysAR296pVRHGA3XCIWJ6mgusZnusT0X5hIiULGFSMel+VPE/bQC/PK+pW9m2PXw9
MBydIEdJPXjz9bWpuUYCvV+lh90Rmbs4U7sJ9AG32QcGq+zG/AiPwDkhJgi8R6TLL8qwLmaFQIX6
uJ7MuAla9auXe3fRZU6Iiii33Dw7r01moZfF7sPyF7pk6rVn21/MvW1FW2VNA3XHNbN/YfLspI01
xDeEOCzoK0y4WYak3142leT2Se/YWPnIYuiOiflLLBLiKwg5Ga/q1/VJspcBWSMnAJgqbjbWwdME
o0rxq3uRfVjIATuikaZcjmHILZY6rkhf4F+GvLbSCgETWd0F6NhTD3I4ZKHQGMQ8UfUrpgFdGvt2
luCoTUZ2YybofP+nK8BG+lzXJp5pXVGFCa087hNzB3arSaaq4VZG+Ohy3aK10qDJy0bFEIvLJd3x
U1dt8Lqpct56HgG35R5/AiAC5HnQoC/PwPplXhhpwZ6hJx2zzRtJPtp0eBNg31T85ao0uNeeVnf4
Ja2uzbL3QeyMeIpN+aRvt+kYd+ZLhLwEenLdfXupPnTIAljBQgI/dhuuSf805mY6GEcNdnkJr0Pe
o39XdjgbR/krw1AqGqrkQjsIklnsyDufbV6Ywv8JvbIA4weS+qAPfAmTWmZ0rm6eAmAlxfntBxTa
kfwWwdbUgsGo6vtCxtAm2G2w5EwqGxGWrXVpg5Y8Cu/c57oxVUkRM9JGjLmqrK9M1VqdLsN93KBT
L5x/dEBpubIGq9cPCSb94aYZPZ52nwgYTL5KKpxgdQVLVnwZQpBsKA+GAUxaaS7UCarDLo/ndmvc
De2V24ToBtxftbsPT0bHqaDh2fc9VS8bh0AmVxazltlapFSR4rRmR6vUEKlANASnJSvtIroNWdtt
po12jST8TL+HfHCM1UzJTmq7mYVODnMwZ9FQspiQLz7Ll3jW7yRdBPHnLuJvyq0FyEnEqx3qDP5c
v2BWsB+nafH26zRNicIGmyjK9P0cydYVc1dCtoE7MBCgPDHHB/aKrguVzWO8df2QpUoP+/vPwXfr
iSW1lYBCLDWdhviLfk7AndmbBvZT5cLbY6EDyF35E5cJsLh9Bk5GJ4EFbvH1bKaMhP3zlJ2eUdrf
NVgq4kSsoqwmkK9TEHvp/T+oPu9Su8kNOSnXfyS2MAvWerOc4vZIJGDvdbfoT0FaWYuplG7J5GY4
8z52N1Cdv/b6ZZ7G+MR2HSvgi5B1B7CHGCrp8S+egIwZCyTxAzU6+rSKmh5qxGafB4NiA46rEYSw
WPhtnoRN8vn9y+beUwjmk5FmDofHJCynOGSNIZ0mMDomU4C+evXWXBgtCPQdFL+7IFaf9QIuYW4G
R/rPqPDN2yy+r9QIZzIZcneuUubHcZIgmoqUYbALKF+WyhSqQFI9j/pY06vo0V48xm/fAb88LRib
7CUSRAtkgSe9LpIbKBR7+aVarX88mLZGg8OmlDz0e9kZGYqzyGVakovinpWhdjgIRQR0DzgtYv21
lPNMW82wNlyIxPhEq5k/b/pKaEXzfYwLtrXIZz98nv6w7Rf8OPGH9gJUI6f1Q5wK3FIPWviiCNRj
+dQdLHIh7xpYbrG7G0qBXCJ+5MqhkVTQMd6w0TJCgHg483Nuvh1D/zkIrLdjXbkn2BKAXZ9nGhmL
STmUrDtUfD2AkDl42kB7Pd35ATAL9Gj/Tx9eAZBzMtD0v4m6p/mc1Hah5azMT/aNcHqr3PalX51T
/KoK7L/cLgtCMkXAlaEKT+QnPZ9cGNLMGvs96CUtMcazuTSoFcYDJgH47Fq6+6wW8fniAYLov5gQ
hWfi7alrht8OB52cI313EyNNl2FW/kgjXl4Zx0VGXVptC2OZAEZbECUIamJTQmrLc6tz9+sBwsWf
9UhkTOPmoM+H409d/KiXHjVGUdx1hRrD+jMgq2KKyeurkJnHnkmt0e/DUzlzb+/PN6an7GEyfza3
yWP24y2REDHg/jjD7bPyTHiP5T+8JOWSpljadYBZ6UF1vzuBOcuFWHbQXXNZXSFaLaM4MYQzqwYB
q8jN5+dCH+5DT5M07dR/23MLpxP+t8BZs9LYDJNFK4CRk4oW5BwoOqzzb6UAf6sSx4JQ3qAHpQQj
xjG0pWURRXKI9irmtbikcgTR6uOYZ9bIrpxUcF6MImpxSCgQw+ZTR/npdJtq6LiLRZhAnvInLeAX
mK99szvHjk/KkLGcQMh4k0VZrCxKcUb9TGvrAh1LVEq3MesNl3R/X5ExL3TXkQIGi+uVqVkbaSQi
s09cVtWozTEJC2+OfLnnWtfLhTZxjppVgpRK8p28vynOO9/NC3K0JzCzrwVQE4QzhvXJ+Icvzd8B
FeVizY+M8s8pICiIx/gCY33ZzDunvbSxpWvviN1KnedvpjCeHhC1mp4bAHmz5dxd4QJ5P3JQ0cQY
AhFnzsi+Rzyx9eNtcTvt2jtfySrAYUEQAhIWbG9lxenAcuUtCMBtROIBUHjxclChcfhNZrRSjUiT
n9zmIOq4YY9mD3r4XeARO0v8rG3kBKZ1M00f7nJzYLNVsyo5F+d+pmMUNiuHL9trRuZT1rzV4NQo
lVxVG5CReJGCXI8COndCirG+PSV51OjZy4tLP8VkP2coglsaWyWBahOVFoCGcJOJwOWMSUn/UToT
dv0J1ull/2mpwqYTPpB/hrDa0R7XHf8aWqvWgtcTkCPxhFpRQc+VGi4XJ4OxpJtuv14PWitZImA0
130DNYlV8gasCJsxwFs326jMQL+qc/3mjYNtHsB/2YYSl7C6hmq3aPi+b+81Vzybr3Dugu56Y9Rz
2gGAal1JHZBrosrnLuNYSLi/NCdSrta1H/+LIxMlLBvngdGClflBhdyUnikPmkIDl9BgB0cGkXXW
1eNT/NI9UwlyBJE5dqW5cnx/Jj8cBO22Ni7NDpwr7m9sDU8P/vd9lEGLWrDC0S8Q4p62v5kYtoJC
HjLUDbOzW1wacaeoSmpO1SfwMpNMZzMsBjFndTjl6jWYTAEZaZxvkw51PWRO8Jdi0wCkVWzdXnnf
paR1z2iLknnM6F81lM9QI6j0rwx5th8l8jqJ/SRBUIKyFgpw9dY0Y47Fx7Dm4Bk/5MrMi5LZvC57
94SPhUILpMR6h2ejVc1EUNswIPOVqvcslUCpjBCwRtqE0EzSmsNxTcXFloIZlyYJnibrKPzYzkZR
UtsDdET/egbO+tMi2DSFyB9Mq45LJnVwhPziSK/F8XfHoJDkqmk6GMoj07ITjRXzEyXlJ5PorfJm
OZhsLl5fi3WVPIhuw9UclJ1LlT2l+bh+2Os1LHeJYbbbw5uATClEBsIiOKcUFXrzs6X7CiY07nks
s4h3TDMTDgZ/V0CykU0MrZgbeSFSuSxrFeLi7997V7blm4nhIgMNRJQZ0NVmEOUCy3LN+OGty6Al
pzx1Sv55DyphnpFKF0Ja7Z4aADtBu5pmCJFyz8t44CEy3erCGXe5FqhcLu2bYjf5Dciw9dIz5sEE
8weFh/bqZJnu4Be4ojXnStA10sxg9qnN+V+fkh/J8qfo9UGEPNv3bvV1OuE9X0UpEBfmGeOcolzv
YLuKZFhIit/KMGM1HHLmMPs34TjMB7T+HwCL1RFiP/Do5we68DgX314gRDdvgxr3oyuoASkLOUUY
/BfwiDYa7TufLeLFpORg5x1Z/KvB2IeNPPSshOSK9NQM+L4ongkag7z3tsleuC8UrB9PNoeM0IqR
c8adQTJ96CfovOVAiH2Ig1VDWnIpoqXd6yvpxrPVg1V0PvGEkTHPNAp1wjgMRQyavr+BhjCizuHO
kvwb4lkjmBvedSDVw/fnlcUHAQQWQy43Gxsu2nAWVYJ2gg5tTBm/lnRDvwBF3tQPXs6MAqRHkv/Q
1+uC9eLBi8hZU7v6ZXxKL9q9Y0SsD/Hu5G6DVYsOBvjvj66qQ0IWggyjIjUPlerb3fGZKMk+ZjpX
Hq5rC7KHGRX+EVdWHjDFNMettLtTowUsZE9AGQW7FZS6/9HEfw0vpQwgEMEK39OY/PTHIEtBA5hX
wCb3npebOKHtUbx2yehm3CzTXOianbeDftLiC1hSCg90AzuSyw78vtrpUDbaFsLD4sPGDUBkXshu
MUBGyQ8M01Ln7agO5OsCfkmbSwdRzm8sBGb/gEsuBIdBEbPZHCFMDdHql/6e5FQW3fH3cYoTMop/
OEJ1G4d9eJY3FHQw56OvQ9omfp3DPjbbPhIZReA5kpXBO9bbSspjfln37E7qQBh+lksJC93blKix
YMURS4MuhMfYLYrY/Q1o308Ji73Zdhpe3+XjD8dlodpMjLCEZH6bPgbZgjkm6n1+gaSrrSlrCOaj
cUOFKZ3LlEyEaqNWOApfugZWYpH3FvgLD61Ss+kuGncwv3+hlz2jZRhLz9yl3IVchqsd0Vc3uAYH
XYu+fVyN+gDogIPSUMjHrmxzoS9DZfaw1dCWW27FtVyCC4UT0Wdekw7kP8VhFWX61otChCWGtJCY
KczaFr+ZGDjxSXx9XoFmBXbnqoFLgOEM6T4l23mQKHs8YB/vmQhxXWpxylN76M3NIGD5U1MG1WqO
dx7PudE/C/jMebXoho87ldJVR6M7R7P8ZeFCCcgJe9VTd+VHZmt24WVbtHrKN3LrG8OgSaTa9jRG
WJw68FyB7/hi3rJktR01C9S4NHnm4U3OZEh8dhO8ISYycxZANDHmmXAhv0PYs7tUmOACWBW1mdnQ
I+cy4rj84LQTnZMTWCiGWBdAikiQyBxu8pE/2njoJNLYZibzfewnSPiqZTEeJ4GO/3C8ddfJpIkL
o8rkvevzOZ0g6tewb0HgFbliCNS+oiLbUSLS1gubCJpdmOcH0ByrNLJUFghsGhK/hVIkldeb06aI
n8lCOBLwsyfIJFDm18fbeF2a5VUb9jS2na8ViqUcKV0Mm6zVmXinpEsM+2aUNvnr13s8tztC71Qa
UYSBkWK3RqEI+n2X/K75FtIi/IO2uwpdOZcWb9hOzQeiz+wkegHTdzw8KH5jQ3rGzT6SIWmkFNem
nCJydQw9nfnBL8EoRse+brqpF1uR870xfNxd95H/SUOaRNKwuu7ISYaXgFz4auP/s7IHK0S8Bew9
Gs+6amkn2/0jvPTpKFjDTk4X90TYvIdLgPReAkoHaMkoGwtTWNB7s8EnEMxaHCHQsr7C7xe2ZR/9
LxEq7wpaCSDV++i64iTLS/WRcusRRIy8V//aXJKP8yRehU4zIRKWQEL0ZbiF6gnR3PoKf1JvbguB
AAj28yv0DxKpmnWomooSc1oFWMrAA0H5w6ioRD7iOVD/WMiLMuuGst0tQi0IyGMp3XaDQoZaWumG
1Gr7jidlpCOQI+VTcj//7sKpK0uAqshAWILVF50DLxEIpPmmy3I211Uy7yVGhgdpssk/XNfZZRSK
SQ9zTandpLLySqjMm8ilQgbUWXBf2N4zZxM/q8JUJB5nY0MyRqGd4VFgfcmUqrU8CfAIgrawdmOx
q7DfXAEjdRFKIpIPlA8qpy1mF28R7hu3j7KBCSwEg6sdvJsr8lLIRHdMFZZRSfO8VglxmNb/z3yo
P6kYsadA9jJgPQgyDdtVJsiOnixrYaHsfuExu646hQCITNiOHCYxdlxumkFbAVGMj3tHZS1y2sG9
EKrMqLHWYGOuhWpcPUGkVILdXCctPeC+DwcQSu8wdcEuok1KWGH6y+khU3kjAvu0xOe2Vx7klnvi
8EfwVJSiKb6hQQdFGueXscC4UQ0kdrpN44nYO4wYbWSVao3HbPhJdj3XcS/9kajus3L3olqdt6eS
YDpInnau8JovuCeTkZX0Cdk6qMfmaJZsc0rc6/cCGl0DtbzyX8jQxoKVA+J9h0fvZ9nNvX+YDcKK
lVBTkL8VfUrmloQ7UOfMvjc9l/LPeBcIFzYNv57KV5z3w9BG2h3FxMEqJqiOTO/zpCkI/ZTDniEN
99BHPE1+f0CC7gxRp3ljttHB7pCEp0PMIFmxsti2LDbhdQuUErgUIGJKyTWJ5jquPFu98hsISqZ4
0dYtXKM0GvuNtELMJ3wfwDnA5BfCOsA/tF9w+RYsCGvouFM4fGG7N+TCgxzylcE3PjZSH6GBDVoY
1cHWhqQdiwKRAyLxnNu4jYVue0vUwwdR+nEGAgq6PX6aUzzILiF0Whtywjk7vrHdDV7zQVZHYUnm
hSvzdXaKNP8Rca33ViV2vs6UDD4ikdotNXokhfutMeaiOSCVvqUHBZFgGSjSbtacnXFhgvIYWnf+
Q1l+JWJaAk5ifO+49MIHJFvP6Mm5Pgk8NSUFOgl3lxYXlQGAPVlMbq6i+0kMNVotPGbYvYyKIvjy
HWr/iUZVVv/swdV8wQywVjWxLjDT18MK5jcz3va3HgHLGPMjQPTs74QAg99ePoP3yNJKler3lo2r
n9FkwvfsRs32JbWK8sxraYNxhXyypu0wZDGPXXQXbxSmsfPD5CjvkblNF3f2U4x38HS00AaUUxxG
LyI8oJd8Oh7hbXDBxLD8Z5Sg/t36FSL2EcVTM50Mh3Fv463MEl1Bv3In4sXG0/3Zy5gudFacQkGk
NzA+UAWnQ3KL3dfnIaRGKAx1SEOY9seMZz7awoki/laE0fjDtlgNncaTVY1AZpnYg9jmP8+K/0pB
+3A4ZGjR9+BNOG85OfAs0qvGcPC8HkpeSnekNdgtQeAm/Xbf7W6LipTLFh/OfsvhKjGGbdUZCtGo
LkyW/l7JaZhRUTS/K+Wax7+t0zl8EepWH/veKVMAw+H/oBixYnn5vFcqIpzNKJDVrQeFTbyaWbmA
etdmU9UGQvw2n2Y3wTtkdf5OIV+9cxbiRQNGtBxG3gACYcF55XelHCvMCU3WqOSL2MhxhGvNt+FK
F0KRH2p/S2eyaSe71say2FQJTyCqWVfjtGpu2JUqwb4RQtPToEXSVvk0N8ZxQXljDoA0llaF06Oa
7FeJyt4c5bNbVa0ycpcHZBthy72pG26QbrXjI1C/+eOsh7v4eGI8DaAjVabHMUniRz988nVf0hnw
5rfnbuOCVahCZIJ6rvNMKj3xUVSVQNnBu4RWkBXqOXA3dwyKH58Lm8Y3onSlEOKy96uy81jy1HgF
/SjD35ZYW28up0M4/uVrSnKwNLlS3Bn+ScrJHF3oGZvHzHacA1EoBxqR8siMzPsBhDgoN7ugxClO
JwBw5v2wKohAxDdBJaOXg275kVSLdvQ6lJE1SIqA7oLdwb+MxvYp3zDSNblNeI/hKOZQ93NaFaTI
OJfWPIP6QsNHkn7XgqIDCyHCV0/tORfn5CLC7+MobLdTlBgSVNt80IedUoMe75Am8jLX/LUGNZf3
4q/kE/m9gBI/exRVuNiiz7ZRg0zX+ON4oxu+JX7OHvTTsyTHYUb0V0IB0C6ffzBzeWVUUnzrtJHC
hQu6Fs359xjdjVuQ9VxA67R2HaCtP3GUthFo7nbPbLqZC4t3SyrXeJqV2eeksjID/E6qJz0BNA44
pdWHY7tjINqKPI86ym9kFiDxx2fikdBeP8mDxx6I5lIY8rdEs5Gz+6Zu1W4ynOflbpRgrCeCJR6e
wwdMXFrJ+hskCoz+Gk5zr3jNY4xGmd+NEK3XK59hNF8niGyVT/jTq+tW6QESPNGVb5zg5cX0NkPD
diK/YPo+8wqLoUCJk30oSMA1Ufq+OoiNy/BdutHP3SiJRNs2geRR56+6psvYvORXn0X3ZuTm0tt/
iLJe3vzAsf3Ineg1jqyOYDI1TkLiX0Que8SVTYSdHL8ceimHmBZ6Z+b6ODmBpFQQHGuXDtTpKdYp
QmlVYXs/QqiIPaOOycEZ+In6oB9iuueAEMXh6cLfWEMXASeCXROwWJyiLt9DZTEIjGbmDk3LjTQJ
JIZ6X6ezNKBNp7SX9mOXZezBYzHwH+icFw1XzLx98b+qn3hlaAhXtUCsNzlLcmJq8R5+d6IIHICC
AlbN6ZCcerxSgMUdWmIEfnl/AzzwdVcsxrLbFP9AoyXF7QIsm4ejh8tSnYB2sDDIv4BUtOSaABQC
Spz+RjlaY+qabSTlNhnF8Vilsw5H1QN/11KNBrIZIxD/WvOXrb1MpQhI5D/hFnLu35ypdxVYW0Fi
Dq09vU5XUYOCPxkjicEq7dUFnyCzoEVy2Zl/8bacWcQgTZbFmE1nrcKygDy3sFLDytDp8OgYYjhk
IkzCAhPAVG7myhrI5E76Pf/O1TupOq/QzBL/v5c0M9VWZAXBTpWDhgn20SNZJl7BjV60M4MH8IwA
PhbZGct56uAiNz/A3wHsXsEFpmK9CSDlRgPU2/MhqQeH2dTpqnBe+i2R8FLSnVKw0rbO77t+yDe8
KQzo9k0MMr4hujN/0XFTVO1VHykM19OE8+L0dumTY7Bc7IEuIeJ28/3BZso80gqY9EF3/ZFNcsdM
GvCi+rrEoxnr7HWkPBEqZxEhngnvngE0Ze7Aqq9BaThJVOB7OGLARNEas44VHcPBveHGTvUTUjdC
L3sUXUhFwN9LYXBfRcid8tZI+tWaie1n0cwhvtwBfNqpToUlBt0A1Uai9i1kE0ywPHlW/fbMNvhs
Gph5E58xR/RTEsc2J1KPe/SueGiV+7ZVvsFa3MWSM4jTvnuiwRFbTDL1H0AUB88agwgF5OKB+a9J
A6h3AqpLXSztRk4avmUnL9OcI7LMHOUzh2LyVGO87CF4hN4fkB8izZkhRn01HH4yJLB6tE+v5Glw
RDM3NTacmkQJTiAbAV+K8EXQ1qrWYVHQRr7MsoTicZbEMsrD6RObw25SW7ooZ8R/H4TooPIEfjpr
REhFfqSmz72+41lQFca1Eb2n9Ib3fRpHhNH9w+blSidAbzt293YKPzta7F7HfHgSnX6a1B+qzm/f
rj9mew/yeH+jfwL4slYInAn0Obsw4ZDLop7DqzR8nlvHSN+6GFBlhcBQAKTdndFswloNufJcJmbf
Wo7ZoQ89ngHYfwSu58slw7uU+lH26ptdrLiWnnHlWYUIwk3+rfMGGT+xpExNZrmL7cNrpdUJMv3G
whlQOKE0KHpJGrOLNvBQGIFVQ2wuK5crwN+kodpxf4E3eNopDEXEKYlnEWYBQz88WDeVejIpi9FR
mq6HBfLHs7F8qYiTtt9xQxdEcq5NCaAANCborcZctkcLJD6nZ8aV27WZF/TDECJ/ymGY7YoU4lDH
dBQjToXYK305R1XHlqBDoeBARg7j6PO932ZLoDuF72gqdFvU2hZIMKXB8G/xR2Ssx0wyKcaqa7WW
HXxyZrOW/jZKsT4X7Vkz7K6sHupgDT/RiJbSG0h1XZloV7XjKuyVlPJ2jcEjCSjATlms14AMG2E3
xxWsKYEXq3GheGMvTRUTpTZC/h+2wD5EGXw28QaXjJbPq5xDmAv2M6oN8GT7iVrtvXh4aFIy0vDY
PsZ4wCP7ciCj52Hu4YZXkZeDqCBK8gHaEAqjHw1hJQlXqVzpvEUQf1qnKxBV7efpEzfbX8l6BAX/
cADNjV7ivyO75hC1sie1Yc8p/536/yOtxm3rkw7kj3LuE2MdlnaIHDP5sGWUuY2PNf2+YG2gCGpm
WRmK98zMmodiFfgArD0n3ZG6Y/w81HaYG1mMfY8Jhk2Q57rl4qKIWuITy6SDlU4y0HDiEtl/+5PG
IvCq8qio97/+lI1KKqhjdXEd1rKBBChadDDUDDaoq9GHF33rh9fcUKer931gERxoDrWkXs/EIGsU
vLVAE6+aUq73+HyjVPfyHBJEEH+ArBBrwgdXkJy1G7a8M2TV6w2SKxcsfkv6qXkh12GPUUQLay9m
Az5wK7W68dB2ikYVo79jHSTx6LZb2b/bmsw4n6618mX49dRTBA/AYzhNjrOTttvqlAiIVr9rBrrl
ep5r/rSKmlNk3YKgC8tUjJFvLmeLOZ6GWUvnICd1RAVwHcbLI5aftDv5zZydNhBreSeXexaotbD8
Pf7kfGlbp0OfgdPvHNEKtGTXxg78WoppVLPZjQWH2FHuE3uNWGl0DDy8K3nVV2qODLxcd64ir1hd
VusjvsckYb7195xY9n5lq1mKVj5nEFcEueSr/iwjGh2T4ONi25LKBH+Tn6pXiqF7qPIhgz3d8I83
LiWpk86yU7Px0ZOR8SuMVgCTy+RZlV3yhGBur0kDG4Z34/E8XPWW60CB34uLnu88kfLAR1hce2bZ
FUN8O65Tu9XPxcz+l9n/kJT/WtHZbWTADaVeJVR8716yvVDlsChNVmbFQrgkKPD3pwb/rK/U9zBE
op7N3U9xojXe2dzAn3T2wKVae2w2d5ejKjz59xhrY57w9Rk1fVdU1NErDCV++lUOlLKqXf8n+y2N
D8Wy7ylh2AyiXFgzCJsAHlJ+Bw4u3wk4+HW9tfP0g3l7m2G08IuZj+Xvooqb3kYt0g6nIG32x/Wl
DX4ZAUJe9SO6kTTV7nmjOtFF3q5m9O3e4UN9OTWZT7TncV+dftxWzJcXnPkmrrFpfYZzKXxNcNyi
ekEjVliBNWl0OsTBpjycZw1bNehiNrmeAXP9QJqAZmJN9rlYP8bk2/2V+ugeGWsTW8P/ppBecRgh
u16tIVvr5DWiIFPjrtacKeDMF6ErgMn8ovNLx0mw/FRWawjlxn+2I2nHu+c7htYspmXiA9Ynu/Gs
aQBw0gpVOf6QdZol1KUm7fLCPemKs+XXjE/d0G3maWQO2NEdeTnqxZNBx8SpR82Uw0a9vIfNMGiY
dK4VopggajlKopPGGUVMeAfWoh68qzIRKKMePS5B1iwmdBDHWYgRNdn5VooXQts+hR/LGkFNrwp7
x4OZl9bRyYsRmNtsIQgFNJLElcqv1kJMKBPiOs30FErVplFhTTbMLYAjOBnyc6HhuPgJMz+wDcQ8
xW6uPS8Bf2CV1nGlbdGb3FBDYVVYJdQwoiV6YqPTITX4az+XsAH/ExMVUI8Q/+CScbn3qyWPFWc+
t5bMKcfEBwY3N1DxWU7KBzjHsViOXsVKphruBWjzLT0gwhwrRiZwC4CKwnSMEYIr1bWe62E9Ve52
YLLDXxRWgSob2G14jL5xLwtEP44V9ehHTPOFZE//bOK+REziUfRrKeZQV3Vk9rf3dwzBgj0WYSBV
BJJuo+2AbzrqIuQBPlv952v3uY+4m+Rxy4Wg3sx98wODZ04HlB77+RKnZ5/ZVncT/7p0OPH5glRt
gbULuWgJOf8wGFcHqqgnjDWZ3iKpnA0uBowdH7mzFGjdTzIALV+BN8jsvag99LxwfLjXkTmc2H/Z
J0ZcUf1jnCF2rTeAUlzHWSH4fxaynh0nTzeBGKzLMz4GC4Wh51XlmEFkwd6y1pkj0+mIzvVUjsYd
9TYxGU/9kz2PsG0XJnp0IT08jn1KLsGxDAL4x1ysyP6lNiCtPLRgmY9UgXbIXZPfT3rYIJ/DzCJ2
hzX1ZiXINDaaZynmA8LDrXbwi9yjnRrTsHWoEpSCxYv4HiCxeZcHTe9IuFhnjTRntgxukGH4LYCm
ijMJnEW7Fz+U1nKwRREEFUvkhPjVakNdnrCQ5NzIdqrnAeR3ssbupNtJLHk7EEOcwkt+Sq+KFM65
x8pjOv8hobxKg6piZrvjvsVodlcp0XV8DpXKneulP2XbamtEPttxr9NtLOEAMTOYI+t1oL5ic+Dt
BrTeg0j7h8WBxR2Ae/qP9zaadcFcMqpn4cBkxpYKAlX7L0Z9pjbAyCWJqozn51cx9j0PPieQ3P4o
HRrDEZspO1PhsObVJdp5I8pcGAkgpUtcKVDSeFouVrX9Qf3nlX3K/VU+U/wliFFWruog/7ocQ/8g
ZH9nZ4rvlQS7zQeenXSYSiinw8ctQVYN2DHaV764nflhviZNHfJf3pggTGQqmKk74EwIYWb7R8Yi
uqirnJWYNSrHvOWcM4zksp4taZLIskWJZWokDkD3D9KUajp9YkpK7Tw03cIRIHNOmuVYZgBWp646
RbyMef0ZuZp4Z2Un2Z8lOyJJa+TkRjWDn+Di27QAz3xMG8bBSraPA5b5u/dbU0BN8ggShaklL05r
29K5DZE06ATV/uSxvUJ6i7fQMAgZfCbuknlBTv+ggWIrFV9/n0B6xskxAaCeMZ8JNMOy2YrUckrZ
TmN180sFlIws/QD7GG6YUHD1z7d0iafx87TVvtQvyIawdMaCu+II+vm8KD1YFGWr3nK+4OvdNXsI
20a0D6cykfOsvKSqUaC73+OqrJWwpnyXYwi2snOd0oRJJjbQQf2j+0LaxS8sHHx6lCGE9O624Yvq
MTzt3PVTLslRJMhaCSeNjjgGYUDf2UdcbwKGCpkm55EGmIXN5zB0H884x2nNjkKxaNTq3IV0dvHu
pHRktV0xCMzS4OIxaukWZqPXCpd/HJ0CtQlBkmhwHs6K9iPrb5OSNRcI4xkFoIB6PwDT+W1YGfoH
FdDhFi1vvoKF8GI231+gqF+tXwiQflCX40U+X/3hr4PwgqBSt5lKzAQynWInDbJNc16bB8zAiwjo
Xgv728+8GaAGC3ZLjMIH8ZyG1Cp6fqelgXqOMB7MLGfgHVZg5Vep1nLpEUI0fMa662I1Bk2ysC2L
b+bcIyQl41DC2D5iuRl/0xLsfMtIdBbs+wsBg4hAQD+ZuiAVrv+PKG1Rsc5Ht835h++gQmQh3ZUL
kg/A/XeyOsxiR8cLv2rpb43/c4eZv42W9hjfJzG4TtDjd+HgccBXMakWrD5mq5RH550OoNWqdeMi
QH7yUQqAIEh6mY74isXbveTsHctxDQf6Q4yEeo7+yPrF2wP5rK5q6WtFcH5BhFgTOYFKkZ7SpXGt
/mviTGX2cK/P0O+LSCX/sB2rWeYEo3oN1VkY2Sk47GKgcJGQQ0DDQNb6VPMc66oLrDB7/ES/c6v2
NoRKCIVApngr6jWYXa1W5kFTj/qXpWvVHHFQxKeOVmzTbL5wTRQOJXHWNFhm/zCkWLieQKOfGbwv
++zzPsgOaRA7a/HSgR46y9d5sQiGYLZE/29qaN3JJ2Qj43sgYo6w6UP6U4l73Wv1qLcavKBEhoib
X5Ie6UeP8FgzCvVA4C1WeVg7tEPpxVMDD5V+nMn14txx9uenjBOR2mD2dLuZTUHXOFknnaYzk0gP
Ee8qwKUSlz11oct+JN7XaQd5j8nkhG2Gc6/GLYwdpWX78bzqLlMmPk9VjP0j9WgIqP5rrdN1XIam
KJOP7CwA13XNVZfcjAYHECsW0T76K/nwo5cq4wnV3xD1r4JcgTzxZjSdzO2wdRmXG8k+5eLEB4ZT
3wHmJd3XMnSO2MPMBBuSs8T+mIOVGTyO1P9vqaguI0Jr6bQj52zjSsBFeuiOiuVJffsL8T5RbFOq
GigiBc1a7a5eA6cHl25qfBL19RpXkOHJ2BQ5XCyHJug8O4+R9ncMc3F0PnGJfvjNvSNwm/0MOGm9
IwtKMRyUXEgD2gaeNBxTqFIljX3NjlEvvDET9gTphcJ1179EKZ83Gj7chDMsK0J5zq9O+rsDJR06
DJ2h9VYMBsEvnOrdjS1tUVKZzxp3/RGsd+Y/i8ycatB9ZXjN/93qFElvFnZ/M4EX1FWbZ6Qq6RlK
yxbe4nxWJJY+staCTkgaEq/8/sYAJBJuhfBcxf/7DWKWv0WczCvzqGCy5m1ujj8jjyBJaotWvdLR
1LUJtEPqFgVZ46tu1KJrZfngTYieySUEiKSIYt8R7nZiwanKmXypULObvSVdUKIY/ZE2S34AR0x8
5ExS81cYmEPtGlEV52p5TeONw+YKj4YVNWmSjLN+AtsAf2krAlV520EWd3/SFc1L2vkt4xAPUgbT
14u0lo/yZpSSlDQEUQkoEsOSwo6To8FYlgfuij1a/bjHLakFv8W/RQogMHXaZXpzmlZvKDRsiI+w
TaD1dxEL4E/FOvl/mLTwcaqDwtKzCApR8rh0qWqT/a9BXCi2jAwOqNtuioRWKzPvVlF5V97y250V
GXeVdsidXicofEt+OH4h0azfZtCc8CeDl/5l9pIwioZ4XWavcqiR6hAeB5DumUBewPcqn0exhGhO
ymWilSu0Dhhuh2npwlfPgAXCbJBhAg/De0HEvL00sDzrz2dBVumh36qcpS8RWPNA/+qIswoGH+4J
tSiwfo0nJV0yaQPB+A4Hb3qdY/DWpBuqe+Z9MBPPKhdlIQ2QWDa+wc40nJIBxOHpDTRHTD8Jni6Q
w+WzUQaMAr/qJQJ6xp2jwr6WE+kIxR6a0SDXSaG4DGhj6JQbcZR0TS/AVsGWdRmDsrqMi/ymwOaJ
wyu26/nPVsZwkHEvrvDLisU/qkj6Nkey59o+ONI7y5Pt/iCaGeuJkAZmoxsgjcbwgfEezE/dciH5
qVQP0Ybf7nfQBUGMV6nvc6J+GV7o4mboIQ8XbKvonX79HY8PP4NkGfBG9TSc6Oc95HKJdsZIzQMM
xdpOfp+CxbZYKLIXD73s+E1CkImz7SYUGNec8p5h76c7DisXKVIFj52gZXfNtAgDYrYYDXLy7ReJ
tddxU857MJxK/LbmV1K3EsLySJMznSTj31LA8a906YwOfqh+AxE5knCJPpLN/NHRecL3efG2nVu+
mRsU4P0o5gWPyqZRYUcuCqC9K5DUgSI1srTBSEs8SustMADwQ+i2QZ5fHeWjdeSqtutdGK1uIDdY
O4CFxiqloXXovGJPXWUVDoKyz7GiL6CUORq+vESg63++xC7HM+Kkt4S3pmCz+t1MsfJN6IE2Cp5K
kD+AuyRFqNYMb4DjBbICI/U1b35I8zXRKa9nW7aG50jLo0VSnmenBnfZ1R/SAYpA14l4gBuGVscs
74gLxCq+tDCNXd5Ozhrc/nQXNeRuklhu9HkZ4HkvwyIXPAjHkTG7IO2MY9fGj3SWmFm6tagceacG
zzrLqxbyxXaSURJSICZ7ZAdJ815h+ABEedU7OGGYFJNTBWOlt8gmuwSlhJqNxOxFwCHmC4XD9sUX
WJ+KJCxtQa8VL5LW23320BK4w5sZOfnLwmg44W/72ZhR3m6mkTFzrf1uX81/ygxNmi0x5maDU3n2
sq8FPaAv0VZeh58LAu2aGxhcmsFalHq4duxGrIpnhBnj2WbBqJKkeFDVuIQabPt7ioVOdFSyx3Ha
a/mFps6D/UH+eOa7YT8PVNP1/tnWuwwDKKa9KBvJohJhXlTMDXw8z2FubSdR/8qRiB8qQyfHmElm
g5hmPf3+J1NOCwNm3JIbrlasIa+tSebJ2dQYHbObxCul/fzvTqEfTtB5zpBCWP3RAbGaXUVdjZHY
lkYkWiNcfFgII8+oErIIigMYBCp+fRLnBm33AEt+gtv/wb+sT3uUeTJiC8igXPYDd6BflPHDf05X
QQfuzNJ/CfzKM5ictqprJNx/N2CTdjWg+cCWs+8B6rUiO0Aw19rVE15HvSgMF6u9sh0O0L9L3ZGh
65q0ZRiFlrYKLrf5Axx5aZZ+hBqTGPerJRCqX3528aMBzkNgSZGeyhNLL6bvZP5GOYubmHIGGBCo
4TY02Q+SiseRxh8u2UZxBbHqvnZRICL5RnDoH/XCDEi1KIfbQmDzwyFgB1CAdC11cC5UYsGf0713
FS6TcTMtsEU05RvwIoQWSF6WH8BxuvIur0WxRvG/vfa4NrL53r3oTt439vDrfWU7v0GAovKMO3gI
E1xSNYI/lijj8uJmf6mRueHaWM5JUv+Rm/Iv+wgtyCstwHJNZRQd2XFnChatBWM0SssaiHZ/WPEA
AXUXVEAtXMwCUIeGR2hBjlgpgQexXUjuoATLQSjUgaqdY+cU6AlbbDV/2B/+e3yOovVVNgzzl4OP
firpK93E78m5GmlkQq1JQ+d6R/OVfeWcCN6WVW0Go/1hAagp414mHS7BLijJBj3m0mbvm97gbev9
g3OFGBXCH+RKTaIWJ+te6COpetbDbd54YeBM2PHVVdzbzsgS6IDaJ3KYYOVVi0R3+GNfNHXkyRER
511RYaijLy5MXUY2RLrpE1JU1c8Vig1jQHJ3EtxfJRpaiBAxjB7t47l5QftWxNtyPBOWI8iAul9m
NeAQCr/CAZV56VdqYC5PugzpfUforDb1Dref6kZZhbjXbR7gWU/32Zm8MXGwifXSKVfaqIVsG18S
j+LQxBx+dvgzvGOzKC8r45hf51v0tzh/9nx/fmiEDjRKw3WtuKQH0tTKJB/I68ZNFhxXdPh248yr
p8EVPBT9U5Q0NBIVMIJR5znxxjngzc1y8XbmfA70K12Ru0DdjTYbI9BISaLL8DHDen6YW4BOfBAB
EpTQzGQsHu8R/dFvaaq4dx+snFYw+jIpXb111hbuFmDjiOg8F1qw/wElLQRhp5YZpnvNwuaS2KNL
EzJfb0QUWSWdNvfq9HJI5rAdzw0SfUOCRL4NunptoguK7bbZzO9QWJGCZbNqYBPjmYXKlwHdcPW4
WhaWmJ5kBPsLs/CGVCURynYmZG72dWQnHAnnCrTumIRjexU24SyJVHYUCj741fBppEIbhaEj9UEM
rCWkiigIZOTOJ4tdAOi/6Ta+5UZmMaQe/Roeb7cvoCtOvN1XnKsusKnKK8YG//QJAfvs1mphbPQi
ExULfgu1C1EAoH7ijHd2mbKOMIPmBNM3jQJk2QiLnaPxA3609UL/Bwkb45zKGbn4vXj90R/JNo5y
ZcEDPJ/9wulY3WP2awL61QQDt3/dEW9lwN7rN2FvTECFTSdeDUiU8xOJn3UKNWF7YIvGHQIUiDrZ
YVtj+ycNupLpHEZvd6KKYYlJTsX7pyDPQOxQ0u/7nwDaPTkCYkZa5AweoToCFhnxx+Tf5UR21HXF
oKhJLiMUlRnHFBTmwEXuavOEHNnvag7XTdR/YCWexGsZcc2uJ6PCIWUJJD9D9yS5RuELiL0ikku3
8L2LMTrsbfCuaiJNH2qPYdQSKLwgehtK7mOY1h+aNOk6u8LByZ3xVci4MSvXEPdsTKB9Hc3o5iXe
mVqX2sp4meWc2h3LSahjQVY9tWsGgKNIvtQlXsw/MTgS4ZrT0t7KWU1rm/KUCd9TUN2bkVrED1i4
520iTp0UpcfEGIcTt2DwJGjc8W6VAyDZNuu+SYgwzyBk5nBIXgT8S2HW3/zjF6lc0q4zS3GFBnmE
5LeJ9YyCwo2KBCqFsUHGT1wTpJGG9uP7NJpKzj7CZi7gbwb6RyPCfxSbX+tCG4t8IBpRiRMADefQ
2nIzH6opVc1qlCyhvfd95pGzi2p3d+1K+arLNRph6ftYjKxHZcxG66F3kso1jKaN0rloWF0iHzFw
2VP/3cVaGRP+0E6AvZiRvxZOwrl/8A2v2eLq9v1VyQfkVIBXm3SucMviJfGPNcTw42iSGhwkwTtD
zarqYNe4u8VT9QOJ3ITchny6woqKyVgUyK68h/Y+eGj1Jiii2viYr4uIXgcK6Nk7RXBgdSGuVFFU
jju0+U2B9Z0GymQ5VbQD/x3Bcki30Ewrtk8FqXGK5Zrsn9EKv4lOTl27ITUXSJKrifJNTIlbE71v
po34PqE7EqbtblSh9q9G/+XFKUz/N02hqdUpA74w2KTStai2nl73PGliHvauTZKUnrKWMcCRsOFz
LwZidj4Qkr9MwoDASoj51tZUe4TcOxtUy46Z/yBFH1TcwCc6nyQeT1AAUp84Uw7USxHSR+e/40Dd
TZFsQzBh1yhEnKX0T6ig37Aj3NsRnMnrNa7dPpmHk8yaGY+W65omsYZ51VP/aJ3WQ9qnaAUUH4n7
hT6qEfD7pEF9X0VHgMLGHIeYB5MzgJAwGVfXktVMGWxdOMOdKsswvjcLpKFRP2t1JEqnrDzaJECI
sSxz900z9OVWjNGNgIQdc649SAIAkyV6D03ldvk+ppdewhFTx4mMFkhIY9igFYQnN/SyloV4YQRr
Wk9A0h0LqxgI0gVKroc6cUGCxUiSunit5j1ce9gK/LQiO8nLHODHCgt0a2bSzf6jyrh1HqUXMhPz
2P6nu+SGv413S8SwQAOMd6Sn9K94volrgBo+2hBsk+pxZ2yVFZdcgM0rlbNAfHNkFtudzma7KEMu
1as1I6vZ80zVHHhqrnNE3j/rn1/YjiGl8NX9O7HZk5VTQo7xO9Dbh/Y61IIa5jATVH7CM97gPK9t
YWKZRR5P22DfKT+s5Ma5/uuNTNw/mjfXpWOs6q8FFcyY7RYTOtD6Yvxr9u2DL9/VrLIbJxL1h2lS
cUt+ZziZnOOxYt21FWuexJiiWqrog1WPZ00pkMiDPFexytUBZZ/cJd3XO5RGKCVJtc0B1AkliiIW
ZvAJN5gZCfUjoxtLthIsId2kG3B8BS88zH9M6UeOjeMvqqRuwKJoB5F/TFtTj0gFwUHqlFOae8qd
1abpazJ10tipTx2eEXw2TxRNX7gYplSPBu/kB0VVumtH5iXiU0OQ7cVF/rFNO4/eVc7cn5jhW53H
6ZS6ExHFbrR1Kd3wbz7VTpDObeszNUJnvgY8qpCPaa2UyG+m9WMiHc0vIAnxIaNVIcs2oX6y9bet
C9lYcUYErq7/1HBkpbA39F2U4soZMZakKwDadpVECqPCJgblQvzY1i8uy76UlYJIls8/EFh+bG71
u/AvgjDatMVpBD2eKwBzirbp+k0YF9Jxx2Uuj2P/N4eLhylbfhQAsExoCFe60O6cGyMAdrpV7tJe
lM51BNOX14Vy/Jd5F76ma9khYN2aO6xJ61dt70XLqMzqMjAwGCJf6esKwtl4pVQdfAgrVkDFlTmx
uQ0e/6fYEBL+45zjVbLK1plvBvXnC7g5nBZX9+On3QCVdUQgw9f/F+OMR7jPzyaw4Z4AA8QrruLb
6+Sc0+1Q11uI4skovjKNeydqUb9BPAJ+YwYqHiFJdu9+QQn5Tw6ioMK7au2ovfcc2KAbUDTqK37r
WVzabNOOA12FSnmeibqSy08PPobqjvR+LsLRFQOvgGOVgAVGS2eHJUg2HXXKpmy+nvvHXJIb03uQ
QAmdZrAASMCWlysFKHFqi+W1gTArBAIKdjz5EbW1Az2oVwiazC3p+pAQYXiw+V49YLQUYJqMqkVM
LLbKA0plJFs0yZKwv9o8Gi7hEP5wHLpshearS+HP3XNwHrLB1toIeEmO1V5bi2/nihHqwU1Q4Qrf
ApQq2UfnCG8GjZcjuEZ82ENE84GBVbXYEKIaMN7eDnzBfx5YEOXQGxsHhIrBAheeYyu2cJ1qtAmG
/9lE9LykLwEBb9oe2dLhix6daORgoJLk5ug+QxMrcC7UjnDAwmeP2gixFWLEzAuMv8nvFbehj5B5
N4f+BrtXpzESyULudbjCMvaTE+CsoTmcrSXS0SlAJ/cLleHQXkLKfijzOPmUIYxf36h4uAGm7pvc
wFkdWZxdUxNbnJeZKs+OH7TNCjCeaf+viGxZ2Kz92vgl5ZGN1iKO5lmG7kzEhFs04d/1wtz7unW8
JV6wIHRrqVOyMGO7YTT6q07NMfxK9jlW4cClHM+ZBdGrPnK0oqSFFhYLcaFiaDGpc0eHGpRrWiKP
k4jHYWkpNfkQUhDohjyjPt+/iPmfINHPpg27Qs6dl7SVNrP4dHwwkkD46dXOWjlQyYrTddgEXC+2
RxDpgBfE2rTgBo4CyJfIiVPbsEkBRfCNc2NYm/CBCc9JNBJjOtbuiw+Hxy6/UAjvPQMf9dLKy7ef
8Cqv+ru7G6idNRxj8jCrNnwqo9xlGLkE0yAs8eN1uzeEXrED+W1r6oKeW/eRUE4jqespLPy1t8YJ
K3EO9Uh5nd0N08GiWcG1Ut2/wJVac78cMo0026cZwkOHNfwQ0RfwMPfb9O+ILmsHASfPUq3UX0Y8
YVJq9yS9NOt4g6XSpga8TFmCvY8p7fKfA5nvwl7IZt0JB5mwL6m1sHDR2bJiYQZuBhJ2AcZz9yCD
TSInDtCqLbrUHGQOCE8bpna+saSZiO65IE9SVAmmYNePRrcbn0kwaYTdGa5WwXlEpTfYb/JVSk/M
1l4nBemjfI6dF16E5v/Vdc51CHR4r8fjbzIPUZzveLx5Yc71CQrfkVPjzBHZ8kUvIwbs+UhLJ8gy
eHzW9FsuLumKRSyL7wuQGzEQ0HHNX/Onk8o2Qrz1HUrHo3Wi2bzQy+nQy8uNLZfGxoOwHPDcXuSm
m7gk9VvnnN6MfglLWLE9Q1l6F6EkgX2ZzkUQ11CEHG6i++qFED/8S/8tx2P9oIiUS+PXPGho0Cli
Gp5+/Qm4b/EphEM3FLU53aIFuje/bfdAwp8O8ZRflsfWpsWtbgcZWILGTrdPD06parFpMvYmai34
Jj/o6g+xqc1YpTmXuJ+ys8GTxh+aUtZAkgV0vUJai+OfC/8XjN4H6Y7m1maZ2M/KnaM6O6VTsv1E
HotVVaq9cb2tsahz2oytsGWYXIna1ajmGqh8O5MfDo0ygLnpq++iJ3Dl6Ues8xH/aGECaIyjbfLx
y3IK9TEUOkXvG+V0i+mvMsWT29TMQOz06HtYAPTncPcL8UtPjrQd1B4xCnCGSIm794sa5QfFtbH5
R3jcNIKEkEmztehybo+kGiDPzNs++FoVZfIo1y25g1kZ49FHS1HJoF9VyYHxbE3NPx+sn9nLHRwQ
CBTOjAOihCRAX4LxMvk+YAASC9Ysj4r1UTXjrBGCyrdaLpCEVltQObDa8MKVU8dLH3HMmMP7LzjD
lD/Og2a0UMut7EQq2/WOLSUC39nx2e/lTYwBmbghq7uZJuQBL0i4R9SXhiONBdL4FuyCjl4IPyGG
iEDZfPAVxtp7GiTRrz5FK7oQRXJV3BFJNQDC5DvofjBuHO03o/hnO5lAom50cNxXMCugSp1Yj2RT
JKMFCJhS0ZiuLo7vPurmx+pxLgi/EqZew36Do+uVTZL2C3caxJqKNDHVDhjbiVqpLVHHXR+e8OoE
YoyrkrXkdVxxDgpzVTIbZ2k3F6aEKHvd60KYZT9td/2UrpTEQOBs0SX8zBfQ60ptwbQgwFK+9Pz1
Oroxy2pDNFNXwivMoObtGzLweJxmPuipVL6Yppvc32pBbbgdNSxAj+uHzTG69eW03N1Xr5IZJa/4
NeGt7kz4tIssj2UQrY9ki1i5Opbr+fnltqK6i+/KsPoC44D2HIkJI+RZrZZFrCD33eC4MeRLMwWv
vDihrmydkspei0YOIGv8/u/uOmjSevFfPCrDFGS+K3WzoxBft/0yXOM+g1zkqQb/NTPBSqVo4jWG
PXpuYcZgq89Ig1BwNC/nTZV56OTf7VDXZjbv9ljxjd3kaWMstpxx7kjD3cUvDQGH36C4CS6HUe+n
haEdAvxVUtGziotj7JyP9auNNN2FpGIqzCMyXr2WTaVcLPxSZ2SS4zxifUvqb4cZtF+nmr1Jjsh+
BwVN1/6ZL9t0hvmNQAKLzBjOm4+mQVg7okXEEmGofm7PNtRJxKGPxacjpM1yysPmyd0Mx5AKBRSf
7wYGMDnj/4hvynmNlXyB+Xw+IFCn1uG4DSmcCGvekaQVynSZg1+XoZjmhsx+Ok/MQPnMVzuGLG1R
EkmT7xqGWQ5R9RPCWkAqf9tBbEpqXNyhU9AsDc9uhJ1TUOi4GxScbRZtqSZ64PqT4n5RhxS0tLlE
hUh4amfcxrzXKvH+7PowIXn2vjaWKUIX6pqv0crdjBLN+BanZ6zQ8Ajs7XhetLO4PNqcHNXrM4sG
CFYbWmMbrK/z0DXMMm+oy8zJIVrhMInKsjHVAikOFDPnGFUJSCpACLFPG6y3IoHvJXRF3PiZKmYm
93CJJCkTbmtzaTG9phBafa0tgYrbNUsWne3QRXBwcgpjrb6ZMY/okTq1j0xBT5Txcf9LPXa36Jrm
xpanSvb2bfMcKVFv50cJmyal7oykB/yafKZ4AvKOHa5QnkobxX/16uxBnU4TSfawilEwlnTDcuYo
Zt7lpOA9uRhLHRryJdNyoPokxXu7pFtC5oBI8G6IlDp0K9TPYLgltGrWwoJnwLi7eraZkRt+qBGL
2Rbw8dbWyuOfWZPREtrDKXIv1Id+CMKRhIyPWzmI0Y0adchrG4N6Cd1YsaviGMHFmpq6/2g1pRQN
FM4KQXv1THTndSiLB6xUM43ygd/ccws4uARNLmcEcJL1wTnFTgvdgiMXToX1vUVqhmFuAANZ6kXl
WtrtqyeZqsz0KuAS6DxVcQg0bjQRnrjIKsO4kklXzcQogXhztTiJVZgiY6rWNyPTWIdUZMa5N20w
bIqQrLq2EbJpFDpDmpm4BPkg9/tHy/B6H/h1Yr8QdaGu5S4aA5q2CRhDE0Dv+Z73zm2w9BRKSMb8
xxLc8Ecwrpn1pT2EkPysY/7FFLdTBT/u0st/yvEWY4pyhb8MXYHohi2rp6Wjo9pxR5OkMI3EMGJq
kLYVkKcrL/0vs4kIBffNR2f53/+ksYGWFks3y6timZ1MtyutiGAJqHb3aRjZ2N0n/kr/a+sdvm66
dGmWooDAfJFvOI3SU4EBpK7+Njn3KJrJQ4n2vV6E5rDv+kdOZ7dU05cq7pO1Xr9ShnX2ZXU6HOAH
WMCltIrd8aFeqsjtsYcWo68SNUvfKwrZztYGmw9fOtsDZunoJZytuRn6n/7vt8QiO+xelqO7kFXr
u4nOQoXYXykEmrkLq8GHAU4sIy5RF1DkPsaifxKS8sluEtLs9d+ID+tN85W8k0cWWhtXyTf5VuaA
c7ReANRTnY4cFBHh1UyXb0vTiUwVy9WL3uCexwM8LqmLx+R1H2pEFebiMRDVe4WxRU1BCvblUdw+
mfYxA+lpYEWsjldodbMOdAQHghyq4K9WneHwTANzv1efufXI/kzTWN0fDZsxSMpNjT7l/upkubTZ
0XbRgvL7tpJglW8+gKM8/uQOsUWvyW145tT5JtUhnWl2RAaNIqj57RLLjujv0U8L6XzSrdN/pn9M
ljjzSwvJtFjWSdWUhdduVFbU79SoJNrwtZ/1UlOB25NWJumQaHx2STtIb9sEShl//spKBIHEp1JE
IvlcWkomAoKHDsC/9EGdhQ5OnNfooZlNxr1o3XvpVgobpPBSJrzrSIv4UKp2rWfbC6I1CY3Xv52+
KFhVjEcO4f/Vwfm8YVdCnt9K8Ib2tjqJjYVJEWnoTM1y7Wol3h/SbeofrEQ0DthQIuZtJChBlQdj
vBFvxjW/9xxLW4d1xEFLN2c/MwvK/QxZlI0GC/0SJBNO4EcFSmYYg7LXS1uLmootjBjoZ/OcNnf3
32nkxtoI1JiiXLx2uobAmcDtu9WDs2lKnF3xyyIjGGYL6tqi7L6cjPfl9sMouM7cQ303FSYQ4l3u
Pu7ITquWBm+dPuvB4nA69Vyz/AtMxnkxcWTWy7+PEcRBLKi5+cdvstREiQZz9NOm/VfdsCexYwzB
iINyGuE4sIEy+UUcNu7ajJXb1VmGXfJErmthrkWoQdH9eJOa9mPA4IB2qYKRmaCaFSJfliSQhOdW
5Yrkq3spEA7kocYbaZFETh+KvuI36AH6moxdyA7x2ktIYX5tjfpR5/DU5k27Vgw2nrxVb3GyT6PY
PNFdNVWncY2PE/rlgQMkyzNhhEj3MbZYs8flxJBUj2hiE9UzjErWEe2wZEeYB2ZrnP34bQrUxx6I
l9Sl563sIXWv2lzA627wTZD+HtdtOCVz5WShc7bREUXs5h9RITvMVg6+SZqbpjiGgDMYtpj/LUeg
FUQbO2hgCZe3Le6w1yKcyXg+4DmkfzOT8vdwqfnxVVOHzpHHXujrrY9Ty2eEELSn/Hntht7DwNLE
9Ql47hzQPtFFchTvSdRGkufM+6aGk8/N5PmuPBHsJT7RUd/4387uTdrGmbgvZhM0tgCvBJwgoCnC
BbOy7AZtqPvtVYmw2GHzCKOHLKp/zLMB6LmhRMVi60OE679UzGadktd1/oGtRoi76Q8vvHrJMrg2
tS+ohPyB36sZ97fH3+ShFNX6vg5+QPR0d0PxoezWt2PHx4mTAIzVU0tDfiNo4YxgOpWiVTI6dxfR
6MLzIlNObkSgmV24rrTIbFgJLEOJyYcaCbS8ZnxStbwyoBxb1voRr1RBTKCA62ZHHAW2RF8Me/RC
qNgaS54G2EQMV53Rt2v+W/34mQmzKmtbrHqNxz+hgRtTAyNlstOnMUx2oZ1cxNPosD5k/PL7qGHZ
kHlpwuj57Yr4amY3hhMKeJ6dyDOIlKjbfDPSaIpFV2PfwtnvyXfE/ljVV4YuPaKJvyr0FAh0Yes4
cfiYpcgaC2rBs620N6ryTwYdU+rm3Nb5qg6cgJHG/ddn2wbkqXOCn38U3For+R8pPDRkMcABM9cA
zdiGGsvykS8dXkqS1lV2BaYcqVp2D/mWl0XIxfZKLn4Al+fI+9GG3lgcTS+sWQ+uk4sa6OYhdpY7
LnWCWL+6MnTr1V0n7ycakLqAk0yRQ8p2+P3oVS6owkQYt5bfytQza9VGl3KnLD+PnEYnKM9dwf6n
zY09dZPETcSTKMgKN5Tzeg/6gsOzOPKBdY6SUwL597Z1dKdZ+BYCRLNmDoamHcVGQiUuEAfRC/Xl
iZZRDkCBu2EmmjdbF7W2E7pePHXsXqXjIq2wbvHKjzTILlJb39g3l17uFgiJxzXEmej57Z2zUs6F
PJ6QXO8indIA5/TbsEAqj8t9TnlFLA6rfay0ZEG6ZJaeRK+JOD057/BVfFpPnrbo7AFZ6X/Nlu+q
BC0V+/T0CbeGAvcIuGXy7zkm0ZQp/whVA4/3JfO5i+8xp2rAK8N0HGIgI3Y4WzG8GhooG4ahbtKx
Eu15tO+ERBMWWQOLbWOkZuziXZJ8dpUPVgZE8Evd5Qnet9nPoqwjgyTkM8tjtSnkrAjT9JvwLBFs
LgBhcMugyE6piN8ZGpbZYpjNDrlI1nIqhxVohMNZeOoAOznnoHmkk7Mz0zfxOENtZNNIrn1kcDBT
+r73i6yzuPOxxs2bDMHrXu8w/AGyZn0lQFHNuzBOHS5UhIptQxB67ObOsyKwMQUNQ97kaVinWR75
9Pl4WRNH+arfEtqDO3QCO7T8lvZ4mrB9/jfPqhXjtp5PKVqgz5PhaRAc6mG9rgiAe83FE/CS7jn3
IB650AxDCwFQ3imtIRv+vfvxAheFMT3mZYQL+IU5nAsl3l4r0HQHTiKhbt8rgCHAYEOP1BjgyjME
okUyLYqdtQaQWFYD1KUXzxRK4dxtfWM8I0bi/0uHfjP10AK6j2LLMZHD5+yuZ7tkx5kQhWKS2R7V
SHdqfgyvIyEUvEIzsJzLobM6cflu026rsLz3/0t23Gor/dYC6EJJNzcWUtCY1nWMyOnInvsjd0vO
XQ1q6TGqTbT2jNM3OCTpiU8IAtm3gag0bv7v3Rx6Dxq0IoZTe+10mwIjXrfQ+b/qSNl6nrYO2Vlq
ZI0ZeHjtKl37WJ5hfS7UYHAUqh6zm6KYnDY84VlRjnrnPn4mZeu6vFwM3pajEnZF1IQ/Z9UEgjAQ
mbOr+nCP68X38Mn4AO96kE9vrot6nZixXm6HD77yjE5pu0X7B6hxJoayCamrfxI10h4ZVBSqIEx8
jzwJHWCRw8lyMVZaLe/pzMGjYzGvewJ4+gl1dDHIWlLTtU/pwrThwlwpR9hLvNNXSswJvWkbDRCc
LNEJQAk4NOL3LFv3f5aDm4xlrcbdZfREiDcTxHFd4/Rjs5waQdVDoW0pohOlnGy4qGmbNI4GEL0k
ISPdV4UCL+801kTWaSoDHp4xJz91BcJT6iZTyMIwYt5jPAxx3YcZnK0pmP7UNSx9Sgt5VZmH3xds
WT2quwG2KTyAWXMqOVM2CTet6oPn8sOTtoC7pmlnCqSm3xRhrEpPNm9QDXpiLX/93UXZ2H7vfnuc
87wT4RVVgLGfrlenHMSK3En9bqvhn2YVlaqiA4HFmpRDJ5gFVVlEM3S7x1RQfCpDONBxURNaTvU2
J8lrzNzIH/EML2e7LzeLZi0hJGRapsPZYGbYbysO0qJhHdVFxylUfOYu6+vG+y7a+pR489KgWL6C
fxt2whWT0OZdnuqIkSVrVRb85+L4duky2BkPdBs+WMCze3Xt7Bau3frGVM7YJd+DM2+5p6XwURuC
s8Iz9wC1L5tXef8KJ+/SqBL9Yg461fnbLk0IxtWhGmYaNi8Tamn4v4KHQOB/dCk8amcsRGiNCQOm
D14OMc57YMJZypW5EmlEyvlRj+f19UoGbZyxIE32xmObOIrTFgOgllw8g4kkCn2lgxEcKhKFOgid
yPCv4FPvyLxL+ME5g0BrmJ4LrAPsiTQPtYE0VQcBbp4UZWnWDgXC86rADBIoqeJmt7TcMuDMqGtk
A3X5z1wU7EXL8d5argYxNsjuy5XRKGrIznk25EeZY4Q5dXpIUfubox/Jb+YnJnJNX8KGnFRaP4CJ
7GVjHzJ4FJ+QKkcsq+x7Me+iJZhFKJSpVpsEwvQajr+19BfisfhKG9QZt1R+DfIWNcHSLEBa2JAr
6UKS15E97hXo60LEr24aaX4Ti1N8jT4CGTDhapivN1yCwDnriJjo17Nt/NOwZMzVIrRM2c9x3l7+
8x+N0PudNNdgBRLr8rHjST0phMoIy5M3iwBhrhT5tu/QlfUQyxp8O1XNh6g1aw2Nh94rJS2vIEWd
xy9zJZSxutYe2X29URXup5ogSbAwPhQXQGGqXS5C2ANtGsUaunuXBjVRhocR8rNwYFhLqITJJHfl
JyfnweUDROsq0nZFFyebVYxru0KowWjoQuuJ70c5N1AwuNfX34NSJAYRGDBqIHMJomPnB/UJDxZV
wC94b829vHisXcQHki9ldsI11/CFaJ5OuFBR4doFc5NGShbuIKyXXOXk8Fo9A2JlDUbcHClTlQoD
yq6TPV/dOD5CYfEFLQBRl6NsIQzDs7bkjiIcCCZWmfgfF/t3KXpAWABUhW9aLP0Rkx7g0Fxb2Aa1
ZP+nQYzvLuM8lnqEwQoZqFoRSgWpw8wW2hWS41uCxEadyo4IqEaxWVzzWq5AWrIDpSzq9PD7wSUV
pkVtvb5uul5mAkA4Hu47FGADk8Eqy2rvH8qXiaUDs26HJ3qj/whYk+a299hpwayeUkcpXOlVbe1f
FQg45Od/QKy90pB4R/XSL7UGgS75LxfOxHczALgO1+ZazBpYF3mvclYjFqRKoR2mhDMEP0GyrA0+
QCxDyBQ7PnkJgXflTsJzpufaHhTyU29VsXQtSTitS58OtNYjP3Kw02BHsPW9ktpAlP4H16namx5T
Gf0mtMnvE+xsyVVJOwTeO+1SR2cV4NHc8j7LbK7Y1Ajk1Wqsb37my+mLAjoehzNTVyS20gDjoxEw
TuNXKffjqGDlDpqaxVxyVmohJwbCb4ZqlfLVzDlGK8uw6xB/eboTt7lpHTv6RJCB0aeqNQnTQ883
LbFuhj2Mk+aJ0uh2xuuqCAhx8nEDzrRwnXMQ+3vOaRo+9Ppc+yXyk46/uAHmZQBYWssjwOA0J42O
5XIpBBXgse/55CtmzcUDUuKt6GJFoyVpo+I9NxXcS6qEoU6GPha0QEuQXQ5CNKXmA6j87b/vTiBi
dWch9gW0+UbsPIJJRubsDr1foo/TKnAgzNTZ6g6bDrRkAVTmgXfn54zfAz7fPf/RfahCOx6iYF5k
68yJldBEeAQCYg1xXYgruYJm0ivOoUsF9lQBY7feMHBpmC5GgV2U6madT74Ub+ejqCVDTcZtYr2m
tyvXgaYWQnoNYEdXkSso3sEJsKCAz0HW4kLGYOsK+v74xNLFheEjKM6o/1WriBGvpw5w0lvDZxhk
p/i0p1/QGTKRH2QLCz5Nby6yT3j5dT9uxyM7sfgsuDPVP4O1C8MseeBQ/yJA7k9uK2l6eFVSGOsx
deiqFWLdFBb/D0xMKzIBxRNL5oWxQAEEMC5AYeAbX/cTz1WU7eJPjvxbD8gOoq8TqaX1qBrgI8pk
IaoaTyIlMiP5nOybsSGlKur3OoeishPtzyiWRD1C50lShw0Jatm11nplqSiJEJEwdJgZmcam5qIS
rvVhimkMZyZ2oaBn5c5+g5dcWo3uhh6Hz6zxTJRdhHy+sS1aeAH1j5J4ibymHIUfWAMLPBkzUUjD
O2F83cGoOkgezbLRoTz6u4aehaAf51mdAru4O9h6XtH5aMn/H8jfLsxNN1643hvEsNDTmKd/CppH
URoJ9cK/kwuE7t2bAqRlyTBTm41MzSVE8KacNPvfAEjG/0p3wWXyzO0fk4gZbShcRKM8ISGrH7I/
vm6Ee+tR/5RY7hehfwe16nvrgaSPQI6oHBuQKvD0xtOguYtNQLKtDE7YvZ0ZhA5vWjMKidIdUdST
67IDcrdBS1RM5medcNIPt27RVDKYB3+6mROdYiLdhq2Y4vPaydmvxfHD+DTSWTWMHa7IEDtAcf+3
av8OsBuoiS1v2RND26Fs7TXA3qRf986aRU4ZZ3TjTMZKK6YDbcsLt+GDuPhvLLDsy1+Uu1ov9bgZ
oJphA+nPaEup359uN5wjeK+UfIB6EXND1rar87vMraplEK2yCTCIDBz+lXMt5J5N3aLfczn5dQpu
esaFVfNhrCzPjLv9ImHQA7/t+8z5Fpirk6m/c5+tsgILoebO0mLh7NrxczcHeYRSZMKKkd3gJ6WS
zJl82Bmh0rbUbH/avJK3ONgc9rax+SXalgvqEVOIUyrnxzm98ixjXP9fukXeIdp5aqsljmyJGb7M
xSVm05byO11rbuNobtWhSNKTRiDz1WIGZTXWuqoharJAQ49XxOsF6bB/Gj4JzNl2WNlMvearhp38
9QqdKv1gDo/YGgvrZn35e9bmDmalc17Ynhves4ZFXgsEGLrF4aRIdlEJJtMhlaAPGiHBZf6mEbw6
rEAQFKb2ZvH9qHcx+n2D+UIJMqWxDFMBJOrpW358ip03n1XQyOczD9rYE+vMuxHjd4Bw5FAfQLab
s8XaW6DwzVa++XHHM/sA+4h8ZV8C/69pFaSFaefabxbh+sGJtm6gzCuDSedblHjoJCf8XkQBLHQe
PdIS5UPEbmJStBt1uWxZBFfYAXH80i6ITLJ/g2REUNnZcGN+9XOJE9Qu6PEuL39hCt27pEJnEdIc
4Pfx8iRmajvg/oZpJcsaxdO2vZCAP5l9iNBXAcmMcJh8cyLs6Z5Z6wGB3YogI7EWyCmswNz43ckC
Rm/OZeFk0xk7UorFFA/g2q71pjTqEk4VOhC+/dBMZnSO1oJTanacz36PBywOkfQIL8wZ4Nvabi8O
2tWanzOzD96+Is3s2y1gSGHVvz6A9wsST40Zsf8L5+qhOcHZ4pjEVpdxcRc94SClrOdTwSr00FRk
Lb4miYPpWUAeKXrTmc3iASOFvBBOo83hlUxmskpQvX2e7NozxLid2R3lOTE542KJnLoXZz1ejTQ8
tsMS8Ew/FHLLG4OiO02S8Jius/U+ARsf1UEa0RXOkONciiJrd+itgm6zMNnTHxeVF2mXZjNJqZ8w
Qq+psp4dvn39lfFn9tnr6r/Ubp+weAczRgHVZ71t3WyPIFi4MslZWZWJDUqr3KEuAEjELixnRxV4
eDf1Lu8AYtBNsZhD6bHvnEdRdwcqwQ9blqUNe21s7tsTIgqY8240piM9IRVtLmivErixnesA6+C8
UnD/qDpjPhMeebOD8/1/2EJ/B67rq1pvH9mQr3gZVjuSNpbLrcgYFaYFQJIFCqoJwXWo9Sie4dbs
Xw2yKninzTD4wfYaML6kSbhg1dVsiMcuZgTbNe5piYNWDsSdFF37KTpq7a2Oa/xfYTQ/OUouKYpU
mk4owE6XlgZ6OJDbd0G0TlQmr1jkhsLzigyAFOyEufubl4ysYuNsu1NLdOxfmrP2x9n4iednxbLK
DGv1uOffYIs9XZiIphhG6//xmFn1bhfN8cvPGIBVE7WIdbEiOGJdcrj2GkKJAVPQXKvtJf6K/DIQ
oGFEBPGbVzCV1OPEPBQbAdkTZTJ61xUf1dgLwfQedBoCkNt1d/aGrOBJi5MIeWjHlpD1E2498DP2
SMIgnvDlSxnCIcGBXSKIwjeVzyRfZKldMElxUwsWyKFG7NnkZRI838fH8sPxE2hL7axGQPyqxAde
rmHIteu176kuAcyUfOE4Pt8uZSsWcXNH6jad/wfXVVptSJSGhlNSyBLrHSMFfDsfE/a89ct+SO8S
6AnxeWozzVHzs70n+1nDYrzxkDLKWVXr4oKUIFxJ4eHo4trry0HS8WejFzzftWW6VkViHJ8XZKKZ
/hxrYOQtS1FYICK+9Ap/6e8+uSpxQmPjBjY1Kcg2Q7v4TTDH+8G8Bgx3Us4Ch3okEzI63SRtc6BQ
gY4tkC7Fe6fuNqUPuDzs+ZNXo2LZ+ojtqwIb3u7A/TlbGgeYHBPZArc3BD4/ZI1H0dBxT6V4m6l2
voWoKo7+B9Dokxl03qi7V3wyh0+7Zz9N9ukO5JpcorXjH7eY1aFJMVtVkJq3CUENqrNctayaSlbC
bJv27on6PjJL9xfvILRP+kbDf1e4AWUNpicl8WmCjD32fwAsagNcJvmc6tmy5C5eMEv7lGTyy+nU
sU1yAmLrYwZT69DMzw9NR5XpROhNAds+jwyI8S1Eav7qE8zpk6nZOA6Yw2ZtO9N8cfLEVVbkUKNK
CWLT+6JK8qB4rO4UEwFYTURh/MF75x7tnMs8/HlC7cG9RNc9hsdevC3ilhfzpfvA1Dn89SAOsrwJ
lc7aRmr/8J6IAwdjouwnXzJt6T1azVVZHEA5/6e5+0ZXYE88uLwJ6mWJUkflRLva/tkLggcSP+uJ
ntTkQINmqhPyqO3LORKHw+rHBNYOfBG830yHpohR7xWOxsQ3XW8nVaasQHJIrntS3i9oJsyY3PoP
26//Umaso0/GEcdVR2x4D8eQ/AE8OTQfCfq1Mi/2MgmLEPb5JKXtoPB7wxC/vLWb76yu2iYU7d2a
2enmWUrh40TVDcB6sJD1cSponoKSuiyRUdb6lpHBZD1R4nznug4reaA5wMvtvQv6wyX6yEIb350K
wZ5jXmT34RpceSnozKf8ATpQD4kN/dKwxOFBEjzUN0mxY6wirFCr4+6BdNckPisUCxZ+wmwWblri
dEuH2LcrT7iaHzcn5En0rdsellpkBPmadymZivLN95uDuUIEoOaklwPOyaBbDiiKgjqSLxhUyZ7o
AcPMOZWCt7BKTA3NLt986Yvwh8OHB2ysxLZmvlWK3KZVZS7nJTrfGXljwJ4Gem5StHRTHdw7gPLx
bS5UD9OoQ8vmpUkvFgGb7QJ/NQZHSz1B/fC83yU5uOdQO+QVAKx/V1W/f/Gr0yKS8slWUKTgJkim
nWV6B0SHKtPt/8I3u8aulMuKaIqnkNeoSTMR+abZM4d1EmAFxDeDgWhcZHRGm7KYkgNBaDwD+a9t
/HEJZSjWaBz/xzM7QofMefyMyPDw4FlijwKlv26plMm02+ue3/wyWs8wvqAzkuoIDua41YutkDqe
jr6VFqep/0iU4nafCPEG2ohKhpXRSL2RilLOdl6jAaVZBhrUvbwMIV3FYM/eupEn0gInZ2WBEjKs
LUsBoMSxCWjIRSPBFOgt3nSJrzKlrLlNKvSMLhEuNMMhX+BfgVqYP1weAzyf5IHo5Zi1mPiOc3g4
Q120n3Q31dxDGAqSI8Krii7p8eZIjVccNdhvFGA2569H0MvNaMdxvPH7WhsfBw1mCUsEa7Hp1S37
dfPED/YXQ+FKN6aWesQkIbJ12NprvWi3rmC6oxUpXSIDgSpo+0ZFEJ4j+wJfw50lkyENjeGDGOHz
fo2Yjex+sJkMER+qGBhpJ5Pd2kzLGRqX3xob3hKi1uCqy6p0WGsh3wqg7rFOLP8LB+4FgzBfE8uQ
HGnjXr4IxlbnA5N64fRJBClrKYQNEvWH8UAeBU2ZlBOjyz6xWG5a1FDGpb8ofiZxdzuxLr3MaLLo
csTBqeGje7UKMWeMug4rmVeYOnVwfqIceuh3YWHV6etQc06rtmn7EFmU0SUFMJxMakmIMfFVZn8Y
EH2kWx0+Oju4pAvcxFeY4BVwCnvHht6aoZtg2vEAAqiKb/BqlvNErdZVK8w+ImU1rrxKDsq1uZcT
/qIn0o5gN4RpKRf/KRMdriG+moQeQX535ZtNg0XPKxaeE/ObC50Wr23rStOEgl5gu6taCTuS84mj
+ASGiyFn2z0Ygv8bPpcvOgCEwt2OklhmJQIV+8jpbaim2hxfTXk41zr8DOobFYdUZUbnaQf5D9Ut
8w4EHaj3uuzuK8AE1VKZfwxSmwldsTMIrQMfVvizCz0M17S869I860sLIpPo7n3DXE3+Z5hBHboq
cF7v6ufHZCKGDk9qZaqWPRyqH9NZeCoAPBgdt6UmDSJdAFU/ThoFT8D5HmSN3vtmF18jF/KLpxhX
x+da/8Q182n4oMrB98aP9p/rPuSlRW23QwZyrRzV6nXsuC/dtKukjQgv4FEoS/aEld7rGMzl1bKy
a8ZaD+kayA33rnuchBRlAnZxR0jFJkcwaFA+YCvGn68clU3DMW2Z6m9gfX8Kz/ERM6Ju8pwTspUD
XIEBpx+QgQZr0q4YQcy+QGNag9xwwCjUcqDzjWlg0dSDozGCBcAUbL1G+ITYYBJPTKc3v8WuFd5r
p2KG4c+jMnq1/6dVSvBfOW6cSn/6H4Tx+Rf00jKVmJYRbLS3ZtqhSCQvKkSRVL9qY9UvOWdAFdpW
2mmskwL+k8x2TWFCwoTNoBJJw6m2m2jRMDzZrFvlSY3pTcFjQkQ0lilCGz2P6ZmqkSPVHafu+MCH
ftlx6rNNCpZPIXX9e82f2DhzsWXXglE/TrTkh0Icrbe4CmgbzJ3soWp2GdFwsPhIrNhxgo9+CRHO
8Wmslc5HJkoeVxON+NACxYYnikykpihyqqI23zxb7Bk6j0lzsyveBYofvEtLUjgz4tKwh/JvVRQZ
jat/XnYe6oBUOuW1IY3OUsekY780OGCuhsUo1Y6xSmZHbj5xD/7g6Ww1c93Qf2VsC7gMJk1VvEG4
qxQXvrQ6/Liw3b3ID5ApHvO+GHZe/aMgnL+UQpdUgT/LwwirAT0JbsPP8kw5vnYwAiMnPNPhQ2hC
UWuzMUUbvVNHL2pSIFg8RN0P8EHEH3B/mPwZLonseNDCCbrhn1GcB91ANsgBsRvsPDxStSDJ3Hhl
N3Y9QKJeabymJW0GRoVxw0rzlYzxfbpvsuPLu267c+D0epyA0WonpfRBf6ll3r36l9dReH+puyxv
utBLH21YOCVdrtvRQf+KKbTmWCGnGLLu4+sxhql5wFJP6DBDsfoou4MvqhJsGcrNupB426DvbFIN
xUPF5omTUDeCf7f+g5TWk7L8tCCGkgqZSwOYN80/w9ALwzcpMt+w8qroiA9NxuEhBdPr3WyG756X
LMy9FElrXSCMElc/F10x+DqUCamYT9z+5a5JbOye/ujRMpWCaHYmiN/NScRtEzTGcA/JktDPs1sp
Aj/JxVieBQpaXZxtq9AXCtmgIzT9gA9AwosvxX2hELQXXQGH/20N0+ehQKdTRtbmKSF9NEFIh4BV
dDARwFLjgrGy1GApZLMrWEL+kRxqHj2swl76lCe+HT9anxL2oyMAdzCObJq5Q38q1R8QFBFUCwE1
8eTebdZnMj27nFS3W6E9KxWIAcFCboRyaLlnlf8IiOT4Y8uy7pJlnh1lh4Mt9A12DHhykF7ONHDH
TUSAbDn/vAy7eJ6xhB3XCqKRyaIqm0nR+J2F0XbZjUDjpnH8y1AEHik7bUJ3fFtCfcZ4cJsmdXMs
eNk7PFJ9S0HFlZmeuU5PWSThTu2cjuK9r4R3e9XXGAmbdNMBdp/Lt/OBEEmeJg6TTQUZ+UbnGPuL
PyxXGByPHtj099iTYlkEWypya1RXEnrvKMOkZRxcbTjsdbBQ9HnXZe5cYNbmgiZCFwhC9MxTnFiZ
/BoKigt590UFYmmKhkBGZS1D82MoeK5YTduvqmS1A730UoeWjtTEpTOqaahkAzJOR74piBmwibMV
/KmSOKa4hP+S/LCBBOJXv2UEChSX5mChiYPjKF5vBqERQVmF3off7TmyQFT9Lr8Z+Lm/noS0M/4a
fbPgOhKWraSsIQIJ29qmgDLX34Q5m+M2D/8VnZLHf+Zimiq1IrN5p6nfnyqgq41l7wS7IW5JcioN
Q04RnS5Nm5MXAvGWgLotMPDzlz0wXd6F4Xj9TRDg0OGU1AY6Wwskivf0bKA2sS4GWP3faolfr41k
rYVxBZVssSfuvTR6RPdwkctVCPUOu9C5E76+DCVkEayq0wT89Iz7jfpu4nr7iWR2X0pfdyEY18Y5
Itgd0rjdSVyKHpC7URFkN4+nbK32k4n5iDWX05i4CPgugoFxkwvv3x5CT2dNsJ/r/a/SUNxdJHGU
MZvHn0xH4l44f4xBJpmjMz8pnZVOs//IyXqRmsV1hIU34QyZQAjzzDR2w1MwDAuUgOKeRdhBG3hI
bEZBNof5/G0Gv/uAUjkkQ5T7gAVeHr37ZtPAW+OiRwHCUAomiSyYYV+e8ff1NGzsYkHuGUH2kLjA
kKiY4tdlBaMuDZ6FrRbcOLe/q6lIN03Omf5Kd3utPI8pr5gQxzaXUf2VpqhQZUjEzzA9iBecHvM5
UwGeI7msP5xjBy2Hus7nG+wVUVbMbx4//IShEF34rpcUx1ugXJJ1vzX/+y2WA2tTYKtJYm+FhOhg
6NVzKobSwZGHgaKko5PQnlMe571Hm4agY/frUb6KABAXFKEHRthw+ICi5ti5gjFMTdm401/ghi+T
KwwYHwbwy3uPg0LLD4cLaEvkEFF6ueAdAv2FxDt78/+Ui6kSRK+4Fae19trqeAQicdPyFDb3kZor
tPYRZcjo1QAVFZYa88YVBgEzVKlyIhYT4Y7AaUzgnpaSwJ0tGqxPt+PhjWGpFAkq/75tQAQOJUPP
1U8hrQRdN1oIpK7PBUeZeDQ/IOXsX3pAlWJ8MXD/1TF6UlUkbhtqutTqqQWFjjo63ZIiBI6ZRBfP
mFrvzVj+3RpSf1qXDx+wuq0wPxFGkibCCQS377/iNLUKAnJ+fNwKIQKGRl66Jz+s22S4pJfB/pHP
IeEAWsbVPcmF8wqK+1ZRT+4oEDxce0+69yf1+gfP/7Nk7KKImHQkFkb/zHWo5B110fsHhY4LlF+F
meDiPsLNmT+up5gAj+QTMzP3UMh/kXxIbbkrX2mTmxcyROtjWdD6ujmaxQIcuYUntivcb9Xnf5mF
y3X+PhoCOk0+FqQ8LRTLpoOtpCsmzAb8Bb7AVkCQJx8sCn39R7MIEG8ZRnitW4AW0jU7mXF/qC9K
gOOa0fB8+SE21FkvGCsETAkJkX4FRG2y25H2Xmr19wmPMq8k0NE3VihZcUtb8/SLOsrybX2Uw8Pd
WlfL5FXTT9YlfeeuF+gEoC5CgotkT2fuSgzXfZvgGfZSyK5Te1HQEfQzeobXJc1JvRB+9bNr3CgV
hje6r1rv6iRi8DyZ1OR7/0QyRoq+BghjvEfZS/ou5fgC8sbhLFkAlVdTip89J7hN6fLhUqHNZYdv
H40vq8XHhOqzX2HAQflb0p0c22y6VebuTBVFwF1X+lWPEWatoj3340oE1xIxvl6PeIrrYN8eE1oV
8YXPzJcS9akJIg/BKF9acwlYX8tL0GTnXwXUCYG4zgW9M2lardVUBcVtiqrs8IZ6h0pKdudeXDf3
ERbj/D89dFf4GvXwUsG9xknsgPGn53QDy7x8nn1IL3qHH7tPcgVWo8VOW7+uZTGI39FxlseMVKwa
JVHj4jjIEyNbF/gMikDTv895psNyxFZSdxiNOAU9eUiTJoIgiuZuOPQtAfAipVh3eK7JkdDWIeid
Nbo29a2aN0dTfpRw7ucpB6hGbDeLJBsYwUx+FL45jPjv6AdWSJGdA6UtTLA32LFanxgpumuhxFNE
ITPPYPdxUPb2o2AxpNqXyVxagLVrSVJOA+5vO9fzv9h5o5cEn0U0xeZjrpHOtL07Msg3i87ZvM6D
u2FsmxzeT1nC/8J7YnREqpSoeJhdUk2uNHIP73bIxFVA0HB4BRIEucAmjJmkLdSv4LwCP6rg+l2H
IXd5rF27teioGoW/9CXEHzmnqot84PKw+aojjClB9DEl0isGoIclMTj01dFEHyf8uQiNxP8k986s
5jBgcdTBiSp7bMUIchfRTkw715zQHpQEZOFgpoXALA1yiH/RXC/q+xMFRnEBVFYVJuNZGWlMLA6h
7IdOd8vP8rU7YINp3bUQmzAsdMnl+Es7hchI/gH7JGnvrptLY1y49qYmLKC7t4WSQukCKjrr0KUV
hzyrmmvbqTILRWq3EY+PFbb2fEdGwzV0CCHqUKPDA9j4fTztk/iaNEckMYudO3N0BfYQ+7q/yf4u
Fs8YBdfSvZFIexEO6VFyMYcrTLR2duAlR7EZJ+QZgbzsmFJHXWUUOUjamB5JO5osgMr8Cy8jZ//F
FWB/jhjdEQIVGA1udWFejT4GO49gjyDfor6G2OozHnMhQKh1pWXaONrE/rrSJ6lE+TVsRGD5lxG6
lRZslOgWuJfhH1CehazRy/2snCgsT0JELnrZMPy+y8Yg+rPQo0IpYEF4L03t0hUcfXWHe91s1WM1
p3jiXfmP0dIeAFmzEcOXEPI019VuTzfMC3PTdULTr088bFbDqplxBuWszqpqP5W15OuvhW4hglT0
051aPaGIPaV/PhEzhPEZaAPqRK4Z8gKyoaznG7xBYLMm9bqCnh61xITQy1K/Jgl4re4jLar5mA0d
5PR0Es51AahqutxIEKEbw6m8G1zbi1DD9V4EWYbAdGVpkjczNHAWcl+vQIaoDovMueucCMfq0oD9
dptu/0Fz+AVw33wH5YXa04OH5c0M+ZPdKSDu7w8w6nouP1WfLBv3QuMWR7HXvm0+9wuKUFLd0t9v
zOMxfZuTxeool+fVxGbGlcyp8DZz9NFe9YkkH9tEUXnG15lkwm7Ftb4WmzGdk8nXnTf2A52/ttAW
nqOEllI/MsYJwIJM/nS+kM+xilB4UT+/Os1Xo8+E+pCJ1whAZVuEdMLZrMzSHpxpOHm4f6f41GVS
y1RGN86xrPxWLj6vS+r6irzGj4MefgxAaO2PjYd2eByh8TrSyUWOIkMc34f1/eRnUhSMMH5/kjWn
h7p1lzPFPYfms31r2HrpX0Z3F9fTfDc8QJmzpe1JUJyjFlrEpRU5Xh6c7mnHND2WP/PkbBdd6cNT
ft5BLiKrsY54MBeulIVt/RWGpQ0TCH3Ny6Zj9SDoHEFxRDuI8fl1E5fDfD0RqSW/t8meYaPOYiy1
N3NNBfcOL9L2UuFebb7PN7sksSuxpimqecSjAfPhPAPI1JMCKfp7DW90moTGmXmJY56ElcOLTkma
E/AeqIje3f3QdoQVOhoOzitmlEyLm5K0iKhQcht/qtWhcILqEteTzbut1nq0Wz+9jbbPifcPNHPL
7VrG4ICV/33p+tB7LoK2/bhuVGXqO1Z+Cikpa1944HAAFKV5A0GbV0zM9mkhk89Te6sYOVF/Bj75
YgyJPJY1xih/ys7URAONeKDOhYWrrqdophp/nNwVguwaioP6Sm+NW9teqENXC+Zj5k50BViWGcbq
vYX+6DBtGPAZQSMlzV4EVEyYPBNztBDZGErsKBnzdFWFYtbGHaR9iMGO+3b+sT/7zZFtrAGOfxCF
r8ZdB49pFQdkDyUzlGkOtI7ywcVTcF75eZ+0Tvqj4dwY70/P0pNoHehyTMGsDDxPO1ba0JaXahRc
wJ6rkLoaWKQhh7xqMaw09mQXELrxBnFr69/oFRFLQDB47k3zFrGpE13lQL+tTs0Jgv5yNy1lNVAi
QdgnApNoQY3G6a11BgvgQxyUJGE1fzQCTNIdR6O2LspDQFCUoMvnmPYoHK9cUDBKekXr9/S0aIfv
e/Ghx76PTnZ3L0CReRX6MuOb/j5KDFOjqXwSyFv/btW1Kht0mRrSykWUGsyqS0/W11skoLCo83QZ
XHE9NjSql7ZZyhPRFaDqPLIY2omhHvvWCEHLbg4EiySuyQtAbjdyupK3iG2UUGLAJohhpdMv0NYp
YLOC1DZFr9bzQ4fLSWYw1e4u5YBTxSxS0yyrBKFvgfiS9GYKhUqBUg99ShJ4LNmQLPIcW+8L9SjB
YPWYbUQ3xtDA29S6chOl+1F0a/g9a8pH7F2bkyLN99CHpaq0tHPp4jC12VzjwejnaH2gTtuu1vda
rD/a2SyVlQX4oYp0QzgfROi6YnXdUU5ZEBaTgJUIrnM6Lv4Sk9k3FWbVvVEGFW/Z7xDUdVYvdxGE
/V3vqQv8iEmP+UUtqdfXj/DMx1jdwQvYy/S8+heAb2uWychSXVF98hIZvamDJmmjWdR98m+8uejr
xqOXRde+5W4I6jgF2Z5/WM5RP+uneYk6WSD6vEaR2MPifpNsPOrFD6WutMcYIID3jDDjKibE02dP
mEbqrkteN1pMjlV371CFQSfxZoJpm4D19f0QCsyFTPg0pZA2Zo7S3b9a3PHPs8mdvj+vbsRc3lpW
ETyOlyw2oo/ZydXq0Xod6sXjLJNm+yatlKdlCiwOMWItPP0hv0WSczSAo6tfoHCgsO3ZSpYvrDVq
gSfq8i2zl5rQnyUMRWW1q8in7hm0WRELjJJLePm30/frk6c4TONzCNqIG/t4xuczKSOnIcuEcxvg
V730SGvblC4q0qaBr9/tZOCeNyTLnRvAb78DUnhRIU3IPGlNnDcVV23Q1YOlVKVlRp/UyK0nOMLO
sfAe4hN3gocBajk8vDTZOxjtalBfk1rHZ3sHBDDz/3P1P2jPWsOb5yPXSIQWQleZwbBD6Lsfr6tx
QQBXh50j/79qmuLpS2T2wvnBXvzj90tVehcRo21/UjsPZOUyNk/x10apJS/Hesop4NBB+1ZtZDi9
6QImNcqNG8AhAQLFzH8lVlw1TcTl61WvebkbqlA45TsuGf5TdsrGJulWGjWV9AkwcOrLLRS/bylO
dhWF14751CJ93YDou7qWWHWCc6MQaRkwPdgY8Z+e5tZUZb3GK1+da4c4uX05waN16XqLYx8RcLcy
OYSuvrbwLcdwx/qwq9sOLnuXIIHNTa/kXylFc/NzuwRI0HEEy5P9bOlT8X7ZreXeATJ4YP9ssCvS
L1M3vjJP7hOa7lG1CNNHRd5yGhjzZE1sd8NO9H4r7rrZavbAi4w6dyuPWl4T1t5b4ynlwCQyztWh
NG7HZPya9XZtm31fMAj4nVGfXTAu+yPO8USsTZx7N7Sv6mgob0/3Fve7gAv+d3nHWd41W19FEb1d
iy1cXo/BFuCAigPUv81VBQ/Ue6cGiiZn26B5r4DKFWtKwBIgAQ8ggnia4ZgQbeziy5SZOU6TPTTo
725Ql9JrpjEdeZ7IfrJ6dWjO7v4Wtf8pLCBqEwQIvTKpV/WArNb3Hid43TT/SPo0bAq11OeJifVZ
7y+WIZwu0yfY0b7F4GZqEaDwRUc1Jy6krlZ0tYtKaLAqVZSEXaKBK9nOf3GuM6TNXMv48lRUmuPg
2JAD1NM0Y/RLxXzWSOtCFdwmSwYjb99AU2yK1PrVFp8VS7vzCBfm9KiUGoI0+D0wvAVG3y8arIFK
0/OJaSdGli5QG2T+dRSqyHf3O3KC0V51c6Kttw83bH870+zpbmylS/PqIUWW+bX/TdrQqlHLUz2T
obIp61F8ffqKqYUcM9GPa3+fj6200XhqAJmo2RGHJxV/rA2buA2rnsPEmUoJBk8yWLM7HqqUHWOh
iaGaBYuLIhbI8Lq3JQjmMEEPX4dc0Dxpxi3t/6lZnKxs8YE/xJeeWmpBEPOCMrYkBToHjHd2p6Uw
TsCk5OHVSvxPVOk9skBoob0V6Rs10MH5H+S0MSJFaePe3pc0V52eC/QsFaGfeGzmqHskpShb5APg
nQMu5oKGNMR/CZBu3ma5KmJhif6WaelNCHihWjxYYhFZ9CTq3BtsPLH+JP0zMVt20l/eMreXCAE1
w4hBWHUutPUSdkeetpKUUDUnnpmddOv/tEyQvCDp2zQ8H01CYSIXjqPVETK0Z0JhAC/WcKHiPa7a
3MtC1TTiFUr2XXW+yqXzPLJ9X8lJlSyi8+adsFwaySBErzAOk584NMLmz7axYjgKojkFELpAN0je
SqyYx6Oxv0OcYVuGi+cRjZFOJ2ELPumbrfv4ssqxRLdQ2AHw0qN1yRJNaK7jUH4e3QxLHKdlg5s1
WUtCvwmPY6mykEvjpM5RprbqfQvvMD1NM8QgYDF3jggzNiFZ27/91+FzsaymR80EotypvT+0vcmn
A3J1LFdcyMUgyegHQHEKg3DnmSQY1/TRsgozepkTpKUQtkDzmzbW48wT68xGJqJniqGfURHcYoJK
Qjl+fOYrSslnDxYo07R5phEoAxq38nEhNJp1a4d5eFEVdUrgpjQ+K9+3KBrLpRiicVBKGpM4LsWb
s7Cbqtlx4ecnjWRaCfYthm6E4jmbrdXURFL3rH9g3Gr4tuUuqHprja2loPZyeJhNrsRwcsBoYpnf
1/MWlDYrYn35+e6+EMmbZq+hq8Ats7qM3TOBTlaqcKWM76hiYIcQ9/rq4m2YuLYUkU3/b7HQtw5c
k86NJueIUHudgNoN78dIGGovglUF2iAKTdAdgdlxqbxiMwayat+xoWEZRFfUEUV5OO5qfOmxlGGE
OGgQJEwn7UTWCwZ3m/b9ugS8fWio2Yc1ZOAMp4eBIIMQvOYQdz3CsVGf6Bao1YWOwyJ0OG3GYlt4
S2R0K8H+mpyezSPocNtwEdz+U1wI0yePYmC994vIWqFGLszXMC4PlFyXzrGv5pBRRaEX+M4ksU4J
k3/kLPB+v9wah3H6zcwi74lRgw89ZL3C7n4wPo5YeD0HvrTB3Paer0BbCl2IWAvT18edEomrMhGJ
8V730wseYTOdPOAfaFzYfTgjSSpzrdQg5q/feQTzw7T2OkXrXMYLkj/oAB2BiTQp9FFpS1zqehHg
xFacp9HLO8JUNebGiNbq6gcXvZBuieS1MbRk8Psq+Jwv5pfgM3a1tMlUboGEi9hAB5e7JHJtSkiP
Lze3w1x/uqWyRuzqE+aXdxNNphrTr+g+o0NaozHFm7Brh64NFziEtyC00+AvJwrRU8/6RBWrWmNJ
ne18A15J2+HH3EJx0kkOuA+fxgFoIs6rbEQKCtQ/w12Cx66ApLnu07OQ1f3gCWC7cjzRNv8AWU7W
RIJ+K7rRhOKEAtQpxhvbiY902t+Orr5/WJCQ/K1+AGlcOEH38p7Wj6pX3NOUMeXnhHRnutjAdmid
Q/gyBmSwMCycocN8UUW4NOqz9fWIkyhMeHJb9Miph9X9V3JMvIlZdmOFp9HC0xsmdm5wVRkiMbv2
HVgA2o06lp3RUHfk0fHqY8IGEco3fXpU/KWBjHKJLa9UBv0kWPTGlEI6sS6XBBTidtmNZPTR5cOH
YdM0zN4/55XYSbvF9SqX6Juleg6QdEZ7UZmVa9lyE8BxYpQRpX9m8MKfHLC33BPwfe1d00gvF6wk
kNcOHnW/rbdO+Y3PPcRXFw3QZZXD4y3rC4UoTIf7XEF7x9ZrMtP827rBdfY5DL0Eg8kQweo4+anf
ofzkjsqcLeo1J/Gfqlv0uE/NZFFA3HMsLIo3hUTmtaMWUjax6zOkLyxI/VjXnzW7wEYhPZldauX+
1/l2aEz389hAmPhFjvBAUvxSu5GyPAWEYMnWq/XEuma30v4BaUFBwV1F+oX0XMGN0+8gD2z83oZ6
lVCdDk5JKaZ1QSC8KV7KZCGjAWtHkOKyfRwnnnJbRrZSjqJ4MpyzrOxo3Xr0MjiyEsOaCP7RPNwk
DQ5kdU0SniyHHN5VHrLraRW4rgmFrIBQnCH6WGt+525TduWs1q1CMa/13xJmSFbV5T0PMZGxuAaU
NhTr5IkyNlt/6t1aj3y3V+xDK6aK0m8/thzECHda2k4Yxblx4QxclmVkGIuf3Mtwpwt32/I43Jv4
PhbRJc3rmxWw1VUe58MxAgFk8MxSxfWX7yYjR+mDT/OzB/i9ZC00q8li30jJ08lov7dwk8qFpI7+
oc3uT4ZBXZmvdb+qTtwrBtjIE5pGpAkpNxV5XeQcXuQGgbVDKZ4JIZjMNMX8vQr9DZPkNctLGd8z
dXLnbO/xa78O4KeePlS6C01o2UjxkPXi1s89dwKIWrLIJmlrZ/bXyjR86TR+UI+MBfvU1YbJvxsq
Oym1TxLngpdpmqX6Sn8qluVYskknKfPJQ+76KcGPWDjyy2mOg1jlIyPE8bq71DYR4I34HwIdOJoI
xYQlLlCB/0TmMf04DAYglgTttRFmIW03K8AB45hHZ38WYkSj20NniLj64ug0kyw3LDD4xI1dFPwp
leycGiSHuWj0pt42HQ03N3AUJm4aFG2J7cnnSAfy7YVgZ7ncnV4nc8GkewVkiXSLoqiajZ9zcDDF
grx0QvVTggnPXzzZQYxutxNBlUTr0VcCEAgXkCXoA/K16hKcqZXXSEpy/voP8tUzBXhs4W9mvBmM
tMJkHWGfzavu8XmJgXAneR3Dr6yQ437A3gEKbbHTq43VIRsj52OrVSSin6ORSxHe++9YYdslIdcM
nZ1YJvvDYnL6nzmuc5mgWKVgDgORjdT9kpWq4pWp3qR1qvq74a07cZBcSRkFEnDQPjf3ZAS6GZL0
2oise6+GSAGUWoqVF4KGT1qBTV10vTlvZVwdmQ0h3FPuOAk2a2pJ04Q7J/dlcET7AokTyf876Yin
EEmA0JaUG/VM0QpWJzd5WTdAUT2yQJjEUnei7HJBvl7cCPwmPoM50uCMAj//3cDVe/gdo+mbjIvW
2QL7KnFtN3y2srJowChHPEB2WCEadZK/e9ycPntuvw2ySGrBXtLVjqcJ8XNHe5fq07KWQjZHwVQp
m1ENfjgUpKd9aALceDZvaEQfMtPx+5L3COZMFSYRcyZ8TMtKgOUwaJpa5Obgh51Jqh53UdD+gDWf
rTg0nT3eXeKi3gbfYcFy0XVf11W2TkG+hvs/jFF73BHEWEZd8qDGX5K1uHyrDz4Kl8wLM+b8rLzX
Dv+7Zp3o6mx+t0R164P936PUY+v0mRD/5CK5zihpe5fi9MTDa5Egkzhj57iQIOS8OMKQBZi36cDm
uDwd1ea4jmPp6dB4/q0jdDYqG+WZopE0BZywsmZfwgHst7N6etLhCX9NTTsZFybjz9QNsLjtoljx
q8XWR4q92Aq0nGoDby8yRHdoWB4wN9SNM5vLHPM1v70I/qX9vrNB4zRx77znJ3u+u7wOpAbiI55m
odeB3OowHK4Qj9N58l0CcvvOw4vYqRFDv9OHhoFBB/EKqg8TNvXwerE3BgOuWUoScMjEY19Av2Of
hgn4xITp3vj+sDOdc/Uj35WNDri2cRzRyLQ8qt1+bTGQsWTJcFfyn1gEB4t/2pi6tDWakBio0Ze6
brlfbWt24mbFIg1KTExXFOVRMsfyySvueJV3LCXjIUgETeS08gGM1iI5YLJKfwycDgb+mXyIxUD3
yy22OarW9+4nS3gPmQ4Zk32aBJj2Vz0zGP5I1cPfrGMQ5KukgjrjKMHoNllTkyNqr6u+IOF29UQA
myJYEcQq+Mx3BkvUuCafOiGQuSatArXd5qM+ghIFTRLtgfJShFUYpiO3H3clnQPyT/RtK+7u8v67
UUQkOe1D6gJZ2xRHauJ0tWzNCJXR55U4fRyqrIvKmOZ7RSf5hsDb1mmiYXi50+ezwZn2dqnhNkav
9pnPvh7CrkQtMo3NV8AS6QhIuq552w6s8qz1aTr4c2k3B99m/1sfRuHVtlaRm6e+PnNzoAU60EE9
+9mjF3Aiavb1mSHGG8bRicEh/0Ab8YeLLxKVy+R2wLjgd4qDqeCC6YVmNvH2iNrUotGQgZTNhHUH
tNs9qQ2GgUEOStq95IqGwl3AYg92sSVQUrjQGI8c++/ni6pRYuNJRhXauoX9wyvU3OGDciy9knBd
xhbZVFK2eKvrVsXTZtz4r5aIG5XfY+KZfIpw4J9B2d5w4Kz6EvnR5GaHpDTF0Fb7igHj4TuAyrzx
eUpdaqgOq6pf9sHYCAg+EIiI+2maASSeV+NVX2OHs43+pNOtrmorbPJpzhOFJ7vvez2D1Y5pKecQ
fqkMeHBcbEQ0ngJENdQ+ZUoyaEcLhLTRb+CxshABm3KZh83O7jig3xPc2KSE/tKwsEsVYgaBv7eS
LcQ01K1IViJ24J9kSFm9p1vkwrJeLtS6fFriQKIPppLmBA0Ys69A0CA31Z3+cYo2wdesvA41MWa4
W03XzjSRzGOkr9/T/eM467ICv5EgalyJ0Wc24c63uTl58Av2WPa0lrpMNm9t6dHlu8JgwvgBWkuy
zbsPKjpmRibRvhTiJU5YQQGpdUmQm0AIYqYmux6IqhEW1mCKpdnLyUxalEj2rdp3ny1uaCyslo7q
x904oMV/ei15CJ080iTJ1tikQSzpFQVuCv2HNunXmh/fZopHdi/lY5lKMJSReXfUoF0KMVH0+ytg
208FTLB7mwwMHJgh9mxXq0gVv0T+2Z1/zy/Lh/AUVVL9GcYXzcLOdjFKCP5FxP8sLLTEr+4ol3Tc
b9nFxWiWT+OlOH6jnpx5SQpTfNkqr9bcii6VgtVvUBzAexp5jePcn/lETd+8gMeyArBuxrwwvu7N
yl99j7QbZFebY8UlGU6KOyd4fRL/SLyXbkXoOtejzQrM7uY5xqQLkHQtAVmBdmxOltCBPUvj0/IO
v++8MYPakin0Hvv/wSPRhIk4a9xMfkyvT3vM59BigC2e0IJxwV+IxrnLecp0nYSw8QdHccl3SJrA
cBqwiOIFkBs4b2vy1HMyusEcxxUADVwTq2ZXXXyuyIKRsNxoDr5seRa1pm1KVqUUB37AwmwLWaIv
egrcYHMdUNYsO0bTO5Qo0PyRol3UtTIDWK8jYBQW83seZEjsY4JyY2o9tCfdkTyvwYB2/g44pqaD
iRv1ut8SrWKYiuhEfWQeyVuhjwlu5hLn5VDjMxH7WGtwUxcA6Ykjiov96XE9ETyEmjO8r58MXbPY
nS5k3JDR/6jz9+tcfMm2eesG2gCZhUyJMxJhGDUSNEeBLtNF7fK0+lfMHOONlXH73Z0aclQDR3Pj
wYOV12x89hbbvNyqB4OHg2Amz81ercH8oqbw8RnVnaKhW5JwxOkifLzO7f15X2442wwOVrBNZ5Wf
6S1diUUmGTac4S7E2jXiV4h6x8g8q75Dzw7eq80CPK7LsV7fv3vKV4RgeH7CZ+QxjqQw4poGYQps
71EvS9IzRW2A9EQBVQADu3494EuZoFVaRLxeCUridpHLDr14AJmEjJN/E9aaPApwiVIXSGroggik
bw/ke1986Jy2i0551UTLagoe43ihYCA92Pk54BvndwlR59Kymc6JWSr+vaUVvAA+k1v67ZSiy2E2
E86s7q8fkghcN3lLP20bKsRmXM8DZJUQZSiJs9ybGElXo5+m9kgV5irXqNduX/Q5Hd57obvlLxwB
u8M9gpVO9dOxh/7yxntmL3dzJ7ySFyKcBrgffeCZPWS8WPgiHrA/QS0gi/02rU0b2TfN7rJhOZKz
XqC9NHVnO0Mt6v6HEFaEpFETPjOBqhD4W8XjIZI38jDAE1M3lAErY5BE0ZldRecxwwXt5xsdruiN
gc1JDsbRQnqeGWivX4nFrA0bxY3O5ncgBo51iVeFbnhC2y0TaeG/yC7DZRQObHVWGh7g89uE6nal
t77hYOcWyzw+D5BW93WXeYpuN/bZw1dLHl2aa1lBK7Y47RiP7fMKwOVPsrIzz52heLLgdDBZLFpt
8bpZhfyumVir2vIO9CGkSpm3czFzEnWXU+XDl9thEYpnkELla//UzjsGKhW3WLuXWSmX7ri7vO2D
vB5FmVjLozahs1tLcIHM0jA9iweBrSfmRP89CaHi47MPPesHzEyqNmcbJp/Kp2DlTjR6Ttp3Lgae
8nNpJOiU85EOtMY97l9q3SUwpCvvFcx7Eg03OqNgxrpP5/bPWcwQDan77yZqCA07uNd7crt1pZeC
5+mgWUwpbNP03Nks1RzxHSiQYKRIHSLzaC6eEj5nLQIAdgcRQ48CTXhdhz77/BLKko17w9e75mN+
Fj8+0s3t7YX+/qReTW17k/UAfQZz+diPRYsmNyEFyADCHEtFicz7+eScYce6HAll2TlMF1oGMNSE
DpsWZPJgg7y9Relnd8aG6oVos7UKTt9QTMtNHZRIU2dEOUbZtTY6f0LbEGCYOs7HEh6E6TeIQAgx
I8giR7HZrx7ONUyxcAStniwCQ7QVorSNUOQnBkPCMg6kCW6nzeYBk5Nc758dX4zR0q/vRPk0M46z
uybHwOlORE6owGa296x/lu80K3Tmdlgjr82pi6Y3mYmdwetCftbPGzhzaoDo/OkuRy0NWAd1ZDMS
TuBFQyjSHyxT0DjJqhWwQiVV9M8mvQxrFTq7GJGQ9agEezV5A5sru1QyInm42J9yr0tmDtPhzTpR
OM/ldWbY4DmGU5S5lDqkI2Mz3AdeVOc9xFwOAkhKZsEmzE732Yh+TOlsVl+mqk51/FnNzAT+f8Hu
tMRo22E3AO/I7P0nZzli+chkJQhNZ6QLFpfv2xB1zgkf3BUv5woSsN7A+tJa0spgX3b2MysljTGr
kByL2/PHX0quggD5YBiHQnN5TPykjmC7WvrKML0oIDkOtZbGINimlCjmIayzindnyRnub9Cp5ufW
SyshPyrCwbu+gEBHo8hVcJBx0TzxQA3Mbispc99PxQbZ6f6jLaArtML0Y/j9HJf+sVykYSDYubYh
Xipe2D3lFpRWgNdgvr+q1oWZ0L+hlMEJD6t/lA1dcSxWw+mY5oZNHuxGaVo7OoNfTnfOeJR8GZ3T
nEj4/JcvvZo56ASMOeDpYH+Z8LG2PcinaM3RS5XCw1Lt1NjUcuJjLGQ0JuYg50K26D9GazVNxlhr
dT+FZyOmCYDdEgnACigCgUdt1SCN1Muz7IbMBHZVtHtKEL31EUgQVoOfMj6z1v3EJEQ9GAh+h0zu
Z/C9Yn//KJdJCSncrz0jispY2FLyh08Ug67cxngRchpkY3U7213emaoxQgiWRipYMoC6HK9ZTxd+
1RIAu8pzsLcWwUlBL4byH7AWAbR7JrkAlXhBRMLva3vyuQCqKY6B24pHUUqQ8IZi8iIRx9sZ43Bc
5ehzfuIuw2F+wc2pMTALdELhXWtH4HJ2KYrNBbSbqFYHWUKJ7sJ3paydTFPgUgPstmik+lmB4tAT
fWJiK++ddCAMD8BkO2M+d94FBuvPT3TC+aeE4SzTwBg5LgiJ3qQKORNVEdpJe69ZtjBwIwbxyj/w
odRHXIsGnihIpEzJzHD0y+VmJRQjmov8o9mJCA0fPJgZ3C7v0s0rRWtKTLmTQazHH9wEQltedP95
tm5fyna4lh8AEHxrDlPWrroGg/xPJ62+iWuhFFOIw70Wdn09q2wTJ7wkuo1WVOxb/rAWNpoC04Tp
ViaDkC8XsyIGmv9V218dsuta60ajnOisyBRdJIRxP4B1Rj9g5ighqXyPk1mSTLvvmXIcUKXsBuX7
B5DFKhEegceQrjIxFjARKU2SMROnxLPT1E6JbW8ofnK1E+duGBNL/8nuIdFQZ9lmqR796Ry1Awm4
cO+u/HnI8gX8y3Q1j9NL83wO+gK9lPIdsNVO6Ca4eKJVx6AGaz9YCXMMKOaAlLV4FsGKiDhU6IRq
7qdr2XeDN7MHoPmJy1Eb7iI5fMMhH7OPReEl0U3iojOfibuXuC4fxi6Slis6kT8UQWtS+IMjUOUX
fpaJWHYDVzQXXylyOytn1pYg5SN5chyDdnNg4wmdy3WPkVnqJn9UDyAL11NzLA0OlDCIiTnwUv6O
tvbrrmfMa4n0pCt5K6tGyDGYr/4+Ullv9gJiMNsz9vE82uw/Lpbet8AluKyfHB5sBTBpEdH910/b
mtMSf/WApEyKc1Js6K3fXeDXG+gL8S4lExgIKiCUaSUX0T5LlY52WjoA4dmBeoY7leKeU+IOrQqU
zCCIeunX3SlJCeDrizFIjeZNKTUwJAyoM+dBW8aoekf30GGz27PwZDkpJaI21bfvqYz4rqZdQY0a
bbdHwfSesRVajibzKhgvQ05LLkDHV44rXpn9wd9ycLHmVlrPu9QR4CD5ji/Qolr0DoF787YQKF1C
QTKck/hCdXXpwZ5YTNAT/E9n/vvjpcNX4biHta9+XO+YmhdM4eJVJhtcDdNps6mGH1/+507YnVaE
U9ZoZfPUz29hPF79dHvE8NHTLaeEXloW37W9JuzVCM71Aq3CTCXWwbiPg3IEZyhWJ3NMAM1KPX6k
CbESpcLyBiOY0tQp+vGmTBC1b9u5HLEh190OyP48UNlzkKuhZLJl7fgCDn3TKTJzd5iOQZzRobOb
AN42zehRo357d7DBdKbL0aCRGAFYSrqgQQJhXibnyBvEiZ2YqWob/m1wErU66J+EzB0wOIjkVq6O
WHWCvLLwfIBh5FQIOxzsFn7HrzTDFljx7L5oqGtTyRdlzB8ZWqMF+SabtGmbDN68G2zDjloGmCMh
6QHeB9aJE1GBmgHzu/EnO77IBZvDltmEFWv0ANEF7+IcxxZdyVkevIlbpDJb5bslqpvREa/ls6Ma
7iSxsogwOGfzLRD72Nh8CczNpU6BBzs35f44w+/TCzI5EnWXiDF66JG8SHSaSQ7Am2l3FLZ0vKQr
6SO/OPtHUH8ZkFNOKJ1b2KuxFGpn3EM27LbkwXUN76eJ+zjye3ZderBquhVLG7Y1Jntx5NnrvCJT
UH6Wrhu39W9ludnvz6Vp53Eyns18nyea6rsaaNXJW25AMBpka757zFr9ZkQZIMv7BIGmrWMNsusD
7O0kltYBQljsygXAesJJykNUbiepHNdhgwtVfUyjEj34lLSLF+CbxOhbfccbUZtTmY0zsgsmXxKv
JAFGIyABb/oRf0rK7rDLoM+wx9OkyG9DZt4IY7y+I2w/D5BSIR7gY8acfCDjZRBxQxwpogxtaGtP
ArsjJ8DRboXyRDhnAs4KHQOz9VudT1L7v8cX6/UP4w1z00ZX1MZz2x/O3J0xS7YX2mLWxzbQO1OM
tzS9SlmoONG+f0oTWAvSb1+9VPqApptFEq4uz9R4oI1BwUcVEi8iEy+H6yyEGl0MOHETMG5Yxe/D
OXqrYc2/8IXuMe/7hLIe72FRPBcQegZq9zf5MNdbWJlY1Sk234CcktJttnyc+CgEq9eASPwnHEzw
FVkcPVm5miRjeowUVNBxGuvNCFkCjxbSryGTJlZ76J8G8DyjqnZjBuE3CtB3ylXKvRm+rKiJa/pZ
tJK/2hSB3f5AQ9pmslJTAlhLv3pPwxh4oXrA0A+mcqG4qUP1/eRUeeB5r+oBz041c5O7jSAwfU2X
dRZWb6IdaF2xG+QpzNDfeQAYu5x1m3E5x2zdlSJERgEUPo6bPr6cl53Ui8mKJSxd+zya1e0ehKdK
/GE/UXMwRq4y7b8o27Km77oVFnZFIq4dqvSK+dOXvBFPcv9vkDomBFdXl28PJHSEd2QvlWM4cRgU
LBZDy8GJStSCGHbV1PTnjQ4hHMHMLP4WBdcjSVyoAE2Hu+WQnqmZGboLwpWhc+bHUzEZ7hpdrXiL
zavWsLozUngAn8vd3gPrKPUz9RBuTLT6RhTF594IqVtOW/O3fCUkKv+zR+OoITFACRbvUOWNtSGh
WWHclLMfmrrz7P0JdEl5UFh89+W8oCpi+LyOP8S152TxghGl2188k73p413jedNV4vxjQRZQnevK
TzbVvoKKrND0HGMtGRdo9ae56XmqAtGKR2T1MnXTds1f9SYRus1n1Ms0aufJ+D3F7r5h4oXj5vRF
cGBA1ZmYIpXaks0WXWTvB+zSSL26Zo79mztJtTvQz6iWpsxI+Zo4JCCDcf6pvP0nFGx8knqwxsty
3AZKpV4qdp54dzayM9ChXM5PeEFyyUBCwrCQm3es+htT5v0T8pzDbWUOH7WQNcbU5sNCvel/o9HY
xIXzAMqhYnGlTXmqQAABl1RbXvgqSJJnrjfBoy03W8ggp5/xiwwZABLauJGXYIAenqf9LqBf3wQN
uqTLzcSWt+CND3ZuGKK8WjJTa0d6EzBtUY80G/Agd1sIc+tC8tR80rLcXI+ZhAbXiN1dH/mozHy4
hrAG1xRLdPIfJEzl14bloZCu4CjOy4uAIeHaduDaWCzqlee+rM5L60DYI5Q9NQ4RFaJpiaifxF7j
g20DZgto7KhcH/2REY1bRFAAbp6Xn7SE+hJQfqOyhwfUMuV3yh2ZL1CUs2FCNMwdhVOvZnyEXafC
XD0Z11EQ3IBU3JQMiCURxFgKZwB+5KJOm0gPFzaJNi0ENanITDanPCthq2WVffi4nGKTdrx4RVpJ
xASS0ylbqLebQYXYOqlTURkWBuI9TsgFGxQXO90TNZVqA9R21P34p9x+2Z3delvWuugkl7JAVz+s
D1WY9eaBMnY0PEhLWYKBB41kBwKobmzdwlQ5zRxTdSlf7Sna/GpjclVzM/KcO5mwzRNwisEknWDC
HZcrXRM/NUy6OpUICMUM/Jx75JgbtZ1cIClFIiRzdVC8BW7s5N0rE16OFBwVVrBcl2p6xac7cO6M
1s1JcbVArFMqUIdS9eWSjnS0A9L/HVViNrUZNyBoTs/pjjak+w7KhS2IgF+6T9O1uvu4NJvIFaYj
EAF7TDzulY0eO9FT+ljLANrRfeidU1szcFl7lkljPGrUmE8YvePAIrixMRsIKY2Gfyx2OE/k9+no
j2DCey8ZaaZD24cnyK8gcWEr6M7uV8kkYg6dmIZrhJFHEXWZOo6ZXK5jLowMT4X4FFjN/bHLuIh9
WABp/scbTcWjqX7rcXvuB9ANIrq9wHlaPNmZ1tk9AL40Hqz2OMRVugCtkEYT93XRZg/wD69DOzAz
pL0sIre3mfQdxfhxfgIu2faxF5QFwbmk+Wdd3DcJ89/gFkq3VXSHbfayrRZoDXTvVdTh0dQSkPki
khDAd+4zsDI/B0Z4hSCYKfBcd1/xlx90bjje8oR4qZ2IXUpcQiq3tC27UpXyWfQbnC7I0LjG4MBO
+uSe1crJgojlUtf49YAtffwIsTnm/G/ocUPbh7IxKigepk2ghoNflaepvVESMLt5gyuuvVcAk7+D
7SJmDqRGR9gnloRZLzF6AJD5NqhbUZko7QNWQv59qVMlTNiQJ3Z6aotKN0he5il9Hpk4j+y8cOXX
vgc1330zyHqDs5brorytd7bSptiwUeR9NpTu3dN+45S2kOlnr2gykZapQfj/ZF/sZDkp7poe7Ymj
PtVjlQTvQ02nr1IiOkQJIYiodnsv4Gxxc0B9O4LaKXasAAUA

`pragma protect end_protected


endmodule
