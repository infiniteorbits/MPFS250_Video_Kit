--=================================================================================================
-- File Name                           : Gamma_Correction.vhd
-- Description						   : Supporting both Native mode and AXI4 Stream mode

-- Targeted device                     : Microsemi-SoC
-- Author                              : India Solutions Team
--
-- COPYRIGHT 2021 BY MICROSEMI
-- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS FROM MICROSEMI
-- CORP. IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM MICROSEMI FOR USE OF THIS
-- FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND NO BACK-UP OF THE FILE SHOULD BE MADE.
--
--=================================================================================================
--=================================================================================================
-- Libraries
--=================================================================================================
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;   
--=================================================================================================
-- Gamma_Correction entity declaration
--=================================================================================================                                                                                                                          
ENTITY Gamma_Correction IS                                                                                                       
  GENERIC(
-- Generic List
	G_PIXELS			: INTEGER := 4;
    -- Specifies the data width
    G_DATA_WIDTH 		: INTEGER RANGE 8 TO 16 := 8;

    G_FORMAT		    : INTEGER := 1   --  0= Gamma_Correction and 1= Gamma_Correction with AXI	
    );
  PORT (
-- Port List
    -- System reset
    RESETN_I 			: IN STD_LOGIC;

    -- System clock
    SYS_CLK_I 			: IN STD_LOGIC;

    -- Specifies the input data is valid or not
    DATA_VALID_I 		: IN STD_LOGIC;  
	
	-- Data input
    TDATA_I             : IN STD_LOGIC_VECTOR(3*G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);
    
	-- Specifies the valid control signal
    TVALID_I            : IN STD_LOGIC;
	
	TUSER_I				: IN STD_LOGIC_VECTOR(3 DOWNTO 0);

	-- ready signal on slave
	TREADY_O			: OUT STD_LOGIC;
	
    -- Red data input	  
    RED_I       		: IN STD_LOGIC_VECTOR ((G_PIXELS*G_DATA_WIDTH - 1) DOWNTO 0);
      
    -- Green data input 
    GREEN_I     		: IN STD_LOGIC_VECTOR ((G_PIXELS*G_DATA_WIDTH - 1) DOWNTO 0);
      
    -- Blue input  
    BLUE_I      		: IN STD_LOGIC_VECTOR ((G_PIXELS*G_DATA_WIDTH - 1) DOWNTO 0);
	
	-- Specifies the valid RGB data
	DATA_VALID_O 		: OUT STD_LOGIC;

    -- Output red colour
    RED_O 				: OUT STD_LOGIC_VECTOR(G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);

    -- Output green colour
    GREEN_O 			: OUT STD_LOGIC_VECTOR(G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);

    -- Output Blue colour
    BLUE_O 				: OUT STD_LOGIC_VECTOR(G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);
	
	-- Data input
    TDATA_O             : OUT STD_LOGIC_VECTOR(3*G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);
	
	TUSER_O				: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	
	TSTRB_O             : OUT STD_LOGIC_VECTOR(G_DATA_WIDTH/8 - 1 DOWNTO 0);

    TKEEP_O             : OUT STD_LOGIC_VECTOR(G_DATA_WIDTH/8 - 1 DOWNTO 0); 

    TLAST_O				: OUT STD_LOGIC;	
	
	-- Specifies the valid control signal
    TVALID_O            : OUT STD_LOGIC
	
    );
END Gamma_Correction;
--=================================================================================================
-- RGB_TO_YCbCr architecture body
--=================================================================================================
ARCHITECTURE rtl OF Gamma_Correction IS
--=================================================================================================
-- Component declarations
--=================================================================================================
COMPONENT Gamma_Correction_Native 
	GENERIC(
		G_DATA_WIDTH : INTEGER RANGE 8 TO 16 := 8                                                                         
		);
		PORT (                                                                                                        
			SYS_CLK_I         				: IN STD_LOGIC;
			RESETN_I        				: IN STD_LOGIC;
			DATA_VALID_I   					: IN STD_LOGIC;
			RED_I       					: IN STD_LOGIC_VECTOR ((G_DATA_WIDTH - 1) DOWNTO 0); 
			GREEN_I     					: IN STD_LOGIC_VECTOR ((G_DATA_WIDTH - 1) DOWNTO 0);
			BLUE_I      					: IN STD_LOGIC_VECTOR ((G_DATA_WIDTH - 1) DOWNTO 0); 
			RED_O							: OUT STD_LOGIC_VECTOR ((G_DATA_WIDTH - 1) DOWNTO 0);
			GREEN_O							: OUT STD_LOGIC_VECTOR ((G_DATA_WIDTH - 1) DOWNTO 0);     
			BLUE_O							: OUT STD_LOGIC_VECTOR ((G_DATA_WIDTH - 1) DOWNTO 0);
			DATA_VALID_O 					: OUT STD_LOGIC
		);
		END COMPONENT;
		
COMPONENT Gamma_Correction_4p 
	GENERIC(
		G_DATA_WIDTH : INTEGER RANGE 8 TO 16 := 8;
		G_PIXELS			: INTEGER := 1
		);
		PORT (                                                                                                        
			SYS_CLK_I         				: IN STD_LOGIC;
			RESETN_I        				: IN STD_LOGIC;
			DATA_VALID_I   					: IN STD_LOGIC;
			RED_I       					: IN STD_LOGIC_VECTOR ((G_PIXELS*G_DATA_WIDTH - 1) DOWNTO 0); 
			GREEN_I     					: IN STD_LOGIC_VECTOR ((G_PIXELS*G_DATA_WIDTH - 1) DOWNTO 0);
			BLUE_I      					: IN STD_LOGIC_VECTOR ((G_PIXELS*G_DATA_WIDTH - 1) DOWNTO 0); 
			RED_O							: OUT STD_LOGIC_VECTOR ((G_PIXELS*G_DATA_WIDTH - 1) DOWNTO 0);
			GREEN_O							: OUT STD_LOGIC_VECTOR ((G_PIXELS*G_DATA_WIDTH - 1) DOWNTO 0);     
			BLUE_O							: OUT STD_LOGIC_VECTOR ((G_PIXELS*G_DATA_WIDTH - 1) DOWNTO 0);
			DATA_VALID_O 					: OUT STD_LOGIC
		);
		END COMPONENT;
		
COMPONENT AXI4S_INITIATOR_GAMMA 
	GENERIC(
		G_DATA_WIDTH         : INTEGER RANGE 8 To 96 := 8; 
		G_PIXELS			: INTEGER := 1
		);
		PORT (    
            SYS_CLK_I         			: IN STD_LOGIC;
			RESETN_I        			: IN STD_LOGIC;		
			DATA_I         				: IN STD_LOGIC_VECTOR(3*G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);
			DATA_VALID_I   				: IN STD_LOGIC;
			EOF_I						: IN STD_LOGIC;
			TUSER_O						: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			TDATA_O                     : OUT STD_LOGIC_VECTOR(3*G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);
			TSTRB_O                     : OUT STD_LOGIC_VECTOR(G_DATA_WIDTH/8 - 1 DOWNTO 0);
			TKEEP_O                     : OUT STD_LOGIC_VECTOR(G_DATA_WIDTH/8 - 1 DOWNTO 0);
			TLAST_O                     : OUT STD_LOGIC;
			TVALID_O                    : OUT STD_LOGIC
		);
		END COMPONENT;
			
COMPONENT AXI4S_TARGET_GAMMA 
	GENERIC(
		G_DATA_WIDTH         : INTEGER RANGE 8 To 96 := 8;  
		G_PIXELS			: INTEGER := 1
		);
		PORT (                                                                                                        
			TDATA_I                       		: IN STD_LOGIC_VECTOR(3*G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);
			TVALID_I                       		: IN STD_LOGIC; 
			TUSER_I								: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			TREADY_O							: OUT STD_LOGIC;
			EOF_O								: OUT STD_LOGIC;
			DATA_O                           	: OUT STD_LOGIC_VECTOR(3*G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);   
			DATA_VALID_O                       	: OUT STD_LOGIC
		);
		END COMPONENT;
--=================================================================================================
-- Synthesis Attributes
--=================================================================================================
--NA--
--=================================================================================================
-- Constant declarations
--=================================================================================================
--NA--
--=================================================================================================
-- Signal declarations
--=================================================================================================
SIGNAL s_dvalid_slv	        : STD_LOGIC;
SIGNAL s_dvalid_mstr        : STD_LOGIC;
SIGNAL s_eof				: STD_LOGIC;
SIGNAL s_data_o				: STD_LOGIC_VECTOR ((3*G_DATA_WIDTH - 1) DOWNTO 0);
SIGNAL s_red_in				: STD_LOGIC_VECTOR (G_DATA_WIDTH-1 DOWNTO 0);
SIGNAL s_green_in			: STD_LOGIC_VECTOR (G_DATA_WIDTH-1 DOWNTO 0);
SIGNAL s_blue_in			: STD_LOGIC_VECTOR (G_DATA_WIDTH-1 DOWNTO 0);
SIGNAL s_red_axi			: STD_LOGIC_VECTOR (G_DATA_WIDTH-1 DOWNTO 0);
SIGNAL s_green_axi			: STD_LOGIC_VECTOR (G_DATA_WIDTH-1 DOWNTO 0);
SIGNAL s_blue_axi			: STD_LOGIC_VECTOR (G_DATA_WIDTH-1 DOWNTO 0);

SIGNAL s_data_4p_o			: STD_LOGIC_VECTOR ((3*G_PIXELS*G_DATA_WIDTH - 1) DOWNTO 0);
SIGNAL s_red_4p_in			: STD_LOGIC_VECTOR (G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);
SIGNAL s_green_4p_in		: STD_LOGIC_VECTOR (G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);
SIGNAL s_blue_4p_in			: STD_LOGIC_VECTOR (G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);
SIGNAL s_red_4p_axi			: STD_LOGIC_VECTOR (G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);
SIGNAL s_green_4p_axi		: STD_LOGIC_VECTOR (G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);
SIGNAL s_blue_4p_axi		: STD_LOGIC_VECTOR (G_PIXELS*G_DATA_WIDTH-1 DOWNTO 0);

SIGNAL s_data_axi			: STD_LOGIC_VECTOR ((3*G_DATA_WIDTH - 1) DOWNTO 0);
SIGNAL s_data_4p_axi			: STD_LOGIC_VECTOR ((3*G_PIXELS*G_DATA_WIDTH - 1) DOWNTO 0);

BEGIN
--=================================================================================================
-- Top level output port assignments
--=================================================================================================
s_data_axi     <= s_red_axi & s_green_axi & s_blue_axi;
s_data_4p_axi  <= s_red_4p_axi & s_green_4p_axi & s_blue_4p_axi;
--=================================================================================================
-- Generate blocks
--=================================================================================================
FOUR_PIXEL: IF G_PIXELS = 4 AND G_FORMAT = 1 GENERATE
s_red_4p_in 		<= s_data_4p_o ((3*G_PIXELS*G_DATA_WIDTH - 1) DOWNTO (3*G_PIXELS*G_DATA_WIDTH - 1)- (G_PIXELS*G_DATA_WIDTH-1));
s_green_4p_in 		<= s_data_4p_o (((3*G_PIXELS*G_DATA_WIDTH - 1) - G_PIXELS*G_DATA_WIDTH) DOWNTO  G_PIXELS*G_DATA_WIDTH);
s_blue_4p_in		<= s_data_4p_o (G_PIXELS*G_DATA_WIDTH - 1 DOWNTO 0);
END GENERATE;

ONE_PIXEL: IF G_PIXELS = 1 AND G_FORMAT = 1 GENERATE
s_red_in 		<= s_data_o ((3*G_DATA_WIDTH - 1) DOWNTO (3*G_DATA_WIDTH - 1)- (G_DATA_WIDTH-1));
s_green_in 		<= s_data_o (((3*G_DATA_WIDTH - 1) - G_DATA_WIDTH) DOWNTO  G_DATA_WIDTH);
s_blue_in		<= s_data_o (G_DATA_WIDTH - 1 DOWNTO 0);
END GENERATE;
--=================================================================================================
-- Asynchronous blocks
--=================================================================================================
--NA--
--=================================================================================================
-- Synchronous blocks
--=================================================================================================
--NA--	
--=================================================================================================
-- Component Instantiations
--=================================================================================================
GC_1p_Native_FORMAT : IF G_PIXELS = 1 AND G_FORMAT = 0 GENERATE
Gamma_Correction_1p_Native_INST: Gamma_Correction_Native
GENERIC MAP(
	G_DATA_WIDTH => G_DATA_WIDTH
)
PORT MAP(
	SYS_CLK_I		=> 		SYS_CLK_I,
	RESETN_I		=>		RESETN_I,
	DATA_VALID_I	=> 		DATA_VALID_I,
	RED_I   		=>		RED_I,
	GREEN_I 		=>      GREEN_I,
	BLUE_I  		=>		BLUE_I,
	RED_O			=>		RED_O,
	GREEN_O			=>      GREEN_O,
    BLUE_O  	    =>      BLUE_O,
	DATA_VALID_O	=>		DATA_VALID_O
);
END GENERATE;

GC_1p_AXI4S_FORMAT : IF G_PIXELS = 1 AND G_FORMAT = 1 GENERATE
Gamma_Correction_1p_AXI4S_INST: Gamma_Correction_Native
GENERIC MAP(
	G_DATA_WIDTH => G_DATA_WIDTH
)
PORT MAP(
	SYS_CLK_I		=> 		SYS_CLK_I,
	RESETN_I		=>		RESETN_I,
	DATA_VALID_I	=> 		s_dvalid_slv,
	RED_I   		=>		s_red_in,
	GREEN_I 		=>      s_green_in,
	BLUE_I  		=>		s_blue_in,
	RED_O			=>		s_red_axi,
	GREEN_O			=>      s_green_axi,
    BLUE_O  	    =>      s_blue_axi,
	DATA_VALID_O	=>		s_dvalid_mstr
);
END GENERATE;

GC_4p_Native_FORMAT : IF G_PIXELS = 4 AND G_FORMAT = 0 GENERATE
Gamma_Correction_4p_Native_INST: Gamma_Correction_4p
GENERIC MAP(
	G_PIXELS	 => G_PIXELS,
	G_DATA_WIDTH => G_DATA_WIDTH
)
PORT MAP(
	SYS_CLK_I		=> 		SYS_CLK_I,
	RESETN_I		=>		RESETN_I,
	DATA_VALID_I	=> 		DATA_VALID_I,
	RED_I   		=>		RED_I,
	GREEN_I 		=>      GREEN_I,
	BLUE_I  		=>		BLUE_I,
	RED_O			=>		RED_O,
	GREEN_O			=>      GREEN_O,
    BLUE_O  	    =>      BLUE_O,
	DATA_VALID_O	=>		DATA_VALID_O
);
END GENERATE;

GC_4p_AXI4S_FORMAT : IF G_PIXELS = 4 AND G_FORMAT = 1 GENERATE
Gamma_Correction_4p_AXI4S_INST: Gamma_Correction_4p
GENERIC MAP(
	G_PIXELS	 => G_PIXELS,
	G_DATA_WIDTH => G_DATA_WIDTH
)
PORT MAP(
	SYS_CLK_I		=> 		SYS_CLK_I,
	RESETN_I		=>		RESETN_I,
	DATA_VALID_I	=> 		s_dvalid_slv,
	RED_I   		=>		s_red_4p_in,
	GREEN_I 		=>      s_green_4p_in,
	BLUE_I  		=>		s_blue_4p_in,
	RED_O			=>		s_red_4p_axi,
	GREEN_O			=>      s_green_4p_axi,
    BLUE_O  	    =>      s_blue_4p_axi,
	DATA_VALID_O	=>		s_dvalid_mstr
);
END GENERATE;

Gamma_slv_1p_FORMAT : IF G_FORMAT = 1 AND G_PIXELS = 1 GENERATE
Gamma_Correction_AXI_SLV_1p_INST: AXI4S_TARGET_GAMMA
GENERIC MAP(
	G_PIXELS		=>  G_PIXELS,
	G_DATA_WIDTH   => G_DATA_WIDTH
)
PORT MAP(
	TVALID_I			=> 		TVALID_I,
	TDATA_I				=> 		TDATA_I,
	TUSER_I				=>		TUSER_I,
	TREADY_O			=>		TREADY_O,
	EOF_O				=>      s_eof,
	DATA_VALID_O		=>      s_dvalid_slv,
	DATA_O 				=>		s_data_o
);
END GENERATE;

Gamma_slv_4p_FORMAT : IF G_FORMAT = 1 AND G_PIXELS = 4 GENERATE
Gamma_Correction_AXI_SLV_4p_INST: AXI4S_TARGET_GAMMA
GENERIC MAP(
	G_PIXELS		=>  G_PIXELS,
	G_DATA_WIDTH   => G_DATA_WIDTH
)
PORT MAP(
	TVALID_I			=> 		TVALID_I,
	TDATA_I				=> 		TDATA_I,
	TUSER_I				=>		TUSER_I,
	TREADY_O			=>		TREADY_O,
	EOF_O				=>      s_eof,
	DATA_VALID_O		=>      s_dvalid_slv,
	DATA_O 				=>		s_data_4p_o
);
END GENERATE;

Gamma_mstr_1p_FORMAT : IF G_FORMAT = 1 AND G_PIXELS = 1 GENERATE
Gamma_Correction_AXI_MSTR_1p_INST: AXI4S_INITIATOR_GAMMA
GENERIC MAP(
	G_PIXELS		=>  G_PIXELS,
	G_DATA_WIDTH   => G_DATA_WIDTH
)
PORT MAP(
    RESETN_I																								=>  RESETN_I,
	SYS_CLK_I																								=>  SYS_CLK_I,
	DATA_VALID_I																							=> 	s_dvalid_mstr,
	DATA_I                                        															=>  s_data_axi,
	EOF_I																									=>  s_eof,
	TLAST_O																								    =>  TLAST_O,
	TUSER_O																									=>  TUSER_O,
	TSTRB_O																		                            =>	TSTRB_O,	
	TKEEP_O																		                            =>  TKEEP_O,		
	TVALID_O																	                            =>  TVALID_O,
	TDATA_O																		                            =>	TDATA_O
);
END GENERATE;

Gamma_mstr_4p_FORMAT : IF G_FORMAT = 1 AND G_PIXELS = 4 GENERATE
Gamma_Correction_AXI_MSTR_4p_INST: AXI4S_INITIATOR_GAMMA
GENERIC MAP(
	G_PIXELS		=>  G_PIXELS,
	G_DATA_WIDTH   => G_DATA_WIDTH
)
PORT MAP(
    RESETN_I																								=>  RESETN_I,
	SYS_CLK_I																								=>  SYS_CLK_I,
	DATA_VALID_I																							=> 	s_dvalid_mstr,
	DATA_I                                         															=> s_data_4p_axi,
	EOF_I																									=>  s_eof,
	TLAST_O																								    =>  TLAST_O,
	TUSER_O																									=>  TUSER_O,
	TSTRB_O																		                            =>	TSTRB_O,	
	TKEEP_O																		                            =>  TKEEP_O,		
	TVALID_O																	                            =>  TVALID_O,
	TDATA_O																		                            =>	TDATA_O
);
END GENERATE;

END rtl;
--=================================================================================================
-- File Name                           : Gamma_Correction_Native.vhd
-- Description						   : This module gives gamma correction of RGB with constant 
-- 										 gamma factor 0.454.

-- Targeted device                     : Microsemi-SoC
-- Author                              : India Solutions Team
--
-- COPYRIGHT 2020 BY MICROSEMI
-- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS FROM MICROSEMI
-- CORP. IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM MICROSEMI FOR USE OF THIS
-- FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND NO BACK-UP OF THE FILE SHOULD BE MADE.
--
--================================================================================================= 

--=================================================================================================
-- Libraries
--=================================================================================================
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

--=================================================================================================
-- Gamma_Correction_Native entity declaration
--=================================================================================================
ENTITY Gamma_Correction_Native IS
  GENERIC(
-- Generic List
    -- Specifies the data width
    G_DATA_WIDTH : INTEGER RANGE 8 TO 16 := 8	

    );
  PORT (
-- Port List
    -- System reset
    RESETN_I : IN STD_LOGIC;

    -- System clock
    SYS_CLK_I : IN STD_LOGIC;

    -- Specifies the input data is valid or not
    DATA_VALID_I : IN STD_LOGIC;  

    -- Red data input	  
    RED_I       : IN STD_LOGIC_VECTOR ((G_DATA_WIDTH - 1) DOWNTO 0);
      
    -- Green data input 
    GREEN_I     : IN STD_LOGIC_VECTOR ((G_DATA_WIDTH - 1) DOWNTO 0);
      
    -- Blue input  
    BLUE_I      : IN STD_LOGIC_VECTOR ((G_DATA_WIDTH - 1) DOWNTO 0);
	
	-- Specifies the valid RGB data
	DATA_VALID_O : OUT STD_LOGIC;

    -- Output red colour
    RED_O : OUT STD_LOGIC_VECTOR(G_DATA_WIDTH-1 DOWNTO 0);

    -- Output green colour
    GREEN_O : OUT STD_LOGIC_VECTOR(G_DATA_WIDTH-1 DOWNTO 0);

    -- Output Blue colour
    BLUE_O : OUT STD_LOGIC_VECTOR(G_DATA_WIDTH-1 DOWNTO 0)
	
    );
END Gamma_Correction_Native;
`protect begin_protected
`protect version=1
`protect author="author-a", author_info="author-a-details"
`protect encrypt_agent="encryptP1735.pl", encrypt_agent_info="Synplify encryption scripts"

`protect key_keyowner="Synplicity", key_keyname="SYNP05_001", key_method="rsa"
`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_block
WBbKVABM8Q1m+AJ/g0wjT+zywGsaPCyn2QxVvxNJ44ev5n/0SYhnisnPVMDkkNX266pSZnBvUZvm
xfLfLQeUHkgTlTedr/9yrsnE02onLouF7OiAeJ7HJfXMy0EG4VzfQUYB05tQf5ZFzYffyzlLJF3+
AkKAvxpZRAoXK76uIsWP+bhzyR4eaS2P/AhkNrsqgz+lONq6QGgAOCq/49jsUAZUvS1x7CrRuw/m
4x9s4iRNDE8vPIbiPJufs6reaKaGwJN4vw1/KO6oCbgCqZ3qzKu82bGk/4e35ZBRWF2XmL/D68fW
M3bn38PsreDWnQW26Mv0DBU+HIqlJbwK6c3fzA==

`protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`protect encoding=(enctype="base64", line_length=76, bytes=128)
`protect key_block
EJ7XVxnWuHboJtTWELv2eSNBX2G5fisZG3Eh23Rg1P+b0zzVt63JUIPjM+pr1kV3podVZV9nlX+f
NQ66WOoTvSkJmeLOpd6xEhc00rYmm19Bx+xXX0wNfgzeKB5tGAdTqnzcGo4uoBpeuHfeD6lUBKq3
YtcbBnUTXbaY/MFEXHk=

`protect key_keyowner="Microsemi Corporation", key_keyname="MSC-IP-KEY-RSA", key_method="rsa"
`protect encoding=(enctype="base64", line_length=76, bytes=960)
`protect key_block
UulpGFwduP+H+6KbCCP95KycyyHijnuZWGTCg/6cp3PkVrbQu9zK6Cje662Q3I/wIXBi5q9jvJzP
rP3BfihytC+J8ARqP4NsX0+BQnJORVPmCN3/QfTJ20biABBnQpJJilYOZTQGG7qWC5GAA8Ea0ZFv
P6UaYKbpczrgA23bLmPwhneqZ7P86WDp9mJqG0QxFi9D8uUzOw/j6EBSzO+e2yTZfCaa5gvbZMb1
CbHXmgtTlnMe89jQSg1mdPz4GEypQb2v2MVyR6UdiMV1sJEEUMrFkqpCWDXLaCPIu+r5KLZWKU99
Bq4S5znpbp45j24AFQxlG+W9SjblxEEMY6+vOJM1ZZjsELNqgZ4g2U+LHbz9u3s2Ij6FRP31yyzc
Knl06CGNCDVqE0GOSxZnMp/H0+0uYnPHEJJyz2kZaBluQKPQ4VPx7sY/+ypcWvWkNWjxBQUBR7aL
DeCL+vd5aS08LJfEwjYTyeaIDx5uiM2s7FEebM5aUouYcktylwYzTG5jFFN2z0KzXKrwlmbnl6e7
rzo988qoSpYd7pw8wZ+U4ThNHrr8N34aPkmPwyQtt/yMsuYvkZqi7/i+LGn77iPA7yHfSbu/NHGm
t3DVeTcR5fIj2+8+zfI19ANdYq+Csfpz8+vpGtv3ZtSUB1CmAaF2zpM0llGD7o//G0Mg2CfnnDGN
UGtU5IrddwL4LF+oMnIdUkVfN5gUk84ADhhEy9ud9JazkyGjyvOA+NhUh39ky1D16NC/2zVGjb2I
+0/15VBzxvdkt3bvOmu2bef8FHV14yoTo3YfTnwYp85XXXLBfhivI3iYOpeDPQ1S0+9YDBjr/uD+
9eZtBjb29xAe9AyNkMppyHl75Ff3yHtNZ0JM9Vd2xkpqFY65mrjYzlz7ld4Ob3iJW3kJW0c37I19
wQ62YcoNVDZ8dAAAAaWU/PZmBrLq38IxwGWyI/RFL+rdba6mRe3yr1joZUL7C3TYStReFZWcuLbQ
ANK1jd/WDUXLqyBETZq9xYqT6U2eJiZsRVVz45nGViTYu0XXd1xjY9iWaHAj/n1SLdflic7WyHf8
jhIyRSwNh1sFCCtNOiNobEN9WaGaRfhJfKnJyUt5eg5Yok9cRUwp3tMOrfIV+aUcZSo+kpwrA2/B
aLW/DmvZ4CVE2tULqfr7iMEznVy885s1PdZ49nUNzGvx1bQocQHZWtG72pWQsfRC5gS7xbXbh5hV
bkj+vYNzbFkELOycNXnJixghGAuCq91v5wQPhdSxcQWOFzyInbLiTK7L1GplXZjX

`protect data_keyowner="ip-vendor-a", data_keyname="fpga-ip", data_method="aes128-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=223808)
`protect data_block
RJS/k3De7FaJvBmK1UQTd/ki+bxjsyCCN3+KL8aX8RfbGmcMsKO0yQMVWL3yzg/caIAVr8vOC6RW
b9itec3gWKKjKu+XXEDKLks8RzbwCF+/6FsoAWIZltgcuibSqdykZdoWK4ob2LQ8InrAJZ1KIpN7
DFBlMNtfHr/TsQB2hXYb7Erz8m9WXvTZO5aqZgtrI/nqRYKRmiX+dvg8tBc2+a0gZunbuKBvifC8
LAXd8hNN4h+vQgJIrjkZL4m6iX8P5JuP8MBR0lhhA7mqr9tDzZnk9j+xOg5xNDcwBlGqWlTGDe45
Z5onR936JFEFmQnayxX316gkH1LIrn0WyChfcDAECOQLaZ3nihUJI2yLM/2MCh9iHdFacdTVAcQ3
oZzIS4road6RMdCrEPULcJnrHxbmjc9bzTr+h+HEWCJhnzpvsbgkhrPluxlxwfBRAj9ezudyyZ/w
RmXt8EoeMxlhGTb5yVQPGW+hq2XwRxLvFfBoLckP/s2W/kI1nb1OrKnKjHNY9v8QT3qLY17BIcxc
xAXW3PqGq+Dg7Ib8Ii0rZPjQpdqt1p1CiN6PeWRyjHppJ/ERg+CtR+LlEfFXwxwIXnoDAVUsRAQa
m4UkuDlszhtUiV8IzddsdPIIhGcdB1fQ7vJQZ87Gg5UkeA4fuNIrzrL6JXfuqoTfhLGr3n1ldY3D
jmHJajEVURQbsosfy9Rcwlh7c0uLnKXqXsD5XiB3EdbEEA1ADWbTAgqkS60Kw01dPSoaqZpwNpoW
ebUdGkQ382Z5R88Ir4pxgkdD/JpbahVSTpEpRKJHWAj9NAh3QIzzGwXPNxn9fCrFlnj+uEf8dVF4
pXrqN99WvFt2jJD+NjhqzVVb8ho40qRNtf7+7N2A6qvCcIG6NjwsZMR56vyMXX1Idg1izrelz5hr
kqhFeGyDK/TSvQLvxIQKEnMoPaPKQ1r9yn4GUaIqCSkxyoiMZiBf7SiN8cYL99PJExCNcO1JP8zz
KMFYCPt1r/Bs7umiqRqrA6zFOSRTeC3amvG62eRN9NaOe2/WI4i8IQ8azbJVRFbz+6qvt9PNmlmv
F4Mtf/OjP8mVfNaEU6uCzBIhPnsb6w7utK0y/ObL56QEKmrmYYG2kRJAZ/b0KEBUK76OIG/MxAXw
MOSqlH5juFMe55llrJ2pTBQtWI/fN8XTu3FOVjPrXDNDoGkkD0gnp7zQGfZEJswH7BDvjoR/6UtF
DM2KVcnxbGJVGBU3h+qSqWP/dt7BvPTjRUOZRejqDBKWJ2pvocTTn+krYUSIyQRiub5UEk7q/Ytm
sLrks+be6Yv+5Zk1+m24m4Za5lcCQOmsIMtVVh3UP/tgXtSIr8ulTrfzyKW383N4BkQuhuU1bqvm
v1nJeIkO7JxJwFemZKZZqwBtrEMwzNwkuvW5E4SaIZb6TcnwIYx8VDV4hpntlKs/GDDsMxhMJjyz
GWPyOQmYwntns0iIXXhV7lYBLoS17jcHJ1/t7fQEdiLkXZGGneJy31NWFpD90eAUMNIyZkbgtas1
H89/XraYHsMpmUU97VyK+aGLmt4zoZ8wTVztYpBeHFHWUvQBezdl26qbwk0zk0Q2zCJTTekD9zsW
Yf6wV+DMvQM9w90Ltk2zLJHqZW6sRAoXnIviJG9hV/D2crPhpY3Ccl+fkmTRdKmAYxqgkUCNs5iJ
4FExb/TCD4AQY0/WZ7kDV5bma71rZyDk7mzTjAKAyE2gn65hQ+mfWmXM5APT43pdrZcI6hjd8+1L
C/BwFdNfAS2VQW9lPN2Xuutni+Z6d2J026J8i/gLFlyeulFRuPkUogC5hhJqRNcDHObjGRMuJ4Iw
l7jyjq9rls8AmG6nP5i6iC+eJFdW7sFlxCAJK3o1amTtQRFYyWqlBmkP1sOSPD1gmuTBGm8LiL5Q
x5ua6BOHzBhNNi6v1v5lFswzz/yrPf2dFEvVKAS1jy8nnS2bUnTOObN7C7oUcKb1w9az+MwqyvK6
bo666n4oRm8nUjRTYW7LnQkh/WGobnC0gcQPZUHsJhXOATFiErLVxKqnKBFipMfvUbHsIQe67Lyb
cI0nBBP/Gock/O1AJ8JQSzGejcpjiumPj1tliC90vGAyHEi0Qoqw3uzQ1PrV2uC1qZdcwiraCku9
Am7pIJf3I/mrA2U74oKvwWA+KK4O+WckYba9Uq6ntJlE8mBZOvnTe6PXp1nRyfzuOOZvq2wExVaB
/4UPEZjZ2f/PfVdquvlQT56cKgC+D5Tooid+EAsuyRSAfsCOFovuDplqIG2RcgXMpbGf3NcK0rlK
GTz3nt6lvJm8UZ+R2UYv1LTCZrCv/4JxghzgI3eHoFaLZQSRrmOhuGu/UMSOdkAA6oNyT+oYOMUN
Igm3SsdDQEL+e4E745nnAxs3IkrF5YzPDxzLTNCc640iRuE4dJCkDTVKxjon8kIdxmFuFNcM8SiO
aBKravRAY58RM8WCjcv+YVtO+RrL0LP6Y0w4jVq77XwkDPQINJh1rolHJzu49LjOfwJRZHj9zpLg
KQrAMKo7yAGljPkI9PGvln5mpTSLO2FBXVvgKG2bbcy64U2Dj35rlCN3qcsuVuDnEpbdLizqan0e
t+/JLdsbT6lpyzQJMYoJKorghnmlyHkZCvt4IaLlFquus27C2XoOL6+XHSxtd1sz4TZwu5HDkeqV
LZgklf+GEc5UCfEDAAN4kJO8xTxyoyr4nqIskyYNojnMyYA92DBc7+GVeqkn+J08unMeYLrhewur
yExku+Tilxs4eaqKZMwSkZbSHwHhnkBJe2q0y707A7drWJfrh2VxxXlz6ZmtUaaTksSZhu/hX7AZ
oKmjZMPDEJ2HFguyJe0iQPaH8V9+cJIuQnUyMOMbNwMngjU8rhmfbolFMM7VnZ6fFh8Gwf7jwf3I
q7bLkADwsnre0ik8tY01Wz/FY6LhDSfSLo/vPcyX2XPYia5NG0ONJDIznBII3vis60C/L3RpoGq/
fZuIE+CSdJK8C0decLoV6pe5+16CTjbUK+K3jW7QHBwSU8nvVGOkldWn7AgqCoUrwcLJmg2bZhCC
VYk9kMbpXzUN2p3ainUzDkAbWQ+bY1FRKcsRs2FOYjQ9Hg03hVALwoukQLdnTwLC+IoM3D9j6AH8
tNAsNYGHXnY6n5gNnKet2V8fzkdC8Yiep+kX5r1SqKkqDTIuWVNMXJOxBvcZKxGRYTDA500/qMo3
YXfGMOHtD1G+mo0jTEUguQ7wiSvl2Gs0+tyxER157tdvO97MV6Mq5vmZt8Nvd1Ib74VGxCxENHtU
e2Z3EYn6dDzl0AmmOmi+YXipH8FPvaiB2053yPPQkG76QEZbZA1pqr4jnoHtO40Evhs7fi0aFXRZ
RDRHkm7DBvjmzG5oSSrb7ZbZO9N4khGChOm6aqEcXloDVcUFW0vPWpEKdDORxV5xvjuJnFlIQDfL
lQ8Bg3XfYLIW3zOc9VIgreVTHpzMUbZds5rKn3ak4BiW/GXd4ied5+0ISNHxlZkYBkN/qpzsYBJk
pBXm7xRhW+ymF4MmKGEbtqc1hld44SHIHMJx+1oLIegewBWF9JiRBJQMSXF5YWpdhI2XPFa4juqd
4rwOJ6zr5O6p1cyzc35U43UATf1IUpWi/4JpNYcTzK/aKO9xgGWukTBRFie+lh1M0QOGTpFpvr7L
8xhzcThUyyLSDo/OkwCVjEIN0YKq9APO/X1ISLonICVIz+GIjZX+ZZ3c/YmlW9IMSJ1oFhFVwZPG
Y3qQThVbsmMn/56HWMRIzNgautM3rRmzzjsiU+7DO2RChL1JI1EzAdumCFRoRf9nMvxsAk2qX9AH
fzIRlKRK7eKeZ4y0IKvMto5ag2BNuHGyYcY7iwGG2XnlN1LObFhww7clWSTV/6IpxYR1dfB/kuJ1
i7mmxs5Ph0XD05xsrk3Y5MW0cTCvfkd3to7ATb4770+ZO7Jokar3Qq3Mn6M11hVrRUZqygEy/iCw
k03q1t8Pft4v35CgJ0HjK9PsjTf+GeW2JjbtgKCf/FnVt2KrOHdfu1/1e6+6srNbuLp6+CjxX93B
RE4f7McGTgh/kab18Hgg2OR9U3Qp57+bQFv6JuubVOtVAnc/C3b3ADnTyXegM0efktcSc1PSjzl5
8rt8SAfVQgvAJNadbmym9htUbJ1dXOEbXwBVFfTbOrLaD0EE/eA6uS5/663fDW5extJjIJtNgFtY
IHe3nDZ2DuCaG+KdWBBlW9zSzf3jgXSYP+MBMilP7n2a7AKyRedQSE6nA8UueoxH0iDlvJnjAXjl
Z/2zfe9GCmlVBwh2w/QaAFTW67AeoR4RX2iFue5LcFNZJcpHBq7cIz+v7dnw5Ha3/+hoKRcWEU4U
3r60O/S9QJnAdiffTroDv7b92mSUarvQr82kYHK+l1cm17cOWSYzxLfK3XpxIHWJNgBKcOnCsl86
amC9jxdpkQGEqJn8lIJCx6OSkvJ1Bih1/JIbTYDiZ4uIKDDw4WwxlU+8k4KAA7ZUtIvR5aKUSD6r
+LvbGtUzfMEsTDD5KQp0ZpwQpEt15t2622rUd9NLfNFRHRdvhicXSIK/4HODDb/kmKthn2b/jXzy
6SkQZEKBgZGwGtYzIQovuoOwaH+d97n96fQRUdT2gvtwTjMR2yVz1SIGnrTD4kC3/bgEEGzsygHK
gE8lC7CoQDqI2slvnzDvWWiyehkCUvfqwjyHq62J2cZ1VajjPDeW04uBhsYhnOfI0pRFPCqaht7p
8CV7HduMtAi09OmgGqpkgli5aUM4fPSBI3LYK8DgUHemVO3k5DP9UWUSZO5Rgbsbbjg/xQp7cu4V
R0pAxovD9N75w10odPHgoo8WiUkMf3OJ24zWU95Aj2UobVIbNHfzIecok1CPvCzER2aO8PUr2036
K/qUbcg2kYy8uN3iPlRjz9kG2mUQ8i3BShfjRQ2/kScLFmq9FjgHosPUKPMtlUWncEXjX/Spomuf
sheJndTY5abHFvCx5K7wf0fnvcknIi89/BUPWHiSwfc62WVP8YT1aJjMzCHIM63OFtuBHXhzL9cq
r21ZUYDwM6PzV23rmlgzZcFGW/6jZEvnn0aZ432ToZOOb/ikHVOOk6TvQ8/vHpvMFPrCaPFwL54p
QnkbyCiBZMj0SOo80qU4LJLUyKSAPZBAieNauzKWOL+LuWuZs6jLd6bweBh47rpOnmTfy+6h3hb1
+QM4qy/YmvXisenlRTH/KMu1fYlcZfGYsIbm1Ocev+ujKiuh73lFIZLNJb3roqvbkoXRKo9aHHVs
GVJ9D/AcSpPLpHEBSdZWMamQ5CZ2XBApW1v9icclA5lnd54ljGNkyui92tWtZfO5/J58iwFZs1Hl
H9Zi8coN/Vaunqsv/q9a69DG0N6FInsCR2xktlFRXl6KKR0KC+oVADKEGpqB7mJw4iqg0y8txllQ
Y+MXGQwSI3DpvJvZMmAMnWNzIB4MPknjchLgFixZo8CB7q3bQGDBTghg1id3mVjoSx7YAv8T5ukU
2nMwFxzPLaNhuCjj+K4QP3nGdcBIRgeZwEDvasJzS2lNE6KJ+tv8t45KZj6MBx9A6nyIgBQAj47i
KFhvp+tvxDnzEMquwArt+boBAEncrqv3N1/OhmTWNkbJ1u+oe6BOhjWyVjgUNZG6OZtWRTCkk3sS
ZE/EUGCetu5adozAkS5vbvBnAfhQgmBE/egq4Ue2hQJ1u77+L0PtfdeaLfH+A4RXrAavQzku9OWl
IESLK4ioY12h4X/reZZZnI4ATzX347kPmidlnjKdeHQL/nFoc1gMwhj6vfPRqjgkfrZBj/54q/yD
7z6N1+AMRsutU6RrX2IJR/vdUvuGYdB6GLGi3+h8Qhl08mvZiLWRhK5WzI/TFLZjcEmh8iavNRsR
3pQohelamlXHiYxsf5bE7aIT5zqEQs9bfy58vq50IRPjDt9gcvlNRNuRClLPzkYWGkygEJ/ympk+
w1ghePXuF1PVaDsauAEOff/6sBkPeXd0DqB5L6XnWacfNapefra0WQ6cz0iEH1Q4PS/wlzkAT9lb
gNSTJHDLX6MsRsS7JaIf6W9GaPDIHPPxczt7HvZY96qsmXYtOb+5lpNOWFBNiUCFf9cp1WBya5fD
Dyhuw47FI7RsgUsfEhk9EGpsI0tE1GkgwbSIjZaLwiRvThmTxP0AIlpEvig7dWYr6OzG3750eQmq
2BIxlGpN9rMrImBC1TGMe5PBp2XN8EpyRQG71YvTzD3CLTMQ0RecWJkqkvROp5s5AtStk13cjFKG
HRsALETseMDuUeW7N0iOPJbVxk+EvcFoPxG2aNgGQ8CUDLEQOZavqgvHHK2tRUPd3dyu12ADA9Ne
5Juf4MVEz38ImxtZfuuE4NuF0F7A3PVwFpRbUXXIQ8U3/q0LtbzTV1VeBnIB7VqSahQkWPZp2/vN
DfZHquU+KL/7W5q4jLfX7b1lsYeXX1WEHuiWKS1/9ppgzbkAOTf45tRDPcFM2tIqgiKVs/4uqqxg
r9j8uMJcj7nHK70XDZd0uV3TOufRwRXe5PQj+oI/INMyibh6mWRPFS6Jv9R72b0oM0qugoPLd+fC
aDtbfLXsl1KQJiJi0xPI1CmNsJodWSqyEi2bI1+7RXwQUQ0wXvPkUfOWvHE9UM/VK08UfeU8DaKy
r7o11K3csDfxaOGeE5GrcJVHfi7dVvZI2G/pOQ/5qKd8SRQUAC8flCED3pCOJgKnCEJ91ZDQAPzS
r7cEqng/eE40i38boqp53vyMzH/T0KYGrQFN3ZFr7pC3LSNEEtQB8ZYgcnfFLU44YJNdzx0B6Fke
zdNCGJejFQj20J6+jXB3BhGPyW6x9xQEHwgMoM4lxW8a3oJzeY/pkl/pQpng89HDbgGWA3tGv4X3
dPVcCwiPBQUCX0T9OzeAchzjKypSJVvM+lTEtAlHKLGRLH6MFeA2SGosO/pV/yhyEy3G+vmiN+YX
wgLFDEVvo2iXbExYk9k0WFdVWt1Z58v/4AUKSjXgmrOPqQin+DILMrWklHEEc3XAoghM7tV8oMoz
VjCXA0BVCV8+kUJMKb39C3UOBboXEnecXeyZNbn5bstwwafzLLQ/Lq5hLom7YPrHIEvxvSb27HMk
7GLTzf1IjTMv45Q2PIzGX3+fG5nVvfoO1exGI+FBQMo2r8Nc9Y61r2omTt8Xa15MkgVHxvWlRiUE
xkmG+00XXLCroxUEPWPBkG5Iaz3hU5QmULbb7w7vr1liRNkJUFgR9rcKlJq5dao6Rrh4uAgINxs/
+9UHEqXMRlUkzRYy4rokcducTPEDu4Kzq5gIG+GWmEM3yY7jQetZHIxzjBTtkxSlxOqTLRRASfCX
GR/eLNBYqegqhifZ2TPI6Qz+kFLqmPCf5kn9V1gGJpBGOeIkoTNx6oCrSVmtQNzzHvCp+lkH85jh
Na4Fc0B/W8YAdfMCKr9+DeE1mf5g7Gs32+6t4aqinPVsuAGZ5UjkamxlA4GtlI14XYFvVM5r2W1u
92LcCowq1wvIqJ5Onodv1AJNN/I7QJ5qf5WAKewZThsBcp/M8uYwIt5Q2QlhxMoZSi7RVc6N5q6R
BQPiJ0L/oT0tqnnPZBxnqmbx4bLUFRmyL6Za6o/0P5CVbQPDc87jPlXGoGuOYXBb2JLbSv1uZ4ae
5X9WDnlinnzl+XbMCXMbvOb++DMzdEjydnid+F7CC+dImqQWvf2/wk2/SyFtFOWpcPWY/nq8TZwM
Xa/DwGADfZGws96+P8LRr4C9lBn0avib3pnUy0FLTabquIXKLSCroKvuRGYhEfdHWtOboFB9+JFG
6Kh5lImebVbEt6fBQSriCOXkGxamAFQfq+RMH4zRJCExUIZENF5fGjoZeVDj/ufr7QOouYiLBZUu
Q4jTlYMPfoRwKwoqbEDbLnMxJsa18sDq9qRm+8HmPD1WgOz0Reid58nQrFLZKKYVcgq2C+b5Fj16
OaIZ2s7xUMUxHvay5ym65OpkS2HfY4ZJr73hRzxF3iiOROKs27f86oFI1pd5tiSxBDkDHc9KKomA
QPSkDqc0EfGGI7od0aR8D07yxGuNaSqZLV9ZxXqEzPqK6P/pwozLfnE5o+GjCO3VIZYMRFvxwuBj
ZQHMiH0BLY6LFILQkPd92W2xOQeZ2Bj3l0/xJfR9xdr4rcsgGi2OdGbRyaiOuT8glpvecvXY2IDu
Zqe05gqJh1BJLrOrr+gH6ooAV/ADRm+orZvV3QKnoivjbRAqvy1BtNqtpQFYw58QtWtfZ6iHsAm2
a130gI2S28x0KuS49OWt3sZBiOJV6DYf9lEHB0kEiH6j8YsDOUIifCYrjKGnDXd1RkQ8b9Hr+YPq
sQxdfGKwv53Q933gYhbxhzxEkLh0QT4T1NsNBH+qojLRbRBeX2pbqlNEY9MJGKMJue2f36cgf5rZ
X5GzuON0Y2mXepxmNKop9DU47NFRjJDmWTuO/Oy4gElUclxoiixLeGA9PhEmNk2vZEb3WC1dy7R5
62PqTrdyOCC+vzeM61eicITPycF84HyRgeQmF05KzeZlkKaILV5Ta/WaeFSYFzCpLwfniJZKCa7Z
ANQavUxL3vdS23ohhzasfXOfoN8GAj4hzkVBrcTfnsLM6WgEkUsiaiorNSeuZ+b79iwHgVuYulMH
dVFmQUsB4qdpJKTYYSK88zvYucrJvere1AlAQpqc8GvkHkq6ZJQDWf41F6a4ijHMyrq9fRrT0osu
+Y6pdVNGmHZc06iiTij3xyOrGZKCgpxcaxm8kk/rrC68ed9G/bxKOdEdh3JO+yJ497zz2/stxh50
9U22Z3GkTojYZIL9VZg5UdNNm+KHpSKf9JRX19eeFyTSmYLtVEwB7BsfIMVvUO/3W3YH6GGiq/Gc
VS30FFpt8dh+zMe8c9xmxjste1DDWTWUoceAKRIdSuO0afg6M+6gKtxk3meNZTA7pMhJcaK/VXYR
Po12DnZWFzrop0koB4SW/PP8WkdY9hJy1qJJIo4d9xqH3k1O30gdmBcivrqT4Z/w8R+E+QaX4wpn
yjH/mMiTV4JuamIMjC2VPj7pP0DuWzFdt9dun82Itz0GWrdO4BzV/PHygiXZ4hTbVLJyFTiJxeQP
0HOfgN9AaXVSEeFCbnvHakCNoe3QeDwjb/NHPLkuwxkQgsl0/AH/TKcJVN5i2so8uEeNRQKkG03A
DedxKJJK2wdWkwIEH1vVjpwHK7OtSWhNujqtBeK4Z6wlYMQmTJgj2/maDt+FCjea9XE9JyR47uQM
j2qkbtOAO0Xwq/9okKOfVHbMlKBoH3xfytzDye1W3naDiGY69akEeU/cPnKn2XrB9BQilfdrflL1
63CSP/3lArq/43SC5AWK5DCklmFheuNJpE9c0thdYBf4+D67/t4cXAxppuXSeWDExaK1k00jqnnh
ILKF6AY/YNUokuSZjVf5OluGeOa0khlbu+H8BN2/YMt1uZfOKr08oRNHb2yl5DvYKoMkabyfOEle
klbz7921rDW+UIVwtcf+GPIB/bs6zdPW/yRnwnivesV1SE7XI03WEsIPqZZV0hZs16T4FPzlQk/D
F85FUUQyWAha8RyQV44sX+nh6AFm2bBuqNTpqlmCgilaVH0zRAYbjTQ0WMcMIZ+cErrtpudPcEUC
V0kqD95sFuwSecUh8kFb0ZWNcESMb1/JKF7ttX7Q2ILCU9/pwdkB/g3r72PHLQhE4Y2Cm2DSQ83K
5+Jh/y2Hy31XkmI/3PVpqi3DQXsf4SO+oLf5zvk7tr7E6ZhPkHzYrhovQRZe/arlWh8psivBpxNn
IxGUf+9A6dZEL+sdv4+jfqIAfQo49EohKnbhuz2z8hi99g2r+nYxKbntjlzTMSpmNbfAWMLRjf9g
tAVAzU/UINVVGE7ICL7U47aMiWcwDG67lT0MA7NlsYpba7/iD8xXpsEp7u1pPR7kJrPjCnJOKfmG
nV/YH+0/KA6R+K44Wm/bfAQsJsrpfG/brxvQqMr9uAnAj8HeBF8OvWvskhTWCZCkE1FkaUpNZrV4
4h1LcN7RMj/v04S7/dHlojYriC4uXup9UcToz/0Lg3IG62V1Vyzg4OpwoYAxVqEK69lrdTWKA03T
pcJl60SOQQ3U0DtBVrrT6zqNTpDcfgHNcnXuHT0EPPBsKwcvrL7RH2IiTaYvKpEpzZCECSlSLSDc
EPuxTcwEPjnXkQe8h/Dc5+atjNpWwCbPOJXNUFvWEpOnyd3+NbqRFPgEC94kBclLbEHb62yQ/pu5
c/Uo+El5OHUrunUxYulfOfB2bNM/I6UjXLmNAD8nH8tgWDYDAvKnGWC5QN5eFfx6d4MI7zvLNk9C
uZlEZlL8hSQB+/qfeVJPQAEybv5XwujY2fJUzIq1Fy8xDlHtcjUpqV6mS6QYGBpIJw7i98mTTujv
xwQysAgqkrr7nQ2/FVAUm1AF+tl8qp6SNBymxbfa1WiU4PK9l9oPo2VyDOPPDAaRgtoNu78x4lNI
HYPxIkaoafkttN3IkltJDAw7a26ziP5M7Kk0taps6AKvVcPFEC09P1tjKfab0d8auhxyFpKTaNPI
5CsSaXozjTLRG2QwRRvhBln4mfwDIIPzPJJ4okRBV7IlpYZza1bhGdaGz1pfHTYttXvXgi3Dwe11
OuJV6Zt9g83OK2R7lwtyNfDsjJPdlBVA/MEDN0fAXo7WnkINLLkbgVd0G3yxiJycCg3SyywNg494
jUaT64fo3OkKiEP+NRLVnXIX31n9YrD/PYm/JgtV1gklrqjWQHliTZ4u+ZWHfRpWe0r6qs2SRKqt
kJZIDxCC4E/ilEy/S/XwCgFQeRGxRuR2x5MxrZEngTq2eBJHEhvEwSpF0I6JKZObVgywB3OMArrN
+VarWLm/VVyZYOWa6EmfJgG6GpFQFU/xJitK7vg9icL9ynPRcP0zFtyKmJiD7IG4ibEf9VfWsbH5
hdmFPFhhJP/E1Q2faDRzcND9wt5QXRuz/KIa/Khp0nVJ/u02ul4l3xe1AxeFi+Zn2Vmovubr4c0C
VGRaxtMh/dZ0CnuZQW9O/JzKkvAElmkaKLXQU/r4rh+A/FiwYxTULmAw5S6prDFkFQQPLqmoPvv4
KnOncFtgCmlTLi4oqmyLBcn8lvpwYVs8OvccgcDwv06qiesFCyTnaoVNeou5PKxgHbsbKQIcsGXI
w3oxLbba96C7T4jr7ie23XWpDbf50U12Mq3DdZGPFO38W7ZTs31cGslaTmwu+ukm6Y4KF6bKWapA
Jg0/PtmVX6hE15FoNAPxtfowYEhLQlg7N25WFH9cpIeILhpKhFsocjbBADy7qVihtg0/u9Ejg9Gu
J8GBR+7Cz3ELOY2gnflkFgu3afFI5e4GdzOI5Tmal+7ocMAiDAufPlaYYQOxLMIYnq3pb2SYtoTd
AT9X/pbcR9vB/VE7igrmDHptv2OdXP/PeJkv577ABv23aF4f1bRgMOHSmhZgedM3tD44hFz5i1k3
eO3InhV4iG79R4HMMe1OpIB+Dprd0PkjYTJCm7HuKY6Ja0/6wJ1qAlcYdWoXqr+BLAoDZFTim48h
rNkQvIlwx39BhoicARPOPX9H5eHBuRodzv6Jc+fPcs9uJ2YcYbnI9tbsL1ZoYSKALWQAzxeukf/z
pqjaZQR6uTmyZJ95vxYbTwE3dVWkL9jG//Nf9Vch7G5ibKghYkFYqBq8CpnSqnN253UGhmv0WM8/
r247B4UcCZV2fhghswEHmvRoUt5xWa06NsS9Ue4OOR353RvzByHqCKZV1B9BDznk2RQ2cLES7Zbs
dTzsMcnpzA/Mtl6sraTFua4z1bAb+U5gkN0c3x1hnag70yZoh7vJngi5Re+SCCgttRBlfpzxr2GN
MvlLST4kvWlEsmlVYClvp9oybCP2TebmwHWeaQVm7YFL5J23QueIx8lDzFDyDCYT8hzvPVlsDxTR
vcSA4xDzY4KUuM2rmVYZrIhTTMgHvvaoiDV6NH9kds/DsMrt3LVNYJiV6A4FIxSLc9B1ZLDZ746/
RTBZX+LPuyN5APfrOXugaUWmmz1aKlesjUgaevnHlqH8P2a3mLjhkWbZG2jcmApI9EJqR6WLM4Fu
hF2MgoSzRMUSmyZ8Ywzyzmtlfk7APmriLOXKSC/7fIZ9TL2AalP4r3T0xSpDJ5oL3uXBREct2l9s
NUT2iDwVq87jzhOZSmbjMPJ41SFAp7AxWvPfdAJfR2A5R0dYJe37eN7M2lIlUBIiGVLYT00xSS/8
Nq7y36WDMefKD9n3Ia1q9E/Q8w6/uXQoPLaRaCf9Qz0cYOuk2FGLGxowMzsT8By7IFQQaWdH+Ixl
kaoDiBQXMS639b1fsX1biVfvx43RA1whDs6q31AZl6wiP2XmEkgpzYizKSFj3SSdxzwV5ESgHsEC
qKoicMRtwOpQUtrOtGIRWADcIk19VDa396+pz2g7W90In/n3XFYdptLvtHb58082eFLvahWp8g1Q
nGyqy1sKFRqtY+JK8ygo84xdNr5rAGK1YK4ZdJRawt/sI5broCCOBMJHga+m1c13doZ9rdSh8EQG
hcmzePbvL487SQzhnIV2+Trx+mN1iO32X7toC8yVIBp5e60xAKBvVnOSBpE8rqV6PtQFVjPttWVy
UnwRZ8oXiFjRS8u6wjJNLsGPiwpr9gngNlkXc9loIcYlZASDTfS9qo0zSqrNsdPZr+hv6IccwVtQ
1NWEWWrbVD1NNABSjqhqNeUEQS7V2pgl4ZFF40mXp4X2Ob3uuoX0YUiCEUMsxdahwVnbV9F99xF3
yyb5iU8ZODduzEgy1YSAkoqUFN5wD13f/ckEymZ1g886FTFBDdUAGi2a6d2dFQA9rmD9g3yS8xeG
BB26xZEIsVdGfTMO1pN492G6KHQ3yBywNNEw6yTmjlseSkleRT+E3X7JF8rHrdEeL3R6Nupa2qv5
EseBtc9j2T3J4iTyigE339pmQnhnZptLcWka+Kx5vbck+yV/bsK/+YplttYAx4G/k9UA61LKe2d9
1aXYQhzc5o6FXjVk7Ke56+zp9FXX4cBgg2TtCW+NykBL/vJPxRtWsbZIa2VT0rGQhLAGpi98X94B
frhQsaVNgSVOXzHRa/UgKNlGwCkVHsy/jqvR/yrBG+9Q2xm0c5h89LWYgB/hseWWmdMvFXNyU3kN
JB3WkRfRUgsKwibo0hSWsl8LE6BronHOFP2gyvO8zg7by+Ge2j/W95Li+yiZafoPd9KottQFzERs
lO2ufJbKIjBV0mqAilitSKgygBkS2NHovuhenwouGRJqwJ5PrSzURm1BhaV6OIZ8n8FiAF8bpiUW
QAEi8tJMkXTEh3IlmjuIhYSFhy7q47GLpXsPkHzDA1GNYuF6ouHY54yWvWBxmGjc15T/7EKKI8Q+
47IPdxwW2SFJBEI/WY0nSJyYg4QFig7JAMwDwcnNHSmeGKupIDlkxhJRp3iIrqQHkPWRHPRQpQ5H
KpLyS7fZpjrb/CKnk0fAIyRmdZgrEbo6OjCrCwUZ6DspBE5lUW1FWq/nnSFYWvVHSACWPznJz76A
e20FFkC24BwEfcwyir0C9kvG44pBTrP1CMUKI9yd0/C5+WRcOc/WynqjjQwaRztgdNWa70nqTIfC
fwuz6Hk9onmn0UiHBD1vpjO2/LRpTPjM9C/XNdAcO/iNeqKB3j+AfVI+GRSChK7bd1bT0NG/Z4xn
pb01EUTopYskTBvgZgfPwVFJJpxN6hd6yYF3h+KwXSE6OjL+NV/8BOokay7JiY5U8+f1XGBpsniE
bmyUOvfSut1x7Py4+qwmBBLhu+otTdPvqYeu1ff7DMZCcTSD4hhVr8EtJVPbuaLP2nFmBJMdTR7p
jMG8h8wcMcEUjG93IrSJxl0HQQGl4/Xv1+7U0L6lU1TRiJTlLDAxq6G1gUUVxbJzB+mX0ehLBFeB
8Ea+ud+TsUGmv7Sla5N0w2hxz/7irkfxqtPTMutqXmIuIl25Qjq/XlWfxy28+fFqUrNyhCNtRGvv
rmzRt1MtueNJwtzO/U8EF0HSYkJh5TGgIs1xMja27zo08nZ1CNtxoahbeAz9JwF/5rl1yayWAWQO
XMEv+FGYuPPNSGDneJIFlBAUc0wwDwyKWfRxLwkIVY9hrdP/aaJP+3dkmlypDUvGqeESQgGqXXPY
rUMj1/47m/yC5NuPyIKJqB0DpuUxxAXqOEOGrehy4AOIehwZ5UKectTyGn7CyV5M03Jg1dvzuQBg
M6KMVKhx8f+eZ8pR4ywhx+NDjafrWJL0UVj/KQw8bqZXVzYEDvQ6lNmgpzxpOf+WlTNAYYMKXnCC
P2wXF3I894zmek4pH2my9lTsUsX46vifBgxaa4Cz37g8YcDx+gZhg9mcEg7/hm2Da4kMvhTFaLO7
kfbeAlor+4TYYAq2P76ZI2UQJo2zDwFdedg4imTgdWAg4MNtxGPE76fgGYyyimp/Aa67JTbcyiNf
1WEoPXIv8cTFiiiyRc7hsTBQMRsUpjiHLv0gww6bBwKS+OuT8RnJy+NPrp9AocC7jBEvs/2kaSke
yabHtTKkScJfJprN07eDFLPBChqlWB7Zm1SK9V/XC+91gviT8Hh1NDjSd/RQhWe++/k7bS5m3Fu+
pBQZosPyjoyBereEfdsamC/jqdX9t6M4jUmTKEAraBvyqke/SIeU+Z7kuGUKsutLKEiifkDGxHsM
JVvCGSQeOPXjz0/95V35av1jskMedvHxmS8d6QZmTZewTlvWSuHb7pfgJlft83voXPX58GM5HUAS
Pu+xazK9xfuKhZqUAeVa3VlpUxGPCTJcmvk+kRpOLA82f0Lu0jZ6IKPXOaYhRAJf3gR/QI45RJq5
9+G1r0tTtaD2a8136j3loo+Fm6XtlV92tYzilLG4+l3qYIgLWGaCwX6ABXC0wdBsUOx0nbaTfVf5
xF7yxanew/JfbveYNOgJtXFPJB4b5IS0yrbm53KUwQgSQ1wSpJq7whioWZY8ZF+6BnNIaNhdLq0k
owe0TXhHK1HbQ20825tSKwUhLj+yKIQKV8ZOKCgCWmIc7yDBrfXyWTAatoic/+keeepfNADoI+Gy
8jSIrk2lrSPjMw+JxmVFQGrq606znhaTFOMAG95oR0lOkON2AZLETM7BsO5zpZ23ixkKJSP5NsQD
jz9cv0HR+W4QM/d3smKjdpXRqTbx6HsA1Z6/Y4V63B1C0/XMu+YG4yo6eJ5cNafUms8itHfxxYHr
38Q0r6SAJO8einTilM7z2P84iYSRFCJBZX9vHiYrtRbVWlI4x6UvYLSJpdNngrB9g6vgyi1rZcx/
LkB83zqfMLGglx7v25ojHdLkN/OzxMur2+7voWjnAjsqmH+t/+RiOA7+H7umXefbNc/erOhra1jj
JVmvVcky8Z/cT5L+gskuBKTemCbNStXUYrCwU01DNrVkwBXtTQw1t2gnjk+PqKAZTJM51F2n+Ga9
FaZwT6aKs2pc0aML1lo1MV3Ptn0mDNtnBbTzpMgLEIs6Y7TnXkUbCcm6eZTzboZ1E4Rdm3jglh5R
+3nw/uUCc6Hv99iNky7nfN3+tlx89l3F10yxlUbQdoDjetKCZw2HJiGTMIw0fw0G/lYoy06HOf2C
rdbgaOKmtKzZcSQ6UJNwb9Cwuw6pSHQgnC3wnQxxDAL8mBZMuNlydutIrCp/7ZN0jxBva5rojOKJ
b7ayRHJ618keiZ1Ex23Y7BNVFG66tbvNOTVEloBwibGx7VBc3cJwCNLR/yTAVpPoI4MlZrcAxPpV
/k7WB+ggrBeRVHlou/1WY2WviQpdjj1RXmpRQ3XKPNVC9nxg6H3TfRu+MNFytPfQwB4g/xMYU6wf
NN1NZFi9IJllGdzInd2cpXLvldIZl2I79YBEACmE8f05I3fckcV1TAdhGo1efwHnuXOw4AAHk3jt
RpUrjL218gjuzSaV9hgH4sBxXZUSk1h6noZovYyDgBAWVbpe56n2BvvAzcH4nG8vTRr6yH5xck5Q
/8P8mfMqNh+2P4bfswEqy4f81VedeLmEu3qU56MoDe+z/AA2tEy0FQOyyVOTlow3VTZmeiZvNtpp
KnHx6mf7PJ0NqBeWJVp7z/BKWGq7ETdicpI6ri6FzalpDP6BVJBhc+y+uCtmyfQa52Y42WEXt95q
oG/h/fsw8Bmvq8YpWcRFNwslja1EZH23qrZMKeoiNjrM5zyzmr0HQ0jr7qZ/hmprNBC09z247Jpx
Jy/tRAOYOxIWlARvNfJyyTOfg4pmaG+RsXzkQ16N09hDp4ZxxTL9tmqbAAxPzXkzDPA03eEb9xQO
QcCAwr3aK+DXgxDXug1wvjkrGmimz37dT5zJf3izh5Chquvx4Soy3XsaxLBuFNnUIyupkPFKN7mA
uADzgzeNB4y3/UxRJmbMoXSfU/s+IjPjnthnKq/FXkYf5+8+UncfHDxaNaCbwx7LZiP4Ab73Uu7Z
lJPxdKKgvrzfvIIWnnORKZQ2cvoKiVzCZEDO+SRGJELFDyjEvftyhHU1PZaIFxEb05kVARVRHgnl
lOgYGlYJkaRCeA9tbSZjDw94stiStqvq4rO+JSXlqOzazo5+Sm1G5r25GTpo0qBIa3Ar6Iz0kpr5
srpjAyfx1MzMB//WKMWE9a69/nYeb8v5z2GN/H/aivS0hZuQ0JbzvNoawbp49Pa9eR9ku+lvW6Mj
834PotekMS0HmObMnJQFf08zPJE0U9yHLmNxV00WV6bx2sVxtNDEtKwKD4JAMU0TmNJij1HZa62w
l9Ho56MdaM28im1vH7P5d1orC7zVeO0alzZaDVcrZ3MM4bML/jTa7yuy453AkgBtNzWzFgvivyJS
O+JziLd0wRUpe01Yp5swUR/FWRhnqgVrWwW54qm5+ch48rAq07cqjI+F4xmybJc7jzFah1Iu29/a
dlNF+EjePolnoJ1vVneKjhHwl07QMmtdEBVayzfD7oeMzmkQxv65II4xKl+AjtIVb1gbVryfX2Nt
EluBYi6l0E7ikwzX92LAqRIiI4LViSmw4A3TAquoD+u2I+nqE4ey/hg4KLEb8WaxqVgNQ8htGowc
28sH81Vsn+siNrRDovqocRr1EzAbM3N6Ye8df1LZEC9zmx1adGPRcNXbVmRl+Y2b2upCkgD4m09L
zIJsoGWbnh/XQC+xMzB3rFrxpD5l35dwRxWhdiHyofx0usMqqPSFGmVZORqKhPS/d8O6ff2/tkCg
t1uEgsmagv5VUm1c/DSnsu7TnC7tufH1qPvl1KCVoaYNSs1Owg33ipeET19KFBAJ9KGeVaQeYOX7
vIETPGkWcbp9Peb1lWt/o8Ydd+rT64ZJl9Hihjrhv7fjiThAEcb/C2DqQk8XFB5OVXvQsqq59InL
afYM+Cs24Fr74PntJqwU9jDHoKxddjK1X5o+Qln6Mftgl6A8fNO7VJ8QKEbECuzj04LTGG42IP3O
46eJG7qRJKW58hkdB7X3PF2+dbvO5DKfXKZ2hvUMjyTIMsX7e9CC4r5rx/62hpMoYcvjzI9POX+k
F9bzuayCGn3zkNVkOGJWTtXE4ke212O2yqf8g/hyLZOxedyt89AaowqIsMcIDH5Mx1vMqwO7wBxN
+LMaryNZze1OxNzY3+y06xfyHymDHOu7l/e1HH6SWzYBj0v6HDyedcA8trd8Q6ZzPRkrClIrs2T2
HcJeWT9iN8xKaO97FeTCkDs1wveyYHH5zEeuVemfk6Re0GIb3HJH6Q6QGLOPVMwpgxbTOWyp7Edl
U6xo8gnHxGwTY4x+j4kIE52OuSKXfRSZpPCpNCUtvs8AQ4uIQCbaszjL7wKjA6zvdMROKVh9bs3C
Ljxz/F977FnaA/fADiP8xD5VYM+HetZa7VH+UbLMNdv32N9YkmOh9ns2C6q1X3+tBP23vH2HzccU
BIzP3elWRRpT1jKU2LSvvR7ioil1yVoYNT7AbvWiXnV4hmQ3L524qvfUrhbZObxSyEQsYRnYmuSI
8dvYiD7ZhQxBsBOfJlDQ4Hp5T7PE3ftO/EL3YUHZPhjqDl4YereOWvjMLxk54Pu1fDhKslbsfj98
kZ1Yo+TCnxS0JXqU3sDV2R9qe/zhTfvuHCAVbVhqYLsEKraIQkKY+5jCvJfRT3yQT2ynmuZSKpV0
orxpoN6qvlC/vS/ewej3Bm1fr97FNeIer8aGZv1a0HQQxrAEJtQ9xfR8FMkkQHQEmzZARBYF3pVM
A1NWYUctf+oEk9pcCTJVp1WYWpAuomCVuNRfN1tMHIjjxM48/5g7srvRqfwte5Hn5ZS5LgDzwieZ
262JTVQOVw7NeKKpYSg0mf6EVe23uFx5gwQ0MUr7dm/Urk2z2qihr7NSw5zDd92DITuC5FA8hiCj
A5CsNmXXZ5Y1+a2N/f6r60l4jzQwhflxdQ/sRUwjbvIrBqoACY8yT6T2VLiU70dIMQNyOpzZSalH
+yBLDb9IZYgbz2fv9RqnUlBw153PkRD2GFhgw5X++k2wPLua6Jiplhh/oc08qWAIAkhvVv3bZUrg
pqQ+KHmv6e1jmnG6zgV8q1OOLcy0rNxujcuBHnMYtkXPUyLbKfBF5fmJbhXjTF+5AQBPeDpmBDcg
bpAVLUVwZGmumUG59vLycDZ2Rn5f57RSmeWWqdjNdRHOTjo8VnF98PDGupm0I1ZWFTQvDajHIBW4
TPYyUUiQDasENmTa535NElD7LD0JdRnZjvFAdzooHc+/ljy55puOZ5X5xM/XCWyd248UVuICZcFI
0/Jj7wWpHupJVIMrXf7z+peDoppePWl/4D4USnV07uAbLAHjUn/1cPAG6o5SmvoCiOQK9jjmefvt
iFfO1iOH5h/g4xn+yeLCUNLhADbBB7hhLB9tYGpuD7G5gi+9yU5bq8ZzEweUpithKjMyKKtxMS/j
14Fg/Ves3Ib+og5SaUMLruBOqdc388mhjsXfrEluQRVGdZavBtDoALkq0BuDMykcBiCN0fXtHk8S
UcWVthmK+uy6Rt8SKpiwt+aG9cbVso/Vcoplvl7mY4EuibydAy5R+EwCJllN5DWG66ugMu8uGCzj
fVJBP65YFijeqsQAt68fI2mloB0ewEGT82b0dc8OrU+Tui+4IUrsMVifs42ylLCHry8dd/2IkuFt
u112VPuDeMOoqsS6uR350KKsKCxp+kt/pnd12YK4KuY6YyHb5atsfeeUnt5ZIS+wXM1VR93xUL+M
YdrsOa9E3jAdhGI2i2C7X7uVYMljqKU/ARE2ND1CNtEdn6wdrsl0xM+m5DfCPJcKXqSe5gx1mcJW
pB4VEZBCUYpbelGTcUEPFxyqW7C8fd93NkV4X3LWLBEqL3P467ybl7XdbzUI/bHZUOn1eqQd9FDq
m2xAdnmGNx9l/eVHvPhODQMaJQcDwuaBa2PMhO84xeijsfzVoAaRSNh61vaqavaj+zhlRXHIfdSH
2PnW/aKprKF75IM13aPBWBw/nguwsQlTxIniMt3mxjYXlfViMuEIKAfx1uNftCI2B5qK4R76kFJZ
qAc1WNT3xYfJDR0XjWFF1iSU7iOOQaJF2SgyKKL22qNIIUwbhiAzekQGCopUklY8RikyPTMfqh2S
BdXaDAAb2VWAjkd/RiFGlSNbARbH27pUOqYRA3CRMEGPloqrDcWsf9Dn4x80tg5Gu9nfPMNhlDzq
d4gWk4gW99HexvCoP2F0lAusxoD76xZY3xqIyuaOzqbB96t3VzYWdn60up+Zh7giRecK3ze4sVPt
naRzMjr6elPXxfuJW/HqoMzAdX7/yUfI1V9jKoyKQvkr6TmpNPcD2tIBROH2/cbkW1XaSvTKE19W
nh0+rPLIj8cHbiTqq0MWjhU3VXe/pBdXziFAzsnzQSd7pz1ly4ddLkVO04wb7a8gAea8AetxDpUp
XWS0FBIQrXHoNVtn+R7/O4LAfPVR2pkYuxHClRBNKm9+fZQaB1K2yAe+3EscreL5XWfqSjW/MzzX
is570zXNz6BdnXKxXXRBDnmVEztYYwMw1hyKnzLE+JkZqW0H0syidF1i5mIWllRhJCogWY1G00Wi
tVIGMPTXACGseDH2GT2gxXFgOZQVxv1Fr+TzJ21VTGrReJ2HUKgN05v/DUNcfc6ERFrDV+fCNqm6
FJqimpsBQgbwg3e2cqVTKoRzbe0AVWTlfHChFjXQjmaqGPsyZ4sju6fi2EfeEgZzC3d2zthZsqjY
OuG7vl8NUz1d0dbiotRZ8sCKLCekrh8T7htwxvwT+vTEUfDOfWdvqUuTiDjMt7dnCgoh3/3XUkAs
LJEPAh6SVDQc5oHFWlisUaLSCPIewu4x6O/i4cRztvmrg1mDKiLKNyBNHshTjCgDd0RgS4dFat+O
9Q+nMTG76orMSVjlzmCUIHry7M9agcCU5KUx9GU52EU3TBNKnX/kwfpZLan9TkSoG0EeFIsafqxz
P81TtuivOodjt5onFr6KKXUmUd/p8tNJDqhkTlw77lflx8pWWVoBxtBFFLKXIxZTc2kCOdpulEps
swULR8/6Ac/pLBRCK7+hZQZ7B/Kai2N/OJ0+QqqPI6eAe3uQpTKMsDxXCGmRVGovCSiYmTMZhQEr
Ag0iav05UC76ym6ls0V1TBLxlYyOY+nIBXdFrAbMzKen/7qxd7tt3hbIJTQQiNhELDg/NKwzzHji
E0SYtJ1K5Pjub5huT3kGQJC9OUM7gynlHi3nKNNi/3DNGaWDinQamcKD1aq27qtMdCRwSSHT7CGM
5hRwf+Z7r7frYk2X5w5B1TVGzc2NMUcIJm7j+417frSleBfjSUlNKKsLwdcuUFcd3XcvqWVrT0tF
Yc+uF6/yV+ku/RDN7yCzW2kG7mi3Xi7wb7p2jecRH5NQuBouqr1uafrBSeZmOp9hwu8tTEyjBjth
B2erDuvbgbQn5sr/lMxwp6sckBThi3YvaSMt+1AnJ/E8/HsxV4BrsAWlFHpZNxXGggpSBNY2Xwrt
O6CPRjCIbFSAAmNndltzfaMIkWjgEURF0JDarUOSlBBnrKa5YyTxGvtQ6HfN7NoUqkyFvSYzpG+K
MkpqYjY62HsY7LpLfIpzVSUwuZSCgHHGBvUYXk++jYhxARCLo+kB09dWa9XnVgWRDLshw+9c+lpG
NcTCz45ae+8xQTFD0p0IfsYKGHA4CsY4UFFDmhJuThmpB2hNfipvWb45KM7k8aUyerT4a2TvvulO
2FORKcaBLiwnL5lYtc+xs1girnJPMxbde9Rk8Y20mGOFCpPpEPuHBE6ZyJ26jmrO92I2DYd6gWMg
PwAfmLds2+7wLwD86/jzfS7yPvR7sgQux6OLsjlen6HgpueS6/ZFxwQkjWnYftl1kF0fGgGoox2x
luXJAqYisYz65n7UwNC0x220L95wcthZRLv5aKvv7fTdYfU7tAdyFw9rT0zn7pu61Vb1KvR7RJfv
SiVLcFfLzhdMR11A6bHcA9nmBVhf7oGhEgOdWgESvyU5SL4dM+kYg4jFtljnVCDr0t2g8jHMWWrm
MvnI6uAVHwQ1va/Ve8F6X639gEuuOwXd+V9NY0Bw+SuBEXmu9yQW3wC8EqYKCONipM5IxtgLWo3D
ue6pShzBL3SublHnr86fIhHOr96Z4lAxUPP82TBdC8z5pBbyyEcINtMm5I5TXvcrKOD1JJ2tkMfb
DIOxNflygBlZMf4u9KASWrouckn+1OznbIUZ8FbYP00lM/wH6TIA8ZQYHIM9eQQO/k2mXCMxNA4E
qmgdmlwfsZubMujAwHx5FaFuRIQMzsBK2mghhrVYzzMqNwujPjD5ph+zdfsUOLeNdetD9W/St66O
XAH2Trx2WrI09qnlPNw4BObTeqeAGgG0yQbcaNRilE4IWxqpIlNLPDBm7YH9mdqv9mc0wKPGWUs/
aoSPePd3uny0oA39BV/6LZje/PmEAkgp7vy5L35eQ/4gNdUMpOMiIMfkkioBTr60Xmew5eu2QC8x
gC7+CmkundPfCnojsincYIv6zkDoUkc28kNI4DEqAFrorMYNedqQ/86WVdMnqlSPXOaUYntjZPiZ
9W7yFCBMB8/nG8bqxzCVAzFXXQ5/kH8ijofeWfm+OOWzKF95HT+CzuFcxf5X4C8JI3kLddECkHGR
3P7cKm4rqsLLMwCXnWuHp7j7+0EyHMD/stTchErQ4nfQ1kiBCoa6lQ2LUMpQo4gKWcdWqSerT5CY
2R01zTxU+P7svrFboaM1NU59Om7zWtCaAFsKC8Z+XuCq/LIGwPmDuKaebx5rb4+2WjtFzHbYsiO9
M/iNib/+LwlGXh2VaLfC+jCCm4U8RrjWj/U03dLkDExQe2Da8Fn2kUPKGZVB+TnPK0H9AX0FyN6P
htJ4AjHotV2xvJ96n7S5ecsDTgbn1FgNpt+j1KVzAxKRmsad2pepsnmzbBroqw2a5nmg9Cazl5Os
lVJa54wHadcVyHUBV5ZaTpqTSp1UkNtIexGDDWuQTyknmG7bSQe7cFk1Y4ESlT5Kzc2nYVzYQc/A
xQN4KEYB+uhoJfE+igKHLt6UhA1fumw6b/S7Wz/uf3b2/cJkqRnHynvqxvowVPj0XzVBGTDtmd8s
nwpz8uvYm7oSu9Z/qbVljtN2jNCpPuGmk8uVTPxJCkRx1mhFp9LCqNCXJUawfvBhh7BleDPI6Gql
M5nY+jYpI7phRhJoA7SwcJjEK40na0BWqx8e3t2F1iNF4MV9wwVF/VQ0H57pngHwGp0QEbcrdwF7
JFYIBBmQ2uNLEWmLMkn6FYfxxi8DN+aBiUJWGsmgiUDNkN1xRFSrazCLrYDuWfBuJrjZAjTVAQNU
oR8mRkc/rZhVOzvLnPriPoo+Pp8wzXpUAAGWoWwQmvc9/QTtVZERHUHUlFY/k1wh7HIgH18UyUbM
E4IotLJmX3lMyHnRL7QlKJbdb7ZoJNbNe7lP8/E3EjDRIiZ0R1E4gf4Mm9XtIFvYwY4usCQmefOU
trz0AFVHk2WnsaIVGVWkMJB5M6NdZyssCb0UgmB7AOEhl2ZJ09LX9LFnSXsyrU/23UWWoKwoSQ2l
wGjjUhSFrldPxG0ypD9eHKzqZspoTLk+Al0YF5srUChrd5c+w+F1AF/fbdI339FS4EJ/pTLwTGdt
/E6FcBos5t+BfE7G80BRbTkQESBegaqk1S3GWUMz3yWF3cRS+s3iWug/3HXBHfirl5zePHro2whJ
Xxcv4UzqVdUlPMxfSRr1p0AQiKLnA+ODSHs1PxZGjRpEadMLlWjKloikad5tm/hbHXnWrLqRdtaX
3EvEuJdPQ7/LzPA96eK0Rskjth52eUSbgWe11AvvyrU/2CyZcQPufTk2r+eFWj9UDwJxtkUL52TN
wzElf0mUwuvRM9egTydfnO0/o7bCtXIqwMsmVh6wbRAeJYGCWBXY7ucfctKWN0zNRmzQtbEDABHd
Lma5pKokxgkY9Kc2XjzwtPQGBayQk57k1mMBTWTZPSerTSMvPL1pEW+wP5RKDiO9UGbITg5P4cqj
rN3UsaGO3g0EQTyW5IOQOaUpm5bkUoL4gsEjAlgVzIMJ+qJtlppfllhnnwDej77JldekFKmy6iBv
kA9v1uN1o33l2S+cvr3BJjoeMN6HkH7TpoEH6S3rk3y+5grzXrifY+mKGXWWggnSd1UMBed7em5V
Dey+NgTYMMQjfGVaoUNNBTir33l+ilWO84/K+IT8hUmwX8/3/YolfzAXtEYKtFxVr79Ej3hRDHtm
DFCdIV7crgCBHmPt46gJ99j227NuYhtEYlKpOqOU9R4vJP1+1pT32uTho/rH2Z18pECGHdNAUz5k
avUIMhFOvYvU0cNqL/K6PqClWmvN29lEbRXnVrSxyXbdKEF5twW3V1FBEER6IznwFJBh1avXQLCj
mwi3QdrCLddmV1BLU1vskzii/HcIOvwBe+ViIiEwEkys6/HS7Adgjgn3f9DqnrHJolQ4LbYvyFnj
ESKTBQli57Pz2hv54HYJD+5QzCIr7bEIPROw1bSRn0rWh40AAo6BzSU35ajBOjkm48gvZ0TFxc2Z
Bak1BTVifn1o2bHmLQwnX/+8AQRFfq/mo8KKLVRzjwDVDIrS+agqHbuAayJ6nhmRgi/krGLOcYtz
56UItVUx+e334H4vuCHOEYU2zba018kBRzbGwH36a1bA1qsZccK3w/fe4xA8G+Bmk/tJA4vESm94
QpyxuU1Fwk3BvixdtOmoU9B1CIPxF1a8c/tQXii13Ov859krNj6APZg+DAvn+227NYc40UlxTsb2
2GK0S+IfIIcPgKU7iANSiT/h6vQihC/QWFvH7a17srS6TO2HZPXSCRoPuAA9y8hOA4ENa8fYJN/+
tbiGNaXrmfQv2RzcmpK1/Ueh0Oqf4wkosT/6cOisRIt0O5HfTK/4r0PT+RfElYV1QPwDKmGrKi8p
lTuo/Jud+CIDiXHneg+th9MNxrqV3xVgy10BBjVVg8tJhnbaICDfyzAzv75Ief+GNHayel5JdJRp
q9GIMjsjWEyCoevv9pjKLHHF1gTT9vnc8B4RenR2tU5L42kYyjCdpre9F2kYMiYwtV1fj9FktuJ+
4w+DEBYQ7bbZgH7KJatLslmD9bMzVpG86nafBW33N4iCogfLSYTPid10k0N5YRNnOkymlrfyopGp
cru0j35cUWiAO3dYm/wGvWy80n9UR5/eAhB1O2W2zgd9LysmFtZkMtACQfoM7UyoyDJLJaKW/Upn
MaNXeJVwB/hj/A1jc6hm4vefF9lZbBVQ888IIKxSAuYYyaO30rViShsTXN3yUJ9vje8wJsajBCu/
4MRbc6+YeeUB7MbaynASVi3LkNQ9CyOY3R0NmvxaK1VZDZcbHvNImXYaEsYevdGiCDBR3XnsrZlN
FlW5+HpwYxmb2J7DvjV/GW6Sxlb2i2R1KL2A4wU/1am2XvN7ssIqbRFm292ieuMFuAxQEjc1Kfe6
xdijMIkOHdgitNc5e2wHVbhxa5p+mPY0g51DhisUfzoYCmjLUeQUVwkxq3Uehe8YT6S54oX6bNMV
2wyx7X0q1LFrI1tcA66g8Hgh1pLOZjnaQhcKcyyJgPCHEPZpdm0Hft0R2Dj/CZpF7mZIMYDnBIzx
3PMMGNg6nEt+FYlnFJRl5ZgSnqb/ITuMdvqGJxZCp0jwagZ4ZnWVQ/ZBLQjLf7mOvNN/eUN5EErp
QNCB7Mxq+IDVZzhaokW0OXC5u2Xz4qQR+uSD8p7q32YkCqnThAZhSRHhsDGE7YZIDWD/x3WGIOSl
zdmd+Qzr7UzBToIxe3v+ynnvvmcf2RzHDDE8mL/uCipdPtfYGygNGKtWKBJZhITiv6ayyp3eClIS
5RPztCYIVN8/1Zg9dTLroVBJco+v9Og5vfeBhrtYqVP447esVa5pSaRi4pyRKwb3oWlXyHWDisk2
Nw4js1Zz23ofIcYe5Vv09qj4cBzjcv+IzFQZJD2kwTwR9pIxHUdEcFRK9IQQFdXoT4zrMXd3mqcA
V4vcvwnAgxjFJOkfBX24fc8wOV6vu+olWhuWwZe1sR5uBeOpf8crtLiNfUUbdPFf7p5AzNmNms7o
y8VHhYiNIrida+2ZaCgSBRSdixbq5wFDIBjRTCY9XTLxKUs/BBphLNeHKhbbZfcjUvbBzT6WoZUm
qjoZVW919+t8E6p8moYNuIHgebmnkBWbHF2ERGtcejHSrTS8lcjKWjDdc+5dNAaeu8XnHvBK6FuY
RtrfwXPqvN0wT1KiIS5BmL+8yYRCwgtoB9RbiGpWp2tYlVuZlfnE4QWoBBj/tXfikRsLIJH5wAbt
ZJngM2l5jIS453OsYjDoCrk90MdpW9EFY06vzyUpdr/pSQoDFVGGBrkjWmgSFuKdY+6TAAh4wXnG
A8Hss7cBjt7geyqu3fn2VMSH36M4zWMbSLxevIC//wttr15e5hIE0qikps2Yo02IJ7TrLIA6u47m
3SF2ACSt6kyMi5hfOizZN85uvCcCoqaUw1TLS2npfv9AlnHprpXHhBwZW/eA5+cYcCua9GfxFvCI
ESkFa5D8jsbjPzT0dWEf3uvWKBfd4DHslTk5Y4AKWNYUwiRKb0FShsqjGYVCLyGLQSEXgZuA2xlJ
vl9vVkjVLIIybLz71V+TwRmQSla911jIcyUZLVnQQgQc6KvoQP3ytcdQRkRU77uKCwUO4YNjAxJ3
MIjV1xJK2Pr+0TsmfXNkn9lB2BoiAZxolGe/kJ8tRMVtb6ADAyX7XbWTbd0D+J3Aop7Uh/H8YUc3
XI2Yz0om0zW7LovsgN8OM7pI+1QCqNq7z6Ccp0zwxwjRc9RkK4yEL7+PtwUPHvD0pdLGJK/umSpS
e7hPymCKAK9i7/07398j+77GWS2dz7Si0hrF9xJSOmQ5QzmCWqoV+ifH2aIaGUj+vo90g/3Zrxuq
Fzy+Ovx2DaDC9xRg+gZ49jrPditAyTOEN8ODXB/0kBOF9f2c7WfQSvjkzv0ZIXgFNrBzQa4ZfawJ
KfgpNgBlLnkFXSrf74kbhpVIZxGGjMdzNWGVvKf4EXng7UcNz032eBSTPRyMMqgyOfY5vUA9Jn3g
N90MkfTJE2DN7u7y+44RhC5ar8zq7FHEyO9kV96WLYJWf6I8Rd40QCXlQJg4sgQLshBFckBbeT/m
Jx5m/Xh8nQWMjSzDuNJMUhmh6CF7l/zXIx1CXtFGLgwrH3E8dbsILN0G1c0ms27LX5JCU0GIaQJD
vsnHshZHDpm1wtT8saCBnt6OHZc2ho31CmVJKDejFtjNn+26vuLsnVkWRYWTgBFOkWWxeFTEXkuu
uIiYo9GL2mI99pwBUNMnQTEMteFakLqxXnvXSpeHC34uNhpM4nWJm6e78wHc7+iieXwrPq0pLcVC
fHhwS/fuuFkb1Sr2a0Q1KkTz2T0+u3UecdHvb/M6CRVHXNNS89rZ3UH0tErI2CNxptDccFDncx7P
Iay+neIuNk6CdNSwBrGeQ6+o6jHkc/bfky9iMPE/famkENEkNaHMO7tcQSY4JTEw5SdmRfre/8Ss
mOxGuyJ7iwxx1cLphmWWwtr8qxcAA4OonqWpxd9N9XjNwX2W0RnYk6o+Xzz+rV3jVELQgJyplNNM
cxu4IyRvEvHqH0Zcy8dozp3dCVmydHFOgtcpO/cLX0vvY9Wi/XEjmTKQ+bxpaNheyub/hJkqCA8L
m1Dd/1EiFAsRKMfpTObhHkvWf6cHcwmnEWQQAe43Uz2EchO63uB2yZ4yFr2Z/7QAgH6CH4Tll29q
eq00aJlcU1i4oSI6fCI20OZCJ4r+GtFPLFjRsGBdrZJt5wbBpOmS4k3w93UuboiSimke3i4YkHzQ
LUzG7LkgR/HdJv2JB/RAgDJdYlzuI91hzi/g3+xyG+K6MguW3iM0t5HgTV1pqpG3Dl3NsdGtvYFU
8rf54liw/ri4+FsuhSQJdIq1Ei515nV5mLtxsR3OW3aiy9k4J2r9X/cTTtmlLgZ0GRn92E6ntOga
l1v8Vbp7c2MJ5+NZoRcu5iQVf0Jm6L5jdjSyAVFh9uxFgiAY40h/QMzIm37Dj3MiXZMjkxCZ6JDQ
Nv0NuuJwYs873xMNyjEF4kIGyXQ5RH+6q9IJqZ88XUKTB5t/Wbu3Cm5WNGwmodYUFOt3eIkxWm63
MWiTtIhHMlQGuxuoCO0n7n0cnqpjdx7EyaMG9AJjAZcggkiqgc1fbyfPB/BhxhmfsWTkDnLnfNWW
JnxebRvKTS5uldNe9ibTPqgWwgu6/yO7ZBrb2nnyo1GxU5b5VuUgxme620MOEvqD7ChA3iGAEMO4
NZWI+KHp3JVK1lPkLqYZBCidsChxAQo5LvsvuhAaripM6TpK6ZMdQDUOf03Z2l3POm8P4M/3jSDe
Y7/aPGSIKkl/R3p838iy56HisdS1Q51ncF6AZZdtQdmymajGCHiGdeNx5Hbh7jMZdJQHvB9Yy6ph
64hnMSq7apfM991Jl7I13LhkHswjm6WCRAWO4jX8ygSveSWy7LMiBGoyw8X5JFwWIJbYvLapOMdR
VtdQRTuTN0hUwPICtEdj7keJ3WjRidb7eyRNP0YDRyrSTz9mljaFhTqF43wOsL7PrasWY5QAv1Oa
bqm/O2ZzwZdiHn198PLpKLLVNtJfioGAqr4ZHjRxBcrnQqhJDFondDljJxbgMviXNr+QKKONOH57
J534pqJjvtvUPAXiu731gG1OjEBr6FCubz+H96vIXpdoz6vSnookifDWaT7RcUDgRVokC9n3z3KU
LzTTBCOvYcXkdZJdwaH8SQGKurLVowh2e6SzXF+k+8fRzg22Aoi3OYEfGVJL2rE+3SjpSOeu4bCL
HAImQzjt907eNv0yl6kxUG69CligYS3ZY60L2XuRQcqA991uQXLo2dSjeJqatuv/UgHcz2EGZtMm
v0QQGZKLrGzLk8olyJjg1Nb9HbnlHtgpGVsIqOSGxGwLdBRICIOF2h62y2gVOiihb7XnHjjIy+d4
SED618nHPt5gW3xpxuIE7lMz/M9W8CKoHQlVtDw8oLzm7xDAvnrOk+yk92tmBnc+QecPPzvLH/TY
odpYQaN7qxPxePszpdUdUvYBPSiOudq6ABAO9n6m/83lf9d0uoYzHS+SeX9Oz5AWFK0zDxCRXxqr
uUlnsG0292k7RQUf+HKjN8a8KVHONWqYg8HljdU/JoF8yXbgMjjxBJ3tWn8R757GZQUENCXFsqYV
XWn2n94rpj0Y6xq5InTLHUrai/W/f/5jcZPZY0c1ZWGE8LZcjAtO8kkZVd4ZdodJjgei2//ovEqa
Uupd6FcJDg6cSxS3h5g7Fa2fnIDBqmN+dcNFS9NuMAkDChOazOJe08fKkpl2Hd3/8XKzDsc3uo1/
arGWm+Bvw95KgQry4X5TEkkGbvE1myK9VtKa34p9uAiE+yVBZ55EL8cTmP1HcxSdTdoubSlPhuEg
zhv4IuejNsu17q+OQ4VCkHtK6o4ASKS7CW5odn+yKXUOfV1c8ghvH499NI1E3lcdV8r+ysIcYiy4
srj4m1GmK//ip46c/CokGUj3aDaYppVt50yrQPiXpBjSYH9GrEO6ZgTyJhYgWHXMDp6S0KTEiZKv
YPnktmRzwRXTvekzeDc082r2tLWWJ8FR9hD1AjwjBWJ5YRPwMxFAddHqJjvAm/CpdtgsYo6Rl58a
DNpSErU+LAu3xeOq8d8bS1rIrQGRqH+o4CuOVpRJoorX71AeEmkMS91QDu0mRU+osvF775fZogI4
O6dh2jgy9y8/gPerdXp8uwfdBrqlzYJmk/NysRDdy0FLiuc1+HY3OFvHayIexLIFxOOypIfJFpxU
BGTnQbkJUz5mY+nNq0vFR532KYZ83iM2pOAYIuIUyR4ZUnwVheIGn0957C14pmwFQkEngOwG6yp5
mRjMP4TsMuHNQyCKvMzrJ8YFGIs6ff5Y2m0+lwXpKoz1pEqc4Zfk3OlG3RW7RjPLfpM+tP2DckYR
+GaDykLC9a5O8Q8qmWBaU1NXdtnYaAD5VYwrkyEobup2Cb/Y6/2PX/QT1ZQLJsS9uzSmHMF+ntLP
J50wszAVuTDBGLJ2hjcF/JSDcFe+SlKxn2xkjVuQOWHx3qYtDACaFSjvm/MGl7dOBPBeiw9nBKOS
7cl8IQDCkOwEh/qF3U5Q9NAMDNxy2EHe7iIkOaSJbK5wPJK3ZVnHBv0RUMETQ3d+i6hBp8Ngcdfa
Hvo3oUhmAXiVhBdlhjopt+zDq6TAkx8g1CWFGaPyyMwNp8/JgZXqqoeuwGbQWuDvqDLvaecUHj2T
SWBFDG/fkUgIK8nzr0L0q+ojmRscAnvMhi48lwsOdqWywCfH6A6EQ0UgKxjdj4baF6ZrXUsyiyiQ
mz+DX2GcngnLB2Q3V4/6gcl09RNKlNQvxiFCLymZng6F+btM9ap6grXY1NYg7DGpj1bhBGsPxMNE
3iDgO/FqFo1Z54Zi5HYDY0VNB5YUNK731B9vSQc8SZPytuMZ3iRR02jsE6tdClmfmgvN6JgRLAhs
YaRQj0N3pDnR25sGPGa9vhTz+IAsoOk5BFIV/Is3HnV1fP/wIq9EMM7bQckeb4DSpkX6J/4iVlVl
YOaTEwmAXGsM2qMmHjOPA5fsoEJ3g2a9yNy1prvQlw0uTC4pjbosVEsaVNDLGicgzhpa84IVNFJ8
Rn+OYgdGMk7tj89Cv/+DQVyYAO/ZrQYNn66WyDC8jQTFFoAUM+dh3GaQxwJYll+91uPwPSDuYsq7
b/tZSuLRYXhAPDlwJs/WPTHOofx3OzPloRc+4eUv1YiRfP6caP16dTma7DFZuDD8Ztg5hbqvqwFu
VyNP05XmaEUWN4p0mdjSbH9o7ZZiy3RkQFZBLKcILo3g5i11sao56/EGLi2naJaFO9wcr0YPvNtU
7tXwJDQNdb7l6ddEyvr1NtfyNE7ZOeFTWN7E/zE2qE++rn98IXMpuSCLyMRHE/H1khdY0Thyga9W
VdN7yQzUwMVmTuJHj7IIjw1s5GZdUOk6Pr6hN7Ljj7zizWbP7e0uQxd1995bQ4xxy7fp21fKsNqY
S40DDSiDzfAxPvA0GD2ASfQ7PrkccsvFkFEsoS3pR53ciOz3T2d+FUEqxVblfJBTxYErdrGL7cg0
tw96ftjiM6q7zOv/LCzEdx6V5yzKz6ij5xPkqwx7PIe8LnBNaB977IFVNl1A7S23VEU63nQB0Zci
nxy82LL5uptybo9b2YbaOuR/M71o3jDivBPt9QrpOLUs/3d5LxZDiC1CdbYOXPHJXDlW/+T0cgBC
MEHFHI9hLC1nHez5ZUYVdLK4eW5m/JrMBQqyR1+jPQnQzNEogrkG9vH934D5ZdlJ37hF5wjZ/F0Y
8q63forMs7Ue0AyF8QnodStPIuq4nn5frTtwENKGdZShLifx1pdy6jbcHboGqXzJxM0dCyjlvvFx
LLK0M1pAV/m57+H52q+mC55GNmC3tzmyguQjR+0DDeCeBIEIJ7jLF0CFnGQEYDYeg+rMDLcdYKYV
URbuPy+by4xwZFoO7PqABuA09ybRxENUOglptyjnqO3x62HGumalw2RTEyjLMtAPDM7Tdho4FJL8
UR8eS58tAb+O4WKHMPw3/1+FYVMie2Iwo4yt4Hx/MtIqIHpMvGTssFKi28P+zAV0j2W7xbitDfS/
xpTSRmRCEEVQnZ0OIq/+Xq8lobflyr5qbH+WZFFg1mrz4XsyTjysg8Lz06smw9Bo5kMaPiLHmsXQ
NHGJaaI9/iAgGvWIghA8a3CtFtUwd1RCu9lA7czUtqpOHSdwfvT/Pob+LpO3hCkzWDZvYvUF9lYM
3tQs96CJK2JnqtG/ENUt4dZejR6nZq7fNlCfWWXRPDMVAIRcNh2qlU9Nxx7qQK4KFZ+HrmFW6JIM
mOU9QaekVvyN90khOscX6+8XMGIcE5KuULG5oxnOlV4thh0VnChKlLAYksvgdhVOg5ut6FsQydlt
C328MmW81k9+Ug+8imxiPG9zW9GUfGrSoAjdIBVUFUV4wrp3riYwBU5sS9LmNmeHmif4iCXX9fZR
S5q4wa6z9BWFVD/zHCDYZ5JWll+nVfcwA/peZ70ltDoiRx3dkFnvroRA/+M5DKIRYysfmZv4REtI
V1K3cjmSSCpbe3DW+KjHAlIH6/9s609e55rOoKSvusmtDFq5VTFpenF5LpOt2IGQ5EZnZbba64g0
lLrOFrmETQYgb5gnIevrFofEqlsISQJt4BtwLa9VKtel2IUTQODBj5IB2IVYqeF0pomGm6Eg47lD
MUsiafE9IwjKuXNfd5JM07fZM7c2g0qiqgLzsmEiZ2uLHhHWwb6ueJZosbrn1GkkqPwkIFwllBsB
FB7jVfByJ1ICIqKXQYDSXm6oBfllEJ6bD2dgy382b4bWAEkoCxxX1HPdey0CDhjy+QpRTtzCSlVw
6N3zwKJnv+q5Bd2ZK1KiSzzToHT/4YXYmSBkFmRPjK/3KfF4yQ3wCaIXjv2VyuX4udhk+gOXoFLJ
BoBX85v0s3K8e6/G3lS0Q+A6oyiYo5ACRKkb/1MclMp4kQYU503tfxZFtpK4H6TKtU/2aHvzrRPW
TTCmfOiYQtYCpo190cseTsc5o/jczfugLvK4dLr3Q9qkYXACieqpqvSisYvx5wmIwS82krSX+jmt
pTi37OrupRu2ioiSZkhGSNa7ACMsA5RpV4xXaRXZKrt5HkQ2j0RessxrazhyOL01r1vMMU3AdO9a
NgwvUxBV6KLgJlxF3IxgKELdCNipO4hzked+ErOKVPtRKCv2aKJ/jsqnoZl+Ncdc9E++NO7Rls6T
uzbL4PAEnRcLaRRDRUrU8637mBbNETbq7zX97mmpcgx3iz6mIQVwznixS6jKlcNUBB3iqGIwlP07
mYZoZsQHUqHvRrwT6XCao9H/OPnxlccDqhKPYRuj8/jND5PajMymMZt4LSILGQK6JMkmlTyGELuC
WPabp0XtO1VqdQ2B7NtDeBzJqKHuZ42lUANnMXCBTRoCYSiA20WN3taJd/4Unl3q4AG7uduhlstI
0cZq4jpwbwWCZUxbecsmCKr5Cj6uxHHfIuLSRUf4ysrJsJ7hW9DEdJhf7hw+aSjfo9ZNg0DpDEf9
talSeWjAFJIbYSxCw24px6PmCMC70n1vFkUayhZpKZc3jG3V9jvzC9eRlq6nTB9FRHKFDqtTZ4A9
IrQRfIpxQrGbenvF586KUGtkK95CofeSpzRbPznO5FIMwyQOt24JCktRs6DsxTkKmx/+fVD3oIAh
i49UP0y6Vqg5VaFqgg9hrKskPiaB1TC0NsJcZTV5ht3BMCZ6zEET50ghctHgoVp2wSgCwbtxpKI2
mEPN9oH57oxosG5vAGasXPDAWDQBGcM2QhQNSBlFIko9733c7TFcLat+lF8MyknCIt1OS06NJ256
CyjtOiQQB/BAsdj5auWNqJdsezDcxPGJDrLifI/VJCginCZrbQvhh6/zGI7bTaiwYNRYzPS2r4dY
4LfpjVI4x0V0Zgh2wL1u747Z+Km3m9i7A8nheV1aOwwC2Ib0QlapowzSwRKQrIw/swo5vPNPBazI
RhcQ5dvGzQJaxAhpDNXVem5b9ZEbXy+TfZ3totK4nE/fIizEhrWerkO0D/H2UbBseBHZsB3bC5vf
l+7dLtoW+9BZ5BQnVsxchnrpeomzkE3eJO88f+SrH52K6AiKProsYxkR/7Jz534YCxUZyWYjJA2k
lHcBVHAs+Q2otGc5x9sa+gQ74ojfmT/Jtg9c3lTkFwnJCU99WiPiZCnYOYJhyIrJc8EtkbCH3vjv
c6YZKuKvi14N3w1Hpb0/az1OR57omVdou0Vm9epMM5dBhRakeM1mAh3IqzAUK/xUyRjrcqxwjxFK
k7GVbLjoUGgfRFS8Bq6FKqvux+uWYtm0Rm3A55D2Vd8pRYUs7FyQLTVv56XLrtYeBuRwBGymvsMQ
biRq48MjFbaw91khi0NC5Ee4RwpVTzfvEWwctrxt8u0BhalkqSNzILyMPjj2r0/6WWGiqMYgwXGG
Ir1p6TCyyUqyIPvibUaV10HEmIkroS5EsSURmfnan5zQTsdkOu8N9sDKwrJsxikxA5vG7suen/ht
PVIBhMIoTp1Dh2+KmeDeMo0advHL63k8hDMihZ7OWgqYn05fYewFYqRUBGOWDDtz9ojtG10j15iC
o4IWDEnzw5NeSi71rHiIMVCsoWcp2y35zt1e/c2imuW98j3vh9kj7chugI8wm+vBvUTo/4fwCYFu
HXikRAaLEJWnjuMWy9uStGONHM7MxbH825KnjsOdco0lH5tHSurLQq22SghqDABOPoH2OG1ygmiY
5/4wQJiiBaniedwURyuDmyl6ongIguIqJydJ6Y3tz9GqiIRclBAliiL9Q06cIZAbD8NlmFFOw001
ysGQooHwAkO8NRBN9XoYwI/NavJdCr59q5NULjLkeaMyI+ppq6Id5m4TaE/i3XWHU7hkxb3Ft/vx
uBMliyx0LyvqSdXjLLijiaT/4cLCQ0rObVgxI/v2it3dqSDcmSE4EyzbxORhITPrDwUnFiDulcmz
H0qVzVxtR9WkndXuFoPIgrEosJ9LzbjyQ0zP9Vb5Ad2Dvx6s8MzegfuLOpyvhMFYqX53dWlvPor1
1XqFiIDcFAx7FrZCLLhq5yXT6C4ZChep0oFCqH3Jjci9vlQ0W/jpSi1AuF2rfkmQ3DIKTdU2FtKz
xgUDZkEBeZx2DVgjYtrXKYNcKTtVGKpXRswqER4GhqML3sFmf1TdMNRpK6XBDuoxSKiyGNd5MPRj
iVyLnPj/3IAAw6WH3SDWaNnNPmwWPxhsEOBVvtA9TOGr08yX6mxZmACuEcntlwkWGrr8YYhZD/tQ
+FVqLy4ldc6ra5Cne4rBdnh/Nq1erDREscqsB+f74Xj7fo+HFbU2BEUyrIyIFwTh1MptoK/9/qVX
eW3tCuKG9f7XE0HHnMCo5va+qHbKHpZyvMpRGdK5F33qaNdUMAi0aUwO1mVWZ/z76YqXCd81VoX7
j0mNUQYFfsJkW4s23AuVdAFdOJOQFIqUbNZSD/A3NRN9nMpF4k4KrN1YJX3v6bt50j+lBmXP/NMb
hi4aTQWPtyjK60187Juiyth8Qhd9FmkKoh10/hqzxaZ42iT2ZN2it+o+x9z9EA7OERUAkU5nUzt5
nSzOoXetaO+R4y2beYhZSGZlOQ3Neaaad747M67UwF0pMNVR6YgEUv5TgNYWmb3PgHTEvdk/he17
XG4PWpeUe606kt8WTn4KtW+oi7HuYfm61ZCBXEMYACmKDYKQMLoonbIfVAvQBFruLTEavOunW5jm
SEbGWbCCgu816n7zCaIEy5QsuFHQK6/llCM3gjWEVgOKU3OE96rSerpUZY5vjxYByKTaNiY8llwG
83fvehyRkCpAfNJKvXJzEQfSbHVmdUNpKWqROggqQ+me6Lnhz06XVvBX+3UJvv4hKfOAOyYhBpoy
kgtrmE/yWv8JvJXA6PfX1S2z4wQIZwRmhF7sV56oGCrRbRJll0BjG2GMTU6ivtsELVVuSeCQFZDD
zlUK7lBTcAzDMkPN6vaOZt4Wh96ywEhvrXtYuVf3ZkyHWDOZ3KHxc7/TnsjST4m7R289vb4BJ/0b
fuM3mFY1bmRAFWI2SoiSJjfSpkXv7B/o7b5SdUT5wggmYGiWBXX4OMyBpTnw+AvCA/Kdtii5rBb9
NLvR3E8hpuRHhv7gumeZMgkoK+fjdZXkHJcUUykVTwehOzPU7PL3+7SKI12lX/1/sJpV6mt8vtD+
dGLnohgi6fPw1v0EVb6p3KaPRhLtxFBwPZniMefYGhgKxsLQTs7XaXRqo4QsH4I3nCUKee4bTYBz
QjXxbBZ6Y1yWzCYTtMIU0ewHtB1QXMGNvXJ+J/4DCU368rWiYlpJd+Ntqeaxmka5lRTTp10Mh1F8
ywML/drPHCEWJQRN/IyJ1TVtA1Gb9epANAUPKJAihE6GzRIq5E1Hra2pv25pvCNaSdPxHb2vLYhM
Xvbvbtimlqs0CHI0VMt2NMwBMUqetFxt9fLLrJQGF2ylx7lo9w/gvl3nBdVHfc4aXlzfXeOLtvJt
dC4CIqANc7H+bynyXCjFsZhOQ7NeOnhnUS+vBKtrd42pe1DWnYL4kSz/39wgRM82PlEk96+zk5L+
i0muRPij7FHevrXqta9sLbmt4HUa/Bbe8UQtXlL3fln0Uv8pyMnKYdAYAoP/ZZMQZ15BzWq2KiGZ
RYKIAq8NJoYhByGyJJyV+7SKLSBYnSOsHKxoXnbNJXoIKx1kmR3cUOMTobXJKxPOzyr6KqW2ZFlZ
WEama6jkehENvrrlvT4x4TMNhzchpCiKveArrcbO4Y4RMpV30JcppruQD2WYzYqlHhXvIv62tcMo
VLQ+iCm15xhkvQ6+BUyADHxUasxYx+WGQd3XFD/ROtorXOSWbMqvOemh6/d0VrIjXdsk24SnSbV4
XBMkTMxpOgqawL19veSt9daNHPZcQ6a9T/xsZfZW+1XlKCkbVrvWzsKN+XE/V1F1WNfZ5JVAlspU
vzz3MhIG2MtfmJcLe3qFnIHoXn7SIWVsjTiO/+UEYmzPCcejxZ1dVcCZ8fDFZ4o7xGfJfPME3Q9C
kpHcR3ul6L914ZHFxKVN/Bp64K4z7rf7+XomDGm7KNsZNMCAcfZ6z/FaJnHPdlzfekp9/zJ59tm3
lwm8ZYGT/T3kZLRwdQDj025wEBISgnDkKGCVr4v299JyHrLr86p1cC244KM7eUtGiX7pDfVcbcsI
N9K6dW+cczvhK6N5ZTbl+yVw3Jjf5E0f0jHSEQuJ+z8rBY2QPC+aFPQ17qbQOQyOGyREwYJvu2M8
qjHX16PzXbCfXm7hBQt4DiLvHa7YTHjImWpkVVt/NxgdAg07ivzkm8DjGK+8tZ9B1L/9GNpoaJr1
2X2sm/1nZ/NxB9wxkwBWEwlE+l3X7HCXtMZcoFgh9xMBrmRMzYfNfvh+wSf+SLnA3ZcOiacQ3ekY
26zzWbRDEwng7CwK2kA0y6VP7SXo4V3GNn79nIyoO4cmmv9bw4VYbW3fAF9ZFRGCtwKaaNGazBhL
5RbuaNnwM8YlkZAUoSKW12JOEooxcWFIUZiK5srRbLITZ4Fr9+0l9yP90PddPlU6glfLM8bNlmyC
JvVJVSLjLbb6knj4Xj2g6q/mJtjyb1Bz56zevm8RawvIumDqUk4QaFzWm7qpOP3Z0YQT4XhaPFrM
NR5yaKjg4+iClC1LGgnGkAPnUAapXyz78I+4Kekv4cOlMGn6SqazVJud8fg9x0HKbgcWctvOd6UM
LBLNZVk1nXkC2JOW0QhwP0jranmZy5oyEQabzs4uejmIEDeui/FNS88+etxqefpqJ3KQb9OpV3W7
lmTXOCYPxhU6aWFgOZ3QYMn5+X4xEgIzTl6ZlvPNTOZA4KMY1ptD+WFGuqvmvgwFR435QthWzkt9
jL3WdhqoSoN4HbJmTZh35rv57a8QBOBSaLCVLUPQ6ALeqqPsI98R/kBRiny8O7fB72vRDFrFnnq4
JesJAGYkwy4d+3opVVF8by4jSNIngjpwcKH3NrU7ErKv/UX7lsTe5I645aVwPliTWoNcEGpc8kMK
wEP9wi0U0qmrNeM/Tu+DFF4FR0Y+ZYgsJIhU3S52DIIjP3ABfMQgXL11jQJZH1hQ1jv2/PdLlsm5
+BreTDb4FtFboUVZ2u1M0P5LhQLglzGKZ+AmqdbJCcYTvAyLDW9RvNYW1Ta8j6ARvu1XOQLz3pT4
6S0GPK5+osDjvX20apKTEDp00a0tCtuw+BVx17LgNunSLZucoWmqxx74i2rFq7YMHeyOaRV+ICkZ
PIr5Z3YsqKhugAE0gn0bOftd0qmScIgWvof1/nfPhb1H6tXZBnensH8pH20MkdiBvj8COf9oWm1M
6Hy/55IS+HdXX2aDmn7oyzH+TUGYnzoFNmvmV8LE3M+jH0kyAby20ydvrqLxfubVoWBsLeDA4rtu
DHlcTGzx9I1aKU9sUCXi4EAYcO0yQM7nIcwv3Hgxy6UYT2J0hWuu5Foa9qdW71k2wHhr+Rv/PB7A
670iin4ajPYfAtEoWCwloQHMou1AYkJUeu4NcmYzUzHvrY5g+KkmTaX6BIjBwLYybYAVuyNiyR07
P9rF+GJldUpOIetgt4M5J4bYUfs7ApNlm2vG5uwLPgqg7YckIGbbwpKFCISC9dyZ6EoJYk+pUOEh
KDPQ2zZ3O3oMsTQ4ajXAErlSOF1VWBOCyX9qNS0iiPFbMksP5oiLhMp0yLfK9EefAIM0A5OejFs2
nWigcYVwlri6PJQxvh/J22tdlpVUQRSJpEgRgZidXxAECWOlCOVQY8m0QYB2SmDiED0TyUzeYON6
/xnkKhxHQ2+PwDu/etljNsOCHWi++0DZ1vcC/D8kUoJktgpf2K347U0u3Nrz2azNLIt4NA3Oxqkx
3AoEo6HMH7lkvLlwwynz0WATiJanQSNqKe74gmKnrSXWIwYxKw99AhidKHpviX9wimj9DOqMzRMY
c4PzmonwbZtWuKUz6VeQnmsEzMFSNiccOt7yP3kH6Tqfyk7+QvnCn3no7qfiwz3JQfH5nnynt8fr
DH7Ie08RqSigbrUQQoBgQeSvLqktH/8eRnxAC0MuDbaUUqEK9cT+3WChD3wpWxTGnLfGAoAWAQrV
jeDTIEyCXdNG58I7Peaf0mG4jPNOSp0KmaZ2KszbHhB/9uz5+pOTuJnR+3p5tggx7yMRr3EeE863
Ke6GC8McHoQbRik5qEygRA/0z/0hEQ5fHWIMoeeocS7+c673uqV0fBxcEhXrwKXE3qmLyqXg4crM
nUyDPylcfyze2c5Y2MrrKvxD6dRvnLHRHyhX08Nvcq80V+mUbkkeOZ6pQ06XIO/A6QaFtCYIJa0H
KKxMY9r099RGpTZdpy7u9Iqe4ojrcZF34GsQ+AdkwmWkAaHjiPyTPnh5uylAXoZlGECpjEcJRU6a
uhz6vcayHCfNl9UOcaG4fE8Kb4LRvt5Oj/ErCORLrN1t78ACBJ2s26c5cNnH5B+xEoNfiqHonNMD
2j8EOqSgHYoqZrEkoTWNJLsbXimELuKM2JjBFNmLc0O3plRF4ckPaA9YlW0VA1vRWzu94emp4IKy
7hKuxhZekeZZKgIUjieuVVFMuYeva6wUi2uUNg16SS/AzqEPVWXNXy2/1u0+BRgJx/5oCV5BIEtL
bmE7mmZTuWqxV6/MR3B+21NKOCdjmEmDXJF/NDiQgrwkqIkOtUeRTq2IMQQvPxR8T9QX9ylJpdBc
NN3uOVeBK2eqJY02KTC+4EqsowuvD2zI4e0z94x7u9P4gmVGpTswRkv9A9SAX7DHiffftg5meSd7
9rDv34k1lr05ZZZTh//IiT5px1tucM2EJgwdlGrSsQYQfMGXHJXZnDjb9KzwdBw10lpMMf4sXryr
w+dBOVr4ZfK95RWGiNSyXxCDpII+5M3ZnhF7zXttwEfjl7iEVoMOqZI+QI2RSY2Y2jApXQPVqxZn
NXsWtIv892VWH3kHTi7ocVqz4pFIyw39dxKaX+BevtyW1jHdxmrVcyPp0zrN+BCffvanxxQk8lfZ
zGaioSHJ9wgtmjb8GP6aZKNhCOm2l8PNWgLJ5os+kI8fh6DfSRDEAcBflVPXPmhG1kjDdOph627z
nZRPC3TxQKtiE1lN1JMahwy4g6Tlnn+1x26rgj169ATFbyuqL8e9vVj3ccxiHr99DcBVWfLRAX1t
YrecRziayYtZnVBgOR5E2XBnvuYcQ1kplq81SbNXS8BO02qGPtHc7CPvOUG/z1j8d52U6pjjrtxE
+CvOXtt5zoHmqcSx8v/Xk/ZOf2SrirDx8zplcfctFm7Vd1QqfOVj4xOFgWgOwOicYzlEYb9cUBh9
aPSPR7r12yQO31kPZB66JZRIEKv9mgpAzNnHZ9k85T74hRcDYtvhDnkqm8a1/l3WUEIH9E2xU+sD
HZAE2F0x3jHwiLjuT93u9MA6AQkvd0APcGcCWjxSo+mz6Ij0MjGuPNgU5HPOm74/50HXWAcUV6sZ
YV8A3Kl7DkaaqwA3lJ4F1xx9jvYMUmAlt6IKyzhpMWi8kP4lBgcB0zcZfkHdbBOWtsEqLacYJBAz
TQTww7mE4zFgiqLpPmLKal5mmGDkcDA6QPWbimS3WL5caWZl6D2KY+bEyvYYfdWH8WPKEEKeTcMQ
2acylQhnmyNz4I2e8qgFgZcFPPNdpBnbCPxZVb4HLxU4LTXDW/1OwzZmvsEcuL5hYBFyjdRBkkIb
EVl88wrPUY7gncJQ7TB0MWr2fSdwpqSC0pclRLVR8cCrErAp3+adpyGjm2wbmlQaXVnZVH3R+BtN
GBdjDTQN6KxJ39lBZZtB5B4PUtsyBwyKWTapLewhSPb29CNdJdAQJQQysj3z1wh7+AcG3Dk95JfF
AVsAd4dt41dk3EM6YNB6RxZVPChKP93j+AfpDD45lLvEvX/sIxd3W/zPztnXIsA8tnv4hdxbChlu
E5yssCitprrb+EoFFKLoD+cPfZ7SS5VLEIkYZDm4vhbY1rzkhvsU68efrYdw9I4n72SKkzanyXUb
TVqOEY77WSh0OlLCzJiSoRJJdVZEZoLP9oU7/Wp9wlRg6Unxt/2Z8nwqgbotUYqdjJoBmA2C6S5N
9P4VFt/wVSHmfpxI/FZdqBQL5XFcJ0hiRxrqMTSF7Ct6qQ0lZ0MebWuZ0WkFPXHtVJDP6ccuhRKd
XMYv2HhYm7XhRzmT210Zzby3mot88ST9NgjCgiv4lWQ8Q1verem9r9tDrA3kNrv6xdKw9xIM21fN
wNbHProZ0CsDfAG2mVuKUx3cq4ZS6gbgfSsmMk51XHuSewchtExWTLHwQV+g9CmUU16Pq5B05SDi
Ojkxz9uj5V4o1/4KgdEKB52CFhBuSW+O5ESQrPcZyapmHLJ7gMfLwt60uBCRsGvwq66P8JfADbNW
+hjqcIYzoejpdOxz5Q2Dv+JWGLFJ8EnQM/z/BT3rgioK+8ePnlJ0VvMMYk3IduSaX8Fhgk8Gpn/m
9r+uNl2RBwVKvFpY0fIyNPgqXaMixnDR7EeXE9Yxe5AFvZganv5eo9cgsIcjXzSf4mmHB7vLNbsz
a8xpIEI4zX1G6AGaag4Gd7IHOmh45rMmYSKh7B9PGsnWBuxApZXSqjCsOOYu9ZKOcC8wcjdRb7io
+VAJDTBALkThgDIm1tPy3dxZmzjkVdmeN2C0Zs4Eq5+TPRufQ8ft+bwcor4DxX63JT9yyLw0SKTp
d8M2GOyBqvaiH1ODURpDcVEEQWgV7fvpJmrVvOtl9lFopzNoJf2hEBUSoCSCGYoMnVmYvVfIaeao
82AsPzy28uiky90t7m7zYSfsXu4sXPh/q45Yh8+HoM94XeRcGr3IuFMoOl9jI88EPZcgkrz1Fg85
C4WRlIXLZT2nlIlbLlQuuzYXZUSclNgTB+BCdUVhAQybNE5EgZNFD72Igw3gV5fpzN2rnascsvz+
KHNZIgdq10/OteIvDqrxOTsfPeCeWPY/4JLN8wNJ0rxRduaB0RngaOliiC6lpFkiL6bNnaLDfuIW
+Aj3/3HwHiP+gDfBTO1puOSv03zSvhLZgZm10ledjbm/g3Cw5Hm82DNsPreYZRiNzScYGoiRa0+E
2rdlkgLUOacePRXxMuYuuf2f2KE6IigcRl2nnRqZsDlzxBhF/hlCrWXGhPIzXHbtUEhcNqj8i+ld
CaBQYZbMkttKkn1pg1ybLOQhPbN8nTP5BYTrTnzAPUdoIfQDO6Q9qu0vgt2XUHsGhtk0nIzCufLc
zlAEg4B9xyIGEilqIJWJNOtD7pCsh1b43ZJFiYGcq+7EEjuE9gQ+Ru7233NM1Mje9IAMumzofqiN
warBWMoVHXMbqqbYMS0Gad6DRcbUWbAk3okaVxKUbclqi8Y3pqIEequlRPKDTAJeLTMVwn6B53ZT
rAczVgKldDsSb17J6rmRacuNjZRBPlYublfPdZNofYx2rnKTrv/RtcjXiqrlEiCBWQT/UIH11MkJ
ym2ojEqe9EWfcPyuDyaA2pBTw14ZfvPmZWQ7OK13pMBub7UMS+wrDzdjxKOR5a+EMrnOxoZcT6tz
5iVVlsuiWJaqen0qb75Mti3GwAcF5p6RGsxm62ZEGlMsmxBsKTQ+NIE1mJwn/uPP8XqSiXZFHuNa
ascyAfWfR1POPYCsxGF/JxazwCBV2SljI8ICc/NnSYXDAU3yugEyf2CFzbGrwu+/QqcIWpY+wvu/
AQsrFCFiSzjb9/hXcRf4hSKyAH6hxqcQOsY3mmOH0m6PYHyqjCww09bYrrAFBK0afllJBzWAAqmO
ZeNW4/+WzrB7kkhbtZ2Bouf4mF14Y61x1ihQDE1BRJKZCTA4UKtydeXTPPUnQKRKvQbapxljeOdb
YaYhNtJHa48XBNyI5jXtKhYDCgu/VJQDMTvE5YVJx83xY9xMiVE2rlLsxFbG1XCKxjRjF6dEPV7y
UKzIA7LiBhpjY41ne2lnht8ldM/3APbGGoCAnjgq3YWEzc7ky+fkIymBG8GEtJJQmxNAdEMXkpLf
YTicYM1jKb+mY6eJOr+cDsHVQus69KOM7e3pGfqgHYVPricHDALIwBudaIgCnW0RyKCBVhsxMWYn
WNcmCfLxQNY5MfMDIIKq5szrfuU2J1L6wVRzISlY69btH14CVmCMun1DAsPXDnOdQkT/kh4Leqje
iKLjV6CbHPF9iWRlNWteL2LUsWQ5TRj3M1BcUvcURp1x9Ll/GdnP3XyAcWNECWNR124Gl6+eDLRO
zUqZAFtzmrEfugGBIaUqqLaVCghSEoLKMYa8l8BWwvU+xiVwzXZEQNpnQfQWR1WzMINUxI0MboUA
/uwHmhDvTw4oC/HA2nNCR/V7aTzkeb7I/ClvF0+sFXFSinfLiOe4XjE1bwtbjQVd0huDxc7uXdeC
nTVGHEBZualmdwpSx2s8C1/mt5TSS7Io4r0uq7jNue0milqGkjL/KegC3QpLbcuwrMoZIZvDqypD
oz1ixHeKlgAwY6+2z+uT8JOhHkYC64maox+HisTGWqEnbogxfl/rWWlglVk+nQITXbHVXZUh1p6/
b4mlmI/ZLHZKNTkfUI7+g4vDZrygvgjg6jWXN5kECb9XzzGgmQr0M1qGrOO7w92FqgnPL0TbImol
A08w1GLVp9iFZ7wRfbCOnR58JXYEDDLk9oZoBa3WUTyKsVOH/0SlAptlnopNsdGlEood1YmVYYxM
DbET7MO5GTgWEajYu5aQe04HrB6m5gosMWpTVdvzOTpAEPDj5v1+XDLmgKLqK573dJ6xMSzBlywg
RgnohWiUbScKQcu7pgH74ReCETJSooDg5axmilPFIqN79mTBB0WRfJ33qZnuzJTtFfyzkJEiB59f
uII8fOLDybZ4QvSE+P0DO7F/otyZ0+EyPkHP5bHCNw4AefN2Btvdc4xKrjEy/3b3RcEuVCN5zQui
CMYX3jSH0NVYtHARfHznvCBOUu19M7q3lS+c76ZscsSI0qNvPJnAzfIhc8XgbhSWdEFBY8kFkr56
RyOLYXEmM2kupU5OU2CAvpr546YlgKXCalt7Q5dYtRM0GP3SUq6QEzJEvKRYXHMdbt9XtVKNFBtS
9ZplYrESGBEqk3xc+RjKFe0ff5P/tpGhgdSstSpxkQsSsyEL1FAGk4PHL45HsfRoK9hRnkohOQCv
za/ZdpHsS7vC+/ZrZH6REJo2rLjDxCPB4Kf4BImn9lBT4Qi4uWFqNJ2dxHR14RC/+LnYaDyvIxLX
frbqujmeq2EtCYOYQZR8WB8+aA/ZgyAuhF4eiOq+3mzxWgk8+NxSmcpCYYz3wuRxt+pbjfo/ltAY
rXyvCgm2qOGm7NpFAeKwq02+/TfJigQLmeE1KUV/aV1laYkAoV69WbtLe1SQO7+EiS+S7ROwYIpX
dx5umJHhwpl/F33q0571RO/6c2jQcvny+rZFd1I+Omstl0XRL0nbldQRusXaSoUnZstzeMlWksMQ
i8HIhz515dCVscDsVmDceAdyMLUf3DZUhqy4haV/BSq/IvWF5AC19h5dqjr2WDP56/uvh+wPwPAE
mf11orHSHz0ukO2bzlbtD0QveWzw+MHXhXoBaJBn1KLOhPJjIuRsHPcrAoMJBCt46K3gn3aQUKJi
rajRMH8veYILjtl8BAMjnol960Qfl/XRPOFXe8w0javsSgVutsPPokYBxlnsVGmq/TzjKBW5R+XJ
PDlb8AqxbJXQxDfCf4cwmZwHZwAzeCpyGClu755shhID8iSJsTgGMCGvdC41tkaNyc6AcoX5Yy86
C8+Ny0Dmmy+H7dKPdHI3nEVnR/KKVcDeVZXIKroTo6xM2pYg5LymKUa7JkypsDcV6I89pCPCwk20
BhHOTcaStrDr87IOwykE1fudU8O0ZUT2uSlUykhFStnSwX+qI6QwVs2DuLEq/nNv11CGM/HSQifi
13o7IoY1YdI/T9STfr/LgyUovpEApNNHJ/8C9N1jUX1DUzBFNKo8SzF8ewwYpXK6CZA8sX30G+No
OOGfTcXlI2J3OwJZejczzZB9AbZr5ByoBvc/WiL1YkxdPT+yxyRj898b+WeM66b0pUUb5O7YAn/2
xDCbCjmazvNTuJyIyJbqWc29FBqo+PH35NOqApuKNLEC+F1jAcX4IuCK0gIM7uVjhrp9xU+HX1Hq
WSPOW5nmX/qx1Qyccw0oxA7uTpOwmOFzZbgNvvj2DJG6sEVeCkupwtHl+ZvdOEdwdiuyuunYIDla
CZ0nEMWc1uNfMBHLOV4mwIjDGq+53BODFm5fRKAv5SO63/qu62gz2D0ecIDg/i0JbdDwqAg5ffWm
VnXYm+0ObDwMrmpl4+VgVZXrfVsHFQBarvTrRlvbYEKOCgvN5boQYfrz52LJ/Ijs7CE/Z4oqbeHx
SGnStzvDabKAO+zmAfB7jB4Y1K21SuKEF2yhHfoFKPH0I6Q7bpZ0jYvNvAu1NfgAgbI5UYvbjSDe
5MMjyyoK6uvthkk8Btlsmj+Le51vMfpAwsTULtQ0Ip+xB63tS/8xGoXYXsWzti5mZKfWqjfyN6NR
Fhyqzum7bpIUcb+UAXGbX/4sHJLmUvmQDTYF6z9EVVHj3EsvuV7s4dDgyu3U1RmWEmIOejMrFYc1
OnUCKsm9yvQx2I4IN2Er5iZwMe4wpHIU3iIRtq6nGj1W7tBHyJiX5fpbgAYpYG+0jq5YpI+TeeNP
SS/UpP3DymL7sMT8gpDnYNVf8TyCnZJXwtWM89cO92pJIOYPijG6v6uilhTIpVdrCkuUbOt1S4zF
leXPyVRYU2q1oIDEPbTvi3SCnWCQgZqn49P5qnun0KZedxJlrhlKp/EfFdMRxBXgK5XdaHUso2/t
IC2IyVmLTFyAgwxjT6N++2vufHLxGx3POfldP9sL36A8qCjK+TNg/qxh7PjQrNK8Clf6/q4aB7tf
cDlez2sdtdF+lSsId5kdj/CoGlCu+8AssSBVyCWtbKlAFNOgKJ/6TYhgyBJXmXUeO+D1NsXg3c0w
WlK4hFxtx5tPtKxQ/JdjUDPWyE+0XsEN9W/+0MmfhBsdh53xUn5uGb8dTsUd8lVmGrkDHaRaFoXw
Ru4rCRPUry2b3elHG4FmLyVNLptS+n5TY9+gpJ1foG4vkJvseCZvUqzQSpR2my7EajboQlm5O9Jl
OsXtg8vGcvkcZTPGyYqM6IZ0A4qT/zT/RcnnEfaPSmc1QyjLaEEnhGhLOOQQwqi4a6KZLv9afw8U
U5VPXWw3u+wZJPLBJQA1Gt6pFu3p4Pva0GTnipi1EMzLk0sECSSgrTBbM9RsWVod7Qq2ph5lGmtP
7eOrn9yAWebNhparEgX4g2fx805D/PjqOuRZgeitIb0qEvz3HcxnArPZFdfBEio+qgn000N2rGrS
oBeNbl6vXKVvhkxQqILSw21R5jQOswJDvg9ndaz05+2PTjNDBqzhGEQjaMKh0BO2weW1AaB021W9
Fv37QSJCMS83lYfknrhRM0DqUSHzG6YWpvhxzypkd/SAwd6SE7RWu8/h5pUqOZgkh6Rrdy/a4dCJ
j+LAgPrjUxBdqHxa9pIspXNJwlY+0o5On9dnepjyR4WABab1nql2pBoDtTAqb7+VSAfZxl48tJ+q
Y4B7kou7kL0RA/Syy/HHBlRYdvg/JYU54j4m8XB1wVKnFF7lLbFlgJgtzIXX5uJ8NkhdAawfVD4m
T4mAmay6Mfrjw5r3qcMto5LcXgGoewLFf25UvaEi9M/YgSzYkAXxnI4M/3T8k64nks7vnz4fQPm4
Log0V74rSWHnmroqO6DPc4WMrUH4AhaQYEWMgjQvrIFo5UKiClV2JWgjRtYwYDFC8jpfwoIa8zQ0
As+2dxQgvzXjoH4N5auZ/VvGd3vz2XS+C4B21OtjZEJzkZPO6TTQ/zNxRH4nkd+G6Rlqd1mJlW3N
+ft1nyFVWTVIqgZriUXqZ4BaohhyK+bWclB9tcFVTJRxDz+yU8kZNTLiQAgEqVLZLkjTIVgh8AdE
54Z+lTC+30MK2A2LKcVpZIishwkRVVe9OTLnoIFSElHJIuggKY+0dnKp5aeXCTKtftmw0FbEgFOw
WGBkiPNoE4OHmTRJMLNehqeIhXohH3mYuJpXalFVIOyYuaI2Z6ZotbVC/A7cHX8crS/anWFGV8qh
rDKGJckI0qvK0GvcAHVISHeVftuwqWyuxTdsF2Oq1Kq+6GUb3tZRTmQ9PVgqku7LxE+iDL7rdg//
g5oUribONhx6QlJfRi0QA0Iz1i07oDvF91LFxI9E8+Kncz6e/JBtTHJn+NgJFxbJPr9FcidxyQGE
Cvy77qqAZ4KejDuB8H9ZDO3IZUQ2DhuXLdLHUBEVsrQYhNiz4wiM7q0TQVHWnobi0A7h8YB5+15K
sRjaMGyvwg+H2DEj47EAwa6WIrGtSNmcQH4qDBi0GG1wKfTU57Z+IOL/bMs28zhfiSO8pfJbvMtC
fgokZapAg7jnyU0vqmHtn/s92i9e2PiSAZK4W3HP3dX+i5lcRqzBRGRzuGpO/B1dZ7lBhhgfMmQ9
5gpf9LHFYWO0yW8kc8SL276zkl/AfnHQDhdxDly9HopRCFP0mHpHFIDuHTzU/kk1HWI6CEZcKLRc
/y9w5fmF7M/h1QYGpeL9UzI3g8TYApu6FhO9nOIZLop3prEG2A7rrrqy+zm8Mx4M0KwX/i0d0kWs
SxmbnrGBUNvnvZItNT5SysFu0U2xD9kl8tC4Ea++26Pj8z7obbeasdVh0WcPqNB874+Sg7iG5q4E
kIh7Z6UdO/zYLt8p3oCEOCvxiAcB2aMez5Dw+L0vY/ErUVTFRfHoGBo9+3hGdQkj+TOVdUPCy9Cq
zcHauTie8sMgMAOC9jXthtgyq14g0Sw4qNYcFIee02z2Ox7gPwMYaCLF8J2jghBcT4p4mbxEMfTV
4wJ1uuoN/2XQUC7T1zV2HyR+hiYig1ofTnR2Va5RFE5EH86oMO7AljhnoVGpXuaFpIJL+wCBnjFy
76ROk7z3L5F1lveAdwLBlkmTWMsrwiwRpNFhuKoOd3ZU4jC7dpcQEPC4ZkdMZW9fL6KlqiqmdK5X
lj/9rs/hTucN5e0pgk+6uxdEkxfV5Ep8MBJXhXufqY8VMEu4Cf839N29gaR9VlRcnSNu91yPS8U0
UZyeOB+m+CS+TscPeRrxBXnRGjIbircy3VB/gBVuedXHEAUZeOvO3xAxUf2xnqffFFeSL0btZ6fN
r/hNC1feJuT+SZx01eT454y42ujJz0aQALnXEeXGnIMiP4ChN0xZQHhahemhXA5S0VI/eSTZrhVz
hg8jKfB4YNAC52mloIo3hyZBRTsx8QX1HHIU8/od0kxYMJsgmsWDJpp9ZkPFkI86tnEqeo4JabLl
NW7uZ5tJSBxxoVeVbrtQc1ThpXHjcD0M6t15u10DHVCLZwKLZky/upLzHW1rDaUk/KasrgtAPHM6
4EbI04+3Dm2VxxBkAWGRnJF0ZZTQkH+dnbUCvCkcKyCoTEtmnDsO64PRDntZPKC4YtRwrGQLaNtT
3QXJk2iamj6NTnx57Sm8N3aVE3RMxdQnk9NIo17WCSkz3qkhYIAO2Q5B50t/pl9dNrEpKoCaI6Tp
T+lM/JHAG2JWTGY0kepBZqnBue8yD/EjGaP2TSMEKCD1U+SWmysZWMskX4VEP9IV9Ngqkng3OGLE
Fq2Eb8t5ZdhZjtqt1nCGQd5G50K49+MlDsLd4RO9FkhhYMUzjxxl8/fMHmhoziDrsW7RvDBTpJ5t
V42cnZhlXYScC3nFIi6LnytRb9lT0ogofSlRP3EvAzGhgBDMBrS1jfx+o2oVXOM38x+FwvnMFJZI
jInuval+FOgsxyHb0SPThXLOClRE0ysqcyA0pf5CuwlDiWdOa3QhPF6qDnw+qOr+NFVcKRcQZOGa
Tx/WiU5fIPh0lLQZuX66dEAbUOdFn/0+QdYls059F/MUDhDTtN2+5n8SSB8lTIXojJvrX2U63KkE
M6uJObKnfsHAJ7FFVwTZaKQIS+X3jKJ6WosFfZ7iXSmAdHH737P9BEi+dyR28NQJ9O5ZLk8GBVNi
1heEc5fDIHIP7an0yigVF0SKZqqmJ3DmmA2NQ6tYXx7aTQh91BigbyVTP3uONOPwgvGl++IQUvAN
Pe+Ik0b+hjbTvOChjrsXFbJ8IEjUgtqE1Kg8DSyv8jngXwdvia/brDC9JGLPY0sWbMrmbSga4yq0
8lYKzo8aaETkBScK5sdeSkJcPMLrQo01kwiEV6qLXvoZdR7lKJv0LTV6kZ4/3XEpB04hqvj1O40W
mE5Mi4jnVWeuLMChjh+xKhoULHkTMS921tWNKQ3iRBLn/UkD8kdw2F/dBxbfjHvQqddk+DjcetBs
5i/NwArz2l6CNwErlq7bYBnsPV/vS+vVRGMGN/QB8k2oB5YV8GBorRvKZrBtPNMDDb7FVBt+Qmax
EYYPOCZqbfxCC383XMHAmO9vc3Gxy1ZnNgz9vA2+MEa/am7/9f7u1ZFsoy3MiXH68+mKrXGig6PH
zZFXca+Atz/IdFuhva8UMO5C3oF6wDBP1zxlYKn8QnfPZf57GC2+RdHMLjQOvdIP125jeJd/jE2P
0dVx6keLMiRGqz7wic7wdatM5uBK0khGGJzKEeA79idE2Xnja88U2u/hFhF2rE0yeufTC1O0DGk8
w6vH1w8Ry5gdYzJXs2pjyfLZQE1RAcwZSdJKdr7SyPkKc/AerRxyj3gFyoLotE4dcZuYxz6/7z/e
gRICYyNMBabwW+uoFiU0nK2VBA5xZ1T+tQkXqCQ+rmiCtCjqaX2irp/MK8cw0iVfrE7dpK7VaIUL
dXitjwmt47FnRlj7RU9OdbtiCQTJlSUgMzhML/4uP8zf84WPfIX2i0gHSHWoRIUsJDQt9rf8BJhx
03knD3+rLKyyLh7QkoIkkaYGX6EUM1NUcXvTlcmo0CnqTEWRmfJ5RrND/5XSS3RWbLtlr7fKVnX6
zDSJdkhXgAhMM4Z/NAbDmVwij7P2FLFycHewMztBKHdsbzr0cVcEtfx3K1BF2nkr/ZGVKsnEI+tx
Ruk/4NoGT70gJUS2ESwTFOlDtviou5Gpx5Xg1iR7T3PHXXHPoa05cE7tcutOTy9sId+fkEYsDmnN
HtTioKAvqn+9X7qBkfSp12gjmJXR5v1G7OEfrsSbq+vnlpcyJYNFs4p19BWO/MPKyan56J1utoNs
NRekXgotKa2FUffHiOUdzLYA7lyJaBejE6z3qz1VR6zcbNTFkb3MoJmZfiqN6WlmKJoXcx/845SR
5yukreTGPghF1FZGWPreRiYTeJ9JENZ/RZhvmKt6kZna5kwWU+6WwUjkAdG+Z7jTbnSx1IlEcZGn
+oKhLLnk8yWrxwUxyeMDWnXZFrJQOnHNYXCttyBR7FdKddrVYnh4XMGBT1hjgqBeUrYyL9M94zol
VOQ1VNKXfOAJbL35rPRwLVR+xupYU9p4ckd0BKQcVlqTOq8mvVvNCqFk342On3YKIcEc4kc8XPi+
goULrXhVcWdnpIW0jl/MvWLLrVq8yKcvPfzbjpEpkyAhwQ/WiaRI2zFK3j0o+2g+OOIXZKJeEokh
JFzMvr1oOgBudXULJqBuZV7v3BKC/aEZgRqs3Y1hDQj1NP+g7Spwb2R9X0dzGyYopCZj6T1p0j0l
fnxBCsmi4CVVsgcWDgYo2RmMw65C6IWHwCZUJTujv4StQfXbjHo6AR9xer0VczgjBGm/bJIXEWe8
MCYQnvHJHG9f3u6qpldkwSAn+2Ote/iqzw1Rjiijw8/4oTNSiNxRqOnHCQ5SujnxY08YslzmNOhD
dJQeGlgTOIxD8SSADw5Q7XjaW4G496l7ndv16LI4dsH5b+EEgPS6FXp91qwBNzIj14KNZ2a9drDT
Q+jCvqeczl1qU0LCclSJ/qbkMxd+7QSMujsa50uBqchlBl70D4wjn622HDxFvIEyUtzsD8S7Z/II
pj39qX2SLkrxQU/cuvPHTTkSF+wBm6YsoHuhvY9DYGR1kTcBf3AvNquWCCR+x28t7zrlQzyblGp0
o+XR4eMSDXtuUEKjIS+iBM1OXJ4TQmMUfxcl5ZPmKlPBTCVsemAmM88RI9Dx7DV1us2iCbfB+69a
yvZYbZOz/nG7p6U8TCDr/x335ZgJa516CDI8M0xws4kBuoNUjE0zPQkLNFcZCMMHL6yQjutrgEtD
JPl9oAJiAMmThmJLCXDCRbYAZgrykT1tD8+qhbccX3Vlu49DQ9hu74dk0rUom560PrgJSJfQn0vC
VFspZcRO5ToVquXFF4n9Lz1ESgm5NrM5F2DZQVLSVyaOnF6hO3jtu2ES+K2hYVQ9jTTUffAy13Xz
fSAQxAakW1FCvvRzMEKFLMoSl5pMhWZob1w+YCOz/M15UH+UuQPzvJgXr/QJpxzXocRISvQBBLbw
E4e+V3fDDwvxrGWEiM7JlWjcurZHx79AziJwq5MM6ZVOpj6oAtp5WEP9xexnhRdk1DjI8b+wCz/0
rMWR8liu8OTsyPAdx70GEZjhKXv8cfmeMzsSAbXLUKH1aSJ8zILvcYzNscIowRzR51FXCcHW7Dy3
V0yckoZNJDNxGVK4XWWR21zpXdJimkrwmls9GaBGc96m83eb/D2/5vklJvKwuFi16YhFAT7FRPgx
gZi9IfMuslJCzR8HgOot4PpJKYIJBoXKcUWxD+8d5Kld8Z+hX40YetDJTNRw5bSVlHGM8HVBJRDx
Y3oAwcua+PIQV2ONmBPlkDc+ilaKEA+wtpW6tJqTKJK69YPX3SvkEJVTgyKhsihZ2O1ISshtPbNi
lQ0Z1TPcjuP1f8lecZY5LX8T+o7xa6ixafZxvl6ItnlOPl2m3idNjzqoHoSJNKl/s8YLcLXjJm3+
fR1CTljBUhu+S6DPk3yPnuHEXDm+o0KOOiecd9FsmTLxeg+ShAHE9NfuPNt2I9xvjR81W6rjbW01
KBExS2SfA8oygiP+wKkNqQJDJDVOoAsAmHB19nJk+83T1O95niwrPx4IVczxAxgJsNXT3/ZEqk3b
Ys4kOwMHPDXYSKMIXACyvlFxN5eTiL3dhvzI6kRFruVnrEOCSgfNOkX9hXDy/gZRiiRYHJX0LY/U
RJ4wJqLDiNjs8uLFhLbM0fKGBNClK3BdaZE3lxyo5iEaaqlYbFoS7gxg8FnaMzmVEavfyf2uQ1gv
0pj+nUdQP97+svenqxeLhPJBom3L/rU7HFLNDK3UppUEjNFxjlgsWT+oZYbqqhM7T/zeNE6JPduV
tBCkOtzSU8YtGiEizd8VW9DPgJXBe90n/MDlLXkCVf0JVjYOtBtOsBSH8xBOr1+zRMhkXGR2wNW4
OEo7OEaTuH1pPbMFKE1rlGt9NCJ+eR+2HDL4nXzewT4uGxLoA0Sz0ViX5uqSb7hwvKCh8JRsoVup
/y45MfXQBBXQmUwqz+ld+41Ky230n87aDZUlMJFoHl2p+3bfQX7pHQSRyd4k1kvIWvzpURjjFytq
pB+KQwc26GYFXHH4yPy8Pc3DMCZuCIosic52byXIb4FoG2z56Z59YwBw3Vh2NnJ0/RUXa/9aZqG2
91wIksyTXnvf6hc5sN9r+fBloQV/FrTpa2mjOeh6IgHpuSHBvhGnYg5r82DtOxrgoA/jc5qHroaI
yeYqDXOxV3NBQNAYg7a+Awfny8RxOaEIGX1Po+Om7AxtAWyOWLUsbV6JMT8Tqkp9i1CJcwfOuym7
7Gv4CFJv8yU8sAz1onY0+cj7db5RsFHKd3G3GC4ePveopbleRT8anxz6mTT87g/03chmOJkCcIGE
hiKpHeHAuFXItBRWtQ89ZmXBCOhtK3VoVqrd+Hpq7JNuuwF8yk/1lcfMYi125AKZfxJJYmgRXalu
X9x7wXm+Jct6IqsIKbsBQKLTJecZhUNxnZUojG+fdl+FoOC+QPz+ljPDjBmlyGmO8g/7cJqgmC1E
TL9ebqK+M1BKm94R6o36i/ZkC8SEybhbh6ulaOUzUyO9FCN47RTOazBUy1CMME+P1kdfw98mb2X4
0iHMjwJjUpbIJPzST/GPoUF98CdbQ7DJW9Zk+Q0789K5+znC2R/G360m30R3KtOC3brxhzNrMJvz
DG61v5BXLFKeREjxi3+CJhHQOLaKYBO1YRo9k5pTA12wN4MB8McjP3bFtps93nJFMPACI59DnI1t
vtP3LJNpEmc3sB/ZDNzWRACkLYr/IpJQoK7IO4C7fOJqrpcoyOkNZuEl+zeddejmTZJ2dMraqL1l
rROFHJMIi+l6I4cHcZkCZ59fqWigLErm2KYUwHGMQQkcCna0tdYcIUugadaIlhTxlnySIoPAmdfd
Ikk4XD8e2SN1LuqDNedh49XGyWmusf+PTwYKA02PcpVNkx/s6kq1ZLU6Z3808oDP47QSXhewlJXI
Y+qmsEEX6h9LgHwlccDV3tWPhThn9RvgUiR386C+Yx59gw3MSFcSG9754w0dIU9ijuXDRA/XN7wf
rVUW5YzDi4dfk0vOryJkPvyRnWkhO07nZ5Ppx7fo7ullcmpvnahCcSu0jI09WstBa/Z9xulgrvQw
JhNQ4gxQ6mB0dKgyE3mfa40w7bgWF28bfUaY84sRUBCc+U0TmX2IDu463rRNDRqMG5+q4tBwCzB/
P8l5LO/7tkzCgdcE428FuvP+83hDvehQAhsNJaEsKca0raW8LCBwFqTGB+m1JRaJJb0aPNEncBnd
0UBDjGoHk8RDBRBOy7nIUAGIgZUDpfRoxjM6qprRBI0pNmOaXustTNFwBMYemKT+wNVFnwxuD8cr
YKFpwO9ul3IAt/CB0nJ/YT6FPAZXvStXNnpR/XO64w4iXhuVyNbm+KRv0OWERKMKABlAOVwbN7+1
4S6L8Ko6CjVerkv+gBgPTWbASisFiCjELiJ56U8Ml/G2348+K9grEfNYcRqx5ul5oyqF+HtBzt89
/VOZpadwY2VTbH1A5x2ZRWWF7qwiqjBVjTEjFR4tgZ1qVbuDxj4mH6QBpn2etTM8npMDg49skC8A
GFQMqBafeUMUyn6hIZCrD7u2URu1kFZoLBCVSwA81ALKkIFcdIufHe7sO/NJJ8dKs86sWpGY1JjJ
aFU8gdMgNkCU/R8wXIaZuZxkDFHjXeg6b1mwyNDbD5zlwub0SxZE82BFRh6h0qDWhJFRnpBUEoR/
X1dCGYRIItwSmomD3VGX/+SElTo+x74dA9h7IVdRYWApDqYH98PhiYn5B00nBKPTQ9ISNF9Yvljl
JAlDJIxWfUdNJoURaw2jHKfWdpxmRsY5SN63mPXcGOXEAQZIAAYMHL68QSLEtjLvZRYXnq5st5tF
RmTZboxWEfa96s87bFo8oensPYf21R4614q/GeC7wDSpKxg5kvPSNoCnrz2P5y2H02aNc8S8plrP
n0PJ5YbbIeqFX2ffDh8rgw8pvXIfgXvwu7L7ofZ7Q7s8vMil7A7xCiLEDoczOuXy5QexLTlzXB+k
h4EknyxBjjjeTExBF3eUaz/qKx9kn3FdYN660W6NyfPd0bj2ltcfCpvM02JBHTKm4laubFJKvjjm
Gg/PmIUvqwwjxYHGFbbINTop4lq1Ga+VihRjB71bMdG+IyIVAMJekTKW067J53nkLVsId7PhY+M6
uRJW7JVbMZPQaUIrZU5rbDPpUZwgH2mtcXh4EB7xhsKpY5tZ7Ctqt4UAdULXLKQDcFSeTU8aMBKz
W6eskQrQwp6HvDgqErbJqFd+bRdV+tBt/2YPAHyFptarjh5ZQlf5oGHDwQycc8Kv7IOKqDgmNPOd
TK+GuO5xtNsGpB7ZpszUP8kt4UPxgki2zbCKYInE6qfL2x7T8o/uLTtKShBi8+vSnIgIN+xOFmie
K1ZQqyI9CRYyH06z5kZ6CQbUEOpmCyRwgJZuysiHqwD6bOUwrlgaTopSODXxxjLF4t0pYAjxpEUS
0fzQOGXnGrbed8XBs57ksxUQSCQUPsiu/DrS8gcqUvo1WXl4dS1cZrJOli/G9fjq9r5nvrZhsX39
24hnLDWzCjS0joDULOSqiMBxgUTqY2TkDFigG3aMk3AU4Boj5MN2dxSfhsU+Bi3ViOwYJjNxGk8u
5MeCuEBKyaUmurXfQN+7rn+y//gT+8yyMqPiiCYsGg0u3+OmTuutdjxC5+sQ3Q+6hShTzxEB80d8
QYVyLAwRWhyzmRoKb+6Zx2jgbcr019TE2/XI9EW15dgYwIWyNdrRP3vxwZqjsog1uFkfYzDtn6Sm
3/uoEySa7A93Ckg/vgFiktBVH6nDPWPfktVpmLXyyw3WwRqmFjUcGQRYbfDc/0uHPChSmybkq9hj
nuHGKgHoRFs6/DK+bcGbYBKyv8w2HD7nO7NSXvuFGpz0D8NS4HGR7YFrS9K2XFbxfMHvKqH+nN+K
2HoGg2CvTZBCqhPKf7lgYaTF7OurReUKPs6HvGNRe5yUBVTa0ABuuljy9DPKHF9LnUB8nOaW+W2H
BLcM1EOHldpKxcH2m/SAdJtv3AnXyg/WW+dNAESmwzvdy3/5kEI/O5zdZUIMaYVlSSulkHfl3Zwp
1s/Qh4WGmFuFcoX2mVlROaqgPqMvXq2a5DPSqiD6LfPH67VUoLh+tRWp5zhQ3SaHTdETgFeypzTd
DuKf29ia1jSuFxxn+zlkIFuL45Nh6G7z9/jioT8N3I5woO6MJqHHep/5aAiuJgZzo+Oo2kgNutoy
pv2cQ7rwvhe5TSkVuk6XEWQvgb+aJeN7LVNargEi0zzdgTBe/TJfu0UqDcYHLuNWZOOT1fAuZoz7
7n7C3JK1EiFXXDDvA04r5/0CWRWtSSE/8pOMukiLRzICRM28xfGhL3Ra+oU0e8sKvM8VfnXSBcgq
U//GBQ0UJNqU2JK8fs+XhjxzB23uZOp98bdulMvgBF8/0RQuoDdmEUJkXJntOH1JVDOctuDZtneK
CVs1oqBxtidqgaAiDBmPPgjpzW2JBBMVWQEdjdNx0JPt0lmTTvhy8w/9cY3aNOCPjNtl40ChRjxb
TqMzd/5Ry9cOAIJwJcmUikSt+bf/YBUiNiV0H/PZChN1ADMXYLX/PqedP9mbglANE57Kh/rlMpHK
BZwxpUJH0D6YJavhD1kq0VdX2WkzTcr8vKrcJrlAXzB/jscgc2H/rfwpbjXiY+pBFx9QUwCalTf7
DSykmtdap4eWrc8UpwfQunExqVEupCxdTlreykqYrqrt43R1qGOce2BVRq7yv4MDGONDK8Xrwhp8
A5uGiVWkGe8CIaIVmL0SAtGQtBOKiP3AJ/rE9MffKvcssiTgW1vvbWvkEiHxtevzTGxHBS+W7XCk
JL5KJV/IrA/W5CyPsvCOeUOE47Qupaw4sXuRBwA5wphJboGtwUjQykaX5i2jdP02U/3cuppAlOAT
2R0V/f2LuQ5mxriO1wZAP5euaRhb5A5S/EwmXzva+/FONJDBXXjd3FBXs0axx9FUcQKgLlaYdZN7
xQWU+QKjSvDfNj1m2K6poeEKvhONLRs2CQ0zJ1BpvGxiZiO/2HImtzDAV8FI7pR+5vlXcoPGjiYu
JL16BibnelmuL3Qgd5IneYsBjKFvskdxezkucUejTmy0LK9AVGETD2EinQ/TOe+PWps6xIQoEybH
eVshU5sQEk/gKorAtFoPmHP2EbKx7YYUd+whAX4T5765pkZ4Mv2yPh85EPw5ucDP/NO2fSA/S6Xx
i8RWGRKZY6oY3xM1ZjC2IEr3rArNk3e7W7L5hRSk2s3FQMFbuhVDMfdGaDuL0jvpoLdi0enD4w5K
zz7ny8DZ7ZK3tsc4qZP6hWVOVq5GKFmMaqZWPtx9Pqfyek14x6eCJFLDDQsMJHP5OT75m125tQZX
uyLWZVDbUQoUtmKN6THuUip3Osibj/bUYSg1LnanWHr5iYhr/u8smZZC3lve5Cpikw56dB21o8M6
uAXkuFvgJDGmx1K2nYcFsk2K6hxdMm2oVC0CMQHkfLMlzBeffuBRPYCwi9ODmHCAs3zimXibj/R2
J7FNzEuv5KKm14OR8ak8zc4aoH3T097rCfi+8S8mIEMduHhLgPNKzb2bQWYWvSILXRom8RLrUPmS
2qDak6U5Ky80a/7yJOMcyRn1STy8UxZunXYUXnW7jWrpgSV9jVX+ZK5wU9DfV34ItyF8Y7Hpc6MN
AeJ+5I+oZI4X8VNV8zsmR153HuNzzXF/kmZ+a4aGoXID75rEaQjTbtAaP5WBnT3CXJIQ3ur2uupR
RVyttePMxkQs403hga4iFtc7gastoX3CBwmB7ipxtaLdRbstC4avG2svapEXnQHK4CzmJS9bfWRh
9hP277yII+iryVPFi35ruIb6Vr+XW1HW4d0pyNqewp4Pspvnoa8L+dXf1SLuIEV5v+qr5fQReN3i
jo+FxM6uM8QinF55gqLoY99srNEASKFMxf4vjYkfnaaBRd4WvSi0doYmdfGvreKONVrsxzpbT7pw
Xcq0xCIs/UtQNSg+81D6gHfdWg0U7Psiaw7gKmNV+apRQFvuK59Fgo4vgBDju6UXerhjxIc40kCS
pZ4nKNEPbTkI6dZTsux2ycSSJaJqKbs9Qa13rzdshEdQxZ2OoOTTzqYD5e3mnyZm8PudFnBzwRO1
LhO3SmY3SVDk+qO8OdzyGGEqknx7uEL7Inb4gFS6Lcde0f5+fSBj0PN5J5I4MUMTJFPaA7/QP+X+
ElOk+ahOtVnafFggGTD/S9lGC18cOXMCf42aESm1dO2wGgV6yN1ST7V5NixNGYjvuJEK7wbm1uoL
ieg7PbnqX1tWPHf3EsAA5i1OO0tgCWcdsowL4+osvP+zg6uIPnCufv43nSSlBrd8DeIfoyz7LM3N
CmXD62dH8NhEZt0VRsNKzewD1cPvzbu6ePTTBxOFTQOT6az7kN9T7ZqR6BE9cTWrFBJxvCj+ji5m
38SYqse1vYg3ZZHJ8ubYfGdComTUI367YETIIFTklJEKkhLnEdXH9zIFcYMHItukPS23Uu5C/a6G
C5zqoH0YDwZah4ChOZ6k6bB9gT1IfNOUd3Wz/aiSbZbWyiWoN8GKqEuC3WVrHRwanwH5tto1PEh8
ah9SjfpI+7wZI0yJRBLsIWvzfoZZ2CBYsRHO+41ICYPrCf9gEih2Xgfxht7yx59+W3GS8fmon5Fz
0iR1flNFwoLoE2RaspjKRZMiteU9OwG3CZqCq+D0r5N2loYzaRYMEQDl8zbfM4ssiHL8kjDHmP0R
kpOTunhq1Mhgu25Wfd03Se4ZTlYv5mNkGLkjxZH9oCYjU0VSHWmguHPdETkBOlEBHHb+4PTL7pfp
iC0DGzduMED4nWFSYOjX7nFwV42qwmWlSE0BEEIgWjE61x7OrlOH2RPiOBaFOkVbZJjLQ5z30I1k
LCzD+rv5CCdvOke+x4oIc4VNmOCCqBflKtSrNqdh9alwBxbSppvM1nANl13XzBuDKJIwhyLjQf+C
4wy+fBm+GOt7AUCAYti/Y7606OBGdlyi9EeWJZAo2y03XT1Nrpoz7Vp8R1Zz5256iWS0ixVmv0RW
BeIot/eI8CApHBCrDG2F2nT5yqCUb0PrDg9l7EpuMkvjOfybgl3VgYNRIVgyNHpVwfuyhL57B9uU
4bb+Q9Fl6y3YnW67Hz06jvg8uLhRaRLtA+17WSFLpkYsgM7cKJ3A/jZtaaMgL10TZwV2rV8xKwSo
O7ros+63jNrHDhU3MDkilFbnVciam6BCLlKmCAPMZhrxfnVtdz3PQf1ROwkr3hdEWz1G9IcAfkgO
rov5ZOz/zsY7HDlUm0SkEIey99d89YWnCyZjU6vXToH/b/FquMKCXEfGDC38G/6+2Bv4H9Xy0u8e
0nDusRzdImn97g5i4Lsk8CgISF0JzVSHM1u81zttxV6OLLGj6E1MxD8ZMMhz4htULIOF1PTPrnMU
YkQKulbApi4j6Lz2JjMwgBQlbsbQncqItWYhFXNNfPKU2WTLDKrPt3t+vFEwEzC2MK9ucLN9535M
sBxMxHpI9hjPfdai4aWSYjzSBswYp8nl/BMSrRPncXIJFaXMgYqTCqTeIuY3rEaJPL96FVtaDrA9
gn253Ft48f7h7hAaYwHaFRHtqSooQppSuXWHWOVj10Jc42BmTvOY7AE9d5C5rEi1cLDPSaC02dLM
aQYgqJ7RmJfb5pmMR+Wg6jNdTaCSi6GyPFBUOwapizR0B1fFM88D5po1/GdZQB2YJIFL/MBnkDz1
TjVT3XUk9PL8zBving+ywEoZ5f32VedA9ZQJVLF5SqvtzRGBSD5Qp/3jrZ6Q7p3o+R5SieHraqme
5Cdka2RLbjREg0Qb0QJApBiWKrgY2TPkqq+wwbyTrKG+VVMWyGK2ftFLmoOWFw2CwymYCyNPeuYm
72vb9SpaeB3QFYprpFInnn/beLvmPor8HOK5i5o2oyURdmnpSUq1obAE0ykmVVIIiH4s6a2kQCKy
oIAysoEyfovchV/qk5zeUzJo9nTkN1ypUs3nZjf6LHoByrKzZQW1zXfnIRQO7zk6a0xiNAo48ONY
JgpaNBRQ6O+sAvLa2nfPgGrMVcBH1YYMMeMpQ9s9lAhTT/F1PHoVlgPJEO17AVb0QDw48XgzuT9C
jCQJPQDOpphRfEEJaZk8hLZb1LD+6AtPNWapXRPkYkjX5imu/htfHSumZ5i2VwhTv0EE7WYKGMfa
/NBzpS1Xx2fK8s1ncWRXVwGemfs6qnWrgCw8tw3E67xqyWbQKpT3H5rG/1TAfh53N4k7O9sJiYeB
qi2lH/07+/hXtNph9b7BQ5yzaDy8xQs/fmHSWhUWu8hIsyHArPsqIlG8DO/8RcPbLH9+F1+8IA8X
oAqE3lE/RCF5o3h9ck2JCszERbeH618eOlAgqT/ABJ9mviq6admlqjOQc4IA559l/19WcOxshist
M2r/PlFWccOM8EQ2nt300Qc+YJVKJRF5+deAYqkWd46EqQTjph+afbMiTFftAYS/m6rSABScbO3T
9GS5dpOA7/QocppVOde2nNgt8rllHooVkAv3duYRJ3df3WxR9ZpQvYdCE8gk0oY2lkywQtR9/xH/
5JiykJ+EbC77XLv2QVhBnmrkAaPMzD+rUmPpONvrpZQV+Snp8DfgxEPUiuvSrLYGzDrx1GAjXeho
ZAR8HzSTgUZ3DJQ6NkEb3QQzN8V2MG/MoTVGyDk4/SgcGC7DAEUdaE7qd85WtPyy6EMFKBvzdHo3
ObCMvieZnshzPNDRVbajD8iVpgMlvJ+AXecS5UfA5CVUbs3IbQ80LeDFv0Qrm3IeywU1cdv2JPg6
gtIpJR9pAcol18Qe6v1LZcnr5shlwhdbMxONgPMfwqBddPiK6ZDUxe8pM97n7V6hykDul1fCfMWO
pCkcp+ecboqvT8lhaA+AFCN4LHp6pxZvArA63qAseTzb9z5ITjJ+9do5WTeg3kytnjKQ3B5PJyiL
ie+q5c8eByimJziFtGo22Mjg3Zxg1SPt/XoI0oYbqKym1DMoDThvUAqKDrTL4IewD98Ci8L3YHBg
VMIfpP6U+Rtl+CKWM/7Aij8+uqalmYdqbnmT34ag6QrTbVUPYBz15VhgvXios9OUJSnE5pfylNcg
im1XOgkYYWuZd93DeNTdydbhedyMd6SdQ0TGql68bCE0N7d+yr7mP1yLF90s74edF307t7cWwQad
C3d/wS7QV17DCG6k4q9MwQ9RzcFymMhuQqCJ8CkFsvL23zQCIQDWUxg4zTw0s7T+M6xvVvn1AIbc
Ux57hT6VnrW3+kEbz9xVMnB6+5QX0jvVTK0tKsIMP8cPwYpeYgAfMOP2rjaDb0n5ZqV6DwWpwvWZ
ax7TfHdxv0rxF41mStYEhhCoWIkQPicBdrslgNE61o5UdATGQTRdTTDOA0Mz2K7gESDFnPGRMBmP
PbaiYL7jFGRPo0lTjS/4dc4DrGThzx5BOhOCMejTCw9BOsI6LtMwrNX6zFRrplDDUkScT1zcMspH
e/uV6IED7YQdiPiQaqS7LDX7thPZX1wunQ1U2ybR6gHZ8mqxfJtkOrvdf6NiWzgLmaO44Sktum9J
jb1s3A9n7+6c9j4GmTcer56/mKZdS+mNbOrbXSPudrUbcFxddgLKl7NSEyCwUgv1suYuXE+TJljR
p3WIjNDLNFb61Eq4UvHJ9UnyAQbB9M+pbZHHD7Q29s6M1dgA4rXKEHnLSKbkMBMYxzVQh2nn/3FX
gZll/Ko9SR+SvfUET8WhB4wucF+Oe7TPkxC9PccmpnInP5ONxV4hy2HNVv4aRw600R4QMnBeQPxd
jOGqvKB7YU9u5nbQ9nCY9bkFJ7bsk6HlY3lQz68jhtOTX+xKKshzgkgscaMaJcY8QRA4sUivYlU1
sHiDNqnFkZgIldRHLcvwSTjRClMj88zAN4tXPpZdXBEs8CHEtArzGriRI4zy+VjGiuOb+nrgashe
StrNVd4C+xAFqwYKobgzwoTl4ylNRp5rP7aM3SFTY7UNwdZwtxMKfs4XbNKNfOFhnlxDCBhIc+RH
15+bI48f1+nVCO+t32mq+Y5OhpsCVDW7p1Hs77BSLuA0Y0lY6F8yXPlPnEWBAPyztasju7CfcFgw
H2LLVwYVRqeoT9zGJVk8BxGGjR62Oi8iNUftGSo/8H883o/CB6tn3RYSXECLftYyTEN1hz5sN7Sk
vK9z4g8z0bYJM+WvjQ3+p8qoJK15bw+TXvLS0bOFH4VLOQK7M7gnoWsRsh4LEglOuMhanNMwVWtF
wErPLKxcZSZQ0/GhJ8BE+0jilfo3ZCITBkeo0lJ9MxZTZpkXy3hl/TbGi/VwM3NvMx2ORFP8HM4S
TLCJJzmy0rwunX3aNAA8lQ34XDumI/pY9RzdcWJyKE2uhp8hJdefbHRBqF4EvmEjdSeBB0V2H1vv
qPjd3dgQz8+zo8vTkVcQUDkkWU0AW0Tj7mEWb7k0zaZkcn9UhBLg7q3abh9hhUiL3gdq+CFsWYSJ
hIvCfgpY+Slu1/HnEP4bojS70lqGQQB7yKOLlSqgBfMfgjM/PBtj1rQQm7I3Xq/m8591XwsU3HRH
Nbju8/kpsFzxJXxDpY4BwHI+FRJHW8LHeTVoAccAAWIaOlRHhJRIHjVPv+VU79OVr+UKU0eObkGX
z2gwK3NB5fTccfbAv2OvCuf/zsLAI74ihvSHWBwcVGdyz7PSIcwx1S/KpgwiJ/biOFVA6N9Uaaf3
xcSV1l2pLyiMxC1zDGEbZ1AW43InDIffrYtAIxT4DOrZxKBQ/jP0u+KEW/gmwi0CUhwM54+2Pghw
l51+KvaQiPKwqe/Rk/6UEcBZef/ll/GCHtIhF8Rm6MhxMWkQoAnwSKyqCMIvJj790EGaTfteYy2h
Fpi/M2G+8jSGoY7HjJE31J5M0b7UEHeqcyPzovnkF6ExXFEiSH1XVVRbLS7myWPe4pjZ0znQOSDI
E9xHYu/PmfR3xzdRDTxHbKoZDqCzva2wnqm8W1x7JHiR3k4/+SAYmhiiO6Tr+NewDy8DI97Gmbel
rNo3+r1sJV+hKB4OieCp7Jvu2AWRo2+9hvvtn3SxbayR1XpsUBMDWc58PDJEr6FYjqQW04TPXPeM
/Qf06XCqCYBxXnjn6Mfar2Ak8j2PCe9triyWglD36Vsi9coO3zUfVfm3GeK0qDoA2Yumkb+pFJe5
dkMaYApukqVVQA3ybdhxTmNDSFGg+/qh+/653X9eDowFXjXr7C8ONSVoPGKVLvRMWGpe9LyPxjkX
3OGmyqFDKHA/QF7KkTLlja53SexLo7XcTXp2nkRYxLY4vu/3rA0xNXuiT71xZZz1hPBugAtleiYD
uhdtH1Y7Fn2oZwBoW0UmlXedsCyyx4siHgkby7rBqESDO2eHu82XLW9SnJzNA8OPva5lCI27m6K8
skbzX6xrHMeX40teMEq0DDzSJp4xW/lmfpdJrwm+JpTWO1wT+lXA5KKid+L1sWhG5oLtAmH0o5G3
WDbrjwHWKGUUkrRsvFVsVGbDJelztrzNlfUtSTeA/7eZlxZQuHZYO1OQI3zhVtyKAnzTzyIIpZaE
UwFflJAAosI8IATfCuNCI9QOxuTFj/3eXOm7AuEAduMV7ijIQaJNpzY0qoraBaQkeTov70oWxKaI
Z84raIae9wdfPPXT6v0qeTNgRYmEbSPHhM35HMSZB/Z10lrDmrY489vUVMRyljAVD6MVYPJnKQp0
EH+GEzTAXR/9LQiclqRzhPl7fWkmriEGt/FOjypb5/96RJIWM2gEx5tLZAGdH7sftI96MfKD9Zgx
gEA6S6UhnRk05u/FLRFEk76cg0EzDWDYI4TdR/Eu5XSMGh9LVv0jaLNfeRtjhPClrZcJ9+gMeJVW
7dSQbYd4mofMQ4C8hTbj3gXFO+iyd339MtiqXsWSw96qLSR3YZ72Eh8ZRByuSlxZtRwDHppcNKjb
iglj2iSRki6UuiunXlyk4fVU6w/NoZh0wHbke8LbmHr7J0f/OR/dEZ6ba5bWxTGn6btKNlHovZBt
f1x1bFwRreze3BjwhDK2sIW/LBCJAbrG/Gef16NX/qqpB5+CAuZG6tSzVeRWGOyFVHay091V/wOX
W3KFbiu6De8bC2XjiTZSH0PVNw8pImrw9Rzer+NksJMVim9zGRF6EFoWAK84+cA1H5Z9iO98n1Vr
iJEhN8CEU6kUkxFQglxaxNJBY+jbad0iwFDpT5LwfSJuNCO+Jum1VtEmNrKbKnBu7Tr7fzZGu+M9
+oZZIJViSCnLWX50C2ZzPYDPHsd/kvf09DVA1JmYRpk2/WYUc6UQhBS1U9zeIbdBXSidSo1AS+Fr
rdjL2lyKkx6Oe3cFpFkL4EDnJ+KO0ULdYmWRkONvNlGZJcy9x3fA1udiG/svk0xgkNnRxz7FcNUj
Sg4ykjjcYV+skoAxaE0iHbidNIWggddY03j452LhGMpAYdMkPbSwvDybOgELmPALW/54MvhYhf4U
foUFyw9LcQJf5k4hJUL0eCUGrZdTGDuB08AelP57aepW6k8ni1c4oiCdMyakJzU6jA5ktS4VjCRc
wLNJVfr5ZxLDzsunOc54NfiuVstLoR4gG0YzTlwdtXZKSeKCSse9lS7I1AEej1O2XUSV8lO1CwU0
NpaY04KrFuDeI7IxgelEO6XpU/1NHTtkUT4MjF+UinfPhamyzJXz7pcNmucC4F9ZomGaYnZQZfK+
v2SFX0FvQfbnsSM/JrEV2+qcUytjUtz4wQPzxxDwLUxs4+6bAsuPc/gwyTs//Bp/ezsB+bgRyqQl
JzCaXA/KlAxoqvNL4Jzt1635xtZq1zRkolzKMmL6BNopTmc3EbR1EcsL5bSrD9u0bB5adcxVLbB0
FEA0+iDISOY8UzE8Vlbf1VrOa4gUHM8eLQyYA7IpzH+959Bd5/ryzzEJKXfznt35INAlVEfcKrtV
ftkqVXvjnT6bCbtRoNx0bTyJB7gNkFmAZJzngi6uA5pVU1ZOCxzb7fiTUPBI0fW6/Ihreos4fCkF
qLC49AxaPO9XUVJp+bGc6gOgUPIP6b7ULs7SRbHmcko/yJ7wzCPD2AE/WkVxjqIA0hDS/Oturpzw
cMZ5GdC8XnrS55w98pdBTiEAZe8AMtYB8vW74LVoX8R94Uncux5fLQHfLjPbUmQF+gSybnJ0uBsS
LVsEMvWkPxgvI1elELwdhog5+Bx+Z5Do9CKz7Z5mSdcFPX84sTA49yPti9C8GkrNqej+JqW//1/X
lPu1YkvTTTynOnsS/MkGNhwZGVlGRNwXd6LmxzMI9lDOJdGBvi0opB78uV6ps15TSokPwq67oNAl
+hlZ+TGKWKox0Vl7oVZ/Th4elIJmSUcvN9Ukd5pgPpBprT3ti6fPeymv23bT5+qx+Oh1ioSJZ2OM
XNneqbpWaMvXZUSqOdPRvoRVYsXLWs22CrzgKGYMKFkH7ebjTVyqHn/VEQWaZ64KYeNZKr4VyhKY
N+0p16u+W9GRu9HsQuzESeqOgdoW8WfrCYodm7rHS9SceGuxtkqyDA0uSdkEVaedKhpIB+Pnco+x
MeUDVTfFZ+NlzzU6rjnT8xnTWL/DiUM+olwYaIBMzXqQh+++uTLSn+vdbpVJ6TuDHHJPF0rVa0AK
oNiMnHVrF4rJmA91cpTeUanmpR1OwhoY+3CWHf3uPyBDJeBYsATkeJRUslGbXnQ4/ms9v22ZEWLU
OshXNE2Xxk9iEV7H3v+88ox//rC7IbeblCflcXV5yvCljI6495K099obATL8o+wTAPQk+e7H0SNW
KXScT0z01U2gFFN8f7WtjrQWmriYcG8ZbquChsrTPSRGbPQcdWyM9Cao2QzrxHJxQZ8PAyq9ZPst
vO93ylirH6xuiAj2cGGLBpABGOZ0DASgrW/x0gfGz2aPumCD84xgYcRwCC9BgNEs6JJJwBghX8FT
vGcUCraZfUZAICvNWzElHcldH99sEV/QbXjpKxD796TBX7Zhfv4eMjntxgq1PAiX3sk6sOcOmQlx
Wf5tE6+lo9kTvX2+rQRKEEvAXnTY+s4Oof6TCTDzhZglLA+nSKuCxoR400v3DRMKmdSvjXF4m3Io
gr+lGFSjj/NpzxgLYEOL6Sj4Y4BP7ucqeGO4kMSbvZBEgi9yhHqc+sS26FNwSDvQYpQNARfloTVz
NR2I4XkHiwIoi9XFMbwY7Zau/U6BbUWWcjE2lD/ylpShyqpp12pZYj7UA4958WVpLMvhnpedLElD
pGbNkL+yRf2Na7HD2aPzE3kE6EQsZURbxB15WWxMLAHMyy/zg6zUmZGF5mxHsdvUMW8E/3tG51Xu
3+QIhWK5t+YyYdHTaMw6yENXKQXI/Si5krhEWx0WoFosCBsHb3YXjH+vH+0KXc8qpYKPdEFe14i2
wcmnKF+jeVPlpLWMdJW/1ho+BxcKWoq8NSrcgX6BjNtki/ZNpJ70sy/2Za17M8QPYQQOwzkD2GmJ
h4Yhy+jJPZ673uKd4NKCHk1NOpiIB+wHu/ScBgFWfy6REmm4VtSCZ5yLO8ZOSyyRkQy9a6tL2Pcb
YB4P8NbZIXQ+rf98dJ2Lq178ZEDxZ8j9dnmYH4BS0iFktnzYU0LUW+GybAJgnV3kYyGX8l2P4uqv
zJFXVrquZ195dRwNmyQJ1XoEVDFM/mneFXnIX5BnKjzI8+KTRW128ITIkf99EHGezFCGk5FeS0KS
qGtPrWWOaej9lmuNlpTlGVLKDIqSdhcpyvUrx+QLy3aSxhHTr3CD5xxmeOmRj0Tu8GAXfKiRBFUJ
gesMNnAYJSainTOjezykoGAvEgiESViErrEk7MymtvX2NZ/58TFKfi6ScITyeMuMZ+gamc1I5lmZ
JoZcyZ1qub2NpLcRFvvEOcqmwg1EtXGLdL6OipY0yuF03mDhtSckLFeuKEIcABcms3sXT77YIrHP
015z3ef/M2Mp9rZDBwmpArO/RyKXXKmjn6OvZp7M2iluoFXfvHnmaLl/qjMoRnl3BKNBjMww7OuS
ZJwaAMbGU6dCHEIZz8liABzAOZtoHd2rw9vt67qYKzG+6pmXw184wbRAR+YGYj7pEqOCw1XkeO/C
dE5ieGKfsB0bi4CBlal6rKrcfFwFidKBsZ8CRRSr7ez2b6Hs89wfT6ROH/jf22S1SXAkou9dIpC5
rYAEpgLnrn1gyN+5GB+2xI7T9U5FjZt22pSLSNAr4C7NSZRoy91I/KiJBQ8x29A15Iw8WZh6ugsa
l/1T29WwKLcG1xrtcUkjzovJPzA6B1wy+SQhOckfZ43293o+PnVqf03wdm9UwQF6nwoi1bJpXmh2
q866PWnuPqaj3Rj773AeslBZI0i5YerXIVC+Jk1qv/xVBfXlfNEnuX9YtddZU5FzhMPS3s+fiqE7
F7yvHrEqgoIXsDvx9xFxVwwhbKjkmXF7oRvHR7nE8s4SamKs+fEeKyuKGC8xL+iCyNvNqaaEa7v2
56YtLAHQdD0ynmYFiBypZ5L4By335qQJd4rnzw6Lmr7HtJtGVhFVP1sPznbRCoa+wxY8WWNU7GRb
ZzBO5KBFUjaCrRIPSy85wsEBMmkv7Rp0XWTMcuE//m6LW0pOjNoVNly1sFgSgKJ43ouQ3KjTG7A6
n7DgxueOAGr0BOH4bw3LO3evSG+sA+BPt1JUllQPPkIoFazxHoUrnfAf9ZqeoFL1oSlvYQBjQ2BT
++apPgXfpJcnNSWIyCmZE2agU5Hj2U/RWcT9TymD98/1YyFsFt/aaQSkruJfsoCM/QUQHtOlLy69
o+baSEwkz0AK4He9Q8LGfwyDnxXL6i4N9ZRZ5y2tuKbW/9lukde2OheQpwh1VM0YbddESHV1SHFO
XbdxfZgv+W2pIex8iarmegkv/3P3dB0CwOYVxDWXcLK6th8Bwpp/mLgk2eL+7CVYTx2J8+g0qSyf
EUygITa47WsgOZpZiE7LpsusX7ppeiQ7pSsFozegLLAI3auEGiQssbHupp7os4LGwvlCNjoEYtMK
+4dwP0U7I2aRl2JRafHGIBU3F7UzBCeZx87eSRKJifEUMXcCghqfmkoLlDQStFmw5aY2dzoJqdpn
6bVB5ltsb2PEvg7QkhURfI1Z0oB8f7ROOPoBtyDYG981FGgNTfUhhKt4Rb6ghYkUaIocUOnqOsK9
SO6XhNwf25pgxTCKMx0aNA8lQKdYXjXughofW7LGOgsg6eMS/HCDu5i/Ta/HKJFjf28HeghzNwzI
9l0afBy1CmifiU9wfxGxJEnK1+VKhu35h0fy4xzNLB2rcyqLnFtmZqAcAxIz5TxdB9jbBEOHLUs0
gue4Ocr2bjiwy4RgU9FFev+b0XAvvCKyc5xe5kRq6b65O9WdmGWwCGttBp6hKGf8GefjkXMRv+Vf
hSqcM0B2DRsfexzmIgiaSt1OzDHnBR3aFDLolpm1FEA6gFVEZjv3HZ+SkZ8gGQTXy9Z8W2EbGH52
eY4pQM3NTioj+Ftnjgda6YjO5gfmc8nK/v2xkgwkRZREUvpzOySPvtt2T2KyRvXPY9D5LjA43D55
VwPGmpQxuZZefyAxcomhqzZGtf18kgehER/LN5c8yKk9e38wp6Z1PbMOfge8rnv6o9huXK9eNnbd
ciI72m7R23Ngi52joxu30f1UKXgMoyG1EWuOI4/DBAft2vdv10el2LAsKepRbEJgi3xqE+g77tDx
mxd4V+WtwNGiCiKAf0XZsHZFru28BKS1KZMTBbag3h57EnKyhyPmIioTZuXoeTeHyFZyj53n5yFE
2uv0nIBXc4U+cUu/ownoN8lRH5ylpwet857a8yhJ10oXnxAnYPPMhHy81ISpVvu3CV6ilejqK2ye
swWmf6fElS82gU9yoxJaRWac7uidWaDtd5WICUOEOmGzn1zzCzP3zrcirseyWX7pBJ2k8CJodCLv
h/nyUPSGd+3wX6Ox+j4ga8oShyTIfLLKPGCYqFeo3d5WR7gQ0v/qrjc+4SxyWlY5mmI6ITzPNE14
CH98ByyNQqMxCOkpH1v6ZmRYrVOfsZA9u8if6rPTAR3IuPkUNqO9CaVcrFf1BrxFJp8vdD4s5vRp
mDJTVrYQo9STcIxxwMAnamb1wQ6vMy5Ta8k5SVnw7XG7NGrZpUODVoiEGnr87h2mKzJ6MBTD8+5d
zKyNO0xZCb+hP/bwuWQ6ISoXKsWwmdwJMnNvkjp/OCtmN0qopZCWs+Tx/xV1G52NRECYTepjkwBy
EG+wucW3uSI3j9Sh3RnEMT6fbofDB+bInuOrFpB8pa0pW2e9H/HzZ7qNWK8SD7c0W5+NlgSbIsV9
pFU9BvSlPKqRAp2MrYJOUV3YYyriAWXEy3tt5pSsN6nr6uNL8BmqvptCN7uEe/8O94AwEkS1AmZF
npMwn6FUmmwCoNGqHIItJiDJAMCzKI1kOaej3PbodGjXFgTiQxXKrJc5ojw2cFZ8xbSvYCX+MxRE
UFuarjzE9i4dJbcMXBEOkr9a/AmpPsu1/7/nPGui3kgsAF4iTbSlqtISjDFcCM/irjuRa1aRt6ge
Ke0QjSevFAhiCG2I1TiydbiIjBEPAQdouw3G+tzKa5PNFL6QHiP3uPCC48YTKGQU2hJAlCFcCC0m
UtFNItISD82U3KQlMZRIwzMTqe1KmiOCiz9WE9B9Em7MEC9TVAkOqLkpSJ39qIhH0muvWvEMu9iQ
UuhVNVBHT6kAYx0zEI5FLm3Gh+mnr8CmJY2/lVYOBoJLs/GVApY6aNoGDikJnEHwhu2PF0L3lF4Y
TG2wFIL8LpO6c1y6JU/c2xU9N6/Zop7fZUvFXby8//tRLRqwDmgE+3iMHEex34WiDvZn75Q2OUwy
p2Smly24dgyoPT4UKVWqReJcaHlp1dbjYdhNCIXqsPb/sCKtnURI1cM/cIhf8eQf7qPdPITgMJ8n
a1dJ5M0DVIdoquofTVEDO+JGdZrMaS87v0LKmLJ2//q8dCCNnBc7SEqFSav3HhYkQNjtXRBZNFCT
7o7syd0eHqBlwsip6aPy3jobGFsl7N/87shIEqF1t55MS5cE6QxY0MM3eoDTGqRVj55e0kNrIf6n
aQU41RQLu62DjpS6TdZnLJ3pffe0yOTih8JR6pwNxb49OV9fvWtObwJeutVwYiD/pg8mQLaiUUgl
agXaxjqBgfOe3tXry+YUfB/p0lT+G289FAMA8BoItuTtfai6cQW8tVNAigq749KqRMuZiLeXG8hP
JFjVJci3m+vlRNY6gCB7+55z1MbJO4cPLMNQnqj0XWc91bvKqM6emhDSpBtYc+jLsT/nof6jqUaa
X41ZaXJuq758h1ANHAGlrwyd7/46wtmEjjOkWxzPYBvl9XWSAiVaUoVQsXo2Eu1n10ab5htbH5Ul
kGvg5ETjWKkwwmF8aqoioSokzCcHpHKdW37ydcDhVwl9cVXwhCotMh7MzBtI7iCaRicpWGNqX7Lx
D0RHBTr5X2WNpn5wkswl/R90VHo3hJ5gvsGv73dG8wsLkERoE2RvuhVetSlHGjG5vj1ZiWTUiKV0
gN+svXr7xvQwwFBm/IkzAvviWR5JOGib7ir1d6fR0w0QdvH3N9PB8EXfHQijy6F2oSEJ5RuLepd1
DnfC7k4np7serRUOjY5lBKPa5IWqveFDiKDSbWV3Uw71PNchyICCaQ/s6aTKcgA7a7k5I0704uF9
vvc1nfeQk8NbB9F/IUMEjcVy8GOcp3vcq4Miws00jlKstUDPlaRtaSjQ4VEneejl6+H/cgRSCm4F
c5uoj7l+OTDaNay7eZ62BsAXcSwL32vp7SW/ES7MyoQCihfI5fUd9L3KClfKffsrcq8bFt+zDfGm
9oZdbnTGrQnY9rnSTkvuoL96TCOL5cfBGIBGmsmugvMzdXpKcbwXTVZ92y71esxtdqET6QVnc5Ia
h2I+1FZ+c/M++B2GWVLNLj6Oi/rWW/MlfAlG7Y9Hbjo4uwlWEXFA6utTAA0su+ggJh3crEewwgUt
YJ4m2LC179xRW6JhaKfdBSGy3fb+JK/GdQGCEaOZdTyEPZgcRNDTuG24QF7GbbVRL6SUL3zM6rYK
ifK9uygx0HEZ9bexNB9XIjGoopNApzPGE8POE7PTTyV4vm1jnWZZipYdqJ9wbazX1vTQG1AF+c9g
cE199vkw7WYO8kjfweTdfVnmSQ8EfRJvfVg8dtj/WWPBkP1Iyh25BGy54+Lhw2AWh/qfmVTFfnQV
3ZHHk9/tqb4BYFoeUUkDLSI07MoSPVin680Q3jWl+gBEX7ZXVqbOwuaZWwb5iOtj/EvM+uY2Xg5m
5ve5mxOKiBlpNQqDfoiGiLXcTgb1Al47CsVDXZm4vBfhjk/9y2SHSCTE1l0IcpZxlu82O8qSmbNu
kzK9/iSFKWpxFKemhmTBLpp1I+BXheli1rjdxTgm+B7AbzrmtrNr0TUDgfUXt6srJRG7Q/uf6ZZ/
CEE+9O2rbPwlUOFoH7GOAERMBIQf0040nVCjR3qs0ylyo9hcnp9RPVGMto7n45Gahgeha45AjlVo
UQ6ITedYsoSHPnZ3WVsg/PFPac0O8nLQ9JlbOG3fP24/rSck4QvYHF6WXZfezpydzYM8N2pbt0Ey
eNcOJyaYdLfmBVB9Dm4Xy+Se6A1ma1UEYHNyqI/CSA4gfSR7ie7B611Z1AwC02xwtyXplkEYD8eQ
Hoq/XPfevSnjpWWDbXA7GzSrIbwzSg1B8AhQExg3DZEW1fwIB6QXyuVpIhtKMYqT7x00J73WKpYM
Piiq0hz5QXactmrlTq2wCYPoaKMbofLvfmD07bUyIOTA9aJtHblqvaqCzILypws7wTV+DvHCyW/6
6SDJFYeAl9h559LhsSC0vXKJUOzzYfgVmfx/3ky3DGjJQ5gOgECb9czH7e/Msjuc9oBhMrHbGnQw
0fFHJOgQCGdfdUNQvQctkyCrxB6L9BBXWqrwHLA0wVyAY/jn/rXt72VPzljkayZWhBgHKO1RjPAJ
x5ovUzyX+M1V0bgRkTo/T+KUTp8iUODWO2WrUcId1t5vWwtLKuE7GkbPqjvrzjKUCXVaEo3gWAoY
6uU57OzTwR2D1bQ6OtJLQqnS8P6PweQoJr8GMWPih3m66jQp/aRQlAAM6BNbEm7xZgsnMw04a0L2
VzUscJds/k5CzzxV5AIKxSZp41syO6ehEzOOhoml0mMNwGzMQ3shuVGg/KwXSGnmV3z3u9igDnps
OPV4wphNBFFLuFPjiYQTp6AgZgNHxIjMQPDLeyFhSUCGQMgj5M3CAUySMg0IMDXhrYPbkfiXBnNu
Elc7E72eiebuiwSki5xPM/ksnXyrWSlQde7t38eezUst1AK9ZYNDSBiUHQslGVpOSzi6XAWILiJc
4g2Wxgl5spJQ1m9WghC58oK3qJlJBRlZSdBJiSTJ6wqFTYoghEH5rYPZhGJeUQgBAyABuzF4hShP
IqxfJYHxER82oL2YLxPEqmNlSoEt9NPkGy3NsPMfg7MatZtWhqTgYQ4fp9l+FB9aAAudNEUUpQ1q
pMTRmz4/DBoiK6wdf1+G72QZ8UoW5F4vrKPc+nxga5X3Yl14wcVeICZzCqIExoEWR/feuNzTGZkC
9nGr6SUCdfVSCTa7wxqg29MPLyKhs7olpCh6LKhSWMbiBsQrpp+19/tCCOn/HwzenpNPDzeiSJXC
q456MputoySozzDVq6eIhQeTLF13+7soJFHVgLZoRyFcttqJ6zQ7AOfhBXrJlqirYGG8ctTk1HfU
QQGaKYx6Jm+qyWm0cKpw6QXzoGYMUC9C1kt1Ds0iVltPm2tQK8NzBW1jpnLUYG6dlf2Onuga6eqY
RvwnIzHGm9stiAcMBTAgRoWSjcdysA+yseFMC7skN6IAXKpuNt4lOaQ0sFRHcLApX6kukUbrOmj9
2FkdCqkslTbegZArH5piPOqhJppFvM0jAcgKO+TUK27TJXJ/kfhJyKP6QCgbsQ0bVd3QQEGOBMvM
hO1mvs1QP2GPHkxdNwxNAaq5OGoNIGjVTug1zRi88xaqgQUJguegD0ZDxxfwrhgm6cMWJzrguNPv
y81gC9h/k5fmp1ZfJHDeLFamPbIsoXRYbifhdo6G6gGC4wvKGCwKPBOfsc2uDgWNOJjaN5uDpM+r
zorpHV0xIK9u1Vy6qlnlCeitfbA35V/+GGb6Mp0bOlRR7+063hsSKX/m0ixL0aDLd+w0w8DK7C3n
zDM0XeCF/Wub/1PLUiyL62amgcOS4FBwrKK065CezvRAg5awzEA1AeL3LoulB8HhwZbjRMSYnmUX
eDhRby967i/iE4goXOyXZANlDQWF0+9Y6tQErf2aJvtFcUnl7IObVAyRvl1GkjCP9wWbooQd/+eB
qGxGCqWj/VI96vCse7xjWIbUXOZNmqCd1NoqEzw4llFyTJCrQCoQ7EZJQXvpms2ZdtTgE7VfGwVK
2hPXAwzNWwc+sjZZfTu3TtBHGrLfBqBKDasL4NdoZoAlgsNrXBbkav/foErqssnrPBXWgoNdCZs6
cU+xJ5xRVWO9UVc01KXquv1whZYZcdeDuv9VtSVWfotra0I4ZCtRpVv/HzsPWcaH1WxNx02HKC6m
yF4vsv6QyZj12+w5CJ2iPXWNv4n/ifAF9BccDrph66Kd+7DopSuLSnc02SCzwAKHtphzvMotyF69
5hBLXz2qVut7gxSN0514vU1laT4cqBbL6CcQOBLKQRlVGrADdWWohWzOXm5MVeRcFSDdPSQtA2LQ
pfy80tOlCtjsnmgiPuARQr+mR1d35Nu5CyCYaoigIDWVP9lFg9vfiuQQgGw14SE+jZmtJsBsA+re
AK0U6gLXddXOl2CWkeO1+R37/ikdNjgfojz7xEtCFoAAbNp1zQPeuigrPM5q0Auyu+cDmnaa5QxB
J9Nlauh7ETiqrvdK0tVLTAkR25lh9pVqq6umYgUfrTG1om6wA9N5wDeRxgGehD6Fw8epCucnXwVl
KrvGT7hnDBuIFWY+a5hHBHHmIMnudnCamTbSYPoiuNm09+KQCSHCwLvhvPfwRA6867OsNDl7bn2p
EMRjWcpNJy6hr+iiuApTWbrZG8sxp7afWfvrJ9GBqrXRS4JqSVd8DCTchJrHDCPM6liI55xEagYY
x8t8sPAmVwyYOqb0QpzmIyhFYrscK3VlpK591FvbUFYkJSSE0LahpCbuXxKC/7RgLu8tFOMXqwI8
Xtrdz9HXUNzbIBA1fuCdtatdRS051mjBdihJE5itIoiRGuLW9VrYv4IPNl5eAk6pKhLVstNNcEjX
FXHrupDfO2ufsqSCsmQUwUpV4k9kstw+64CkXYr3IoiiIX/WV0YWZb9WdsOsCLB01jQsLzwCwNGA
vSID669+teRRjRs6Ja/HHKdxjaTB5hzo//txQey5jiIqLlOtRLG62uZmMpqqCxPpAbHY7XExg5Cm
HTThv8zZrtT/RaCPDLKuNim2hF2Kyp/jmcZV+/A546j8V/mcTulqkWcXi81y1VQ80O7kyk6wcu3J
dfbOymFdcjmQLL7pmrkar+upOmmMgX3t6omQ7teLzRs28Ej0ZM/rkFjZy06JeNMBN1BuIGTc8g4L
kN4E5It6THqG1Ov/8mxpFdAY4MsI8pO3zAcfQ04HMSyh5d3QXo0n2J7EM+T2VE1p8r7cX3snA2GC
gmWR2eJQaqC8F/SBeaQaSg5Mry2xqzVHgvHUB+U/048d89YcOkDzrwLsU42TWDEnczLOkDLE11Cd
TLyrJzNivmkYxbLe3h5Q71m7iFq0CxWsNcFaxz5jbRMlRJIhK08ua8fpwRPq33IGYbbB/CfhkWge
0FEYxR6hTti1069OonQdsDzGJUX4Cn2HzR7ea+br7z5AdKrkSKq9NAN8SNrUkUYKBjN9BzstEVRK
XbnJ5XU9xyxU++R9k4Vjz9bAY/soeXumZo+ZgNpoPKPmixIYPmZ1vU+sAbA8gUEF4rNP6cq8HDEg
ZQcSc6tD5EXIo46e3ghovYRLQtg1S37j3lcMijO61d8p0HjV4sUGCI/FjDhVCU86gGSnfQMe4Ylg
PMSuc9Me8eOILi7EN09XmCcX+VehTz7yiv2nAPadiCW678F8uP8kNU28lIVFWev6lUkHkUJ9ZTtO
C2ZKfTfhGnXEV/y+PXk5kM7cxdujKVh0xCEXylL1QBmOutd/keiR9wGctuGtL3gJNKnHUFH/PRAL
I4KH53JB0KURaWtOuCD3bC8/M+amJCNdLSo/Q6YigJarV4aPc9IeSOYwyDlb0OfrpHglrniVZnCb
r3fcjX42zg1ldpDeVvY9EOI+3Fl6OUUVhMx8EB5hxNnSXKEPUSqhRlO9F1ufKeiGCCicJk785D6C
Pn+u3xLcsW5QlLSTO/EDnl0NsMBseaP1v7cmVUf3qzmV3BJvGCKE/wdTGZhUbVl+i138y17r7Q+F
RhFlz72SxsG/P3RDZkYZEHnV2gnqWGdfiqeCD1FmZzbWu7VjFWtkZpsl8nAVMp4UytjoVROW5htz
FOBlknB32FHJUI4qeoezTa2io1jUZS9ViC4UOmRRHVUV3RRuceIvs2xkTruhb7gUZspRjcGr0FCb
ZTpdm6k4UQ1SxqLB2uctd7E0RrJsVsFMyems0d9dF5Z5MAk6qrb5xwZzoNTHVvKx58tGjsUC8sqF
MQVsJxBKWTO3ZJxMyUeN1X1a7KUl52AdKqZt/iktkjy0P2LYobms15Ydms90XPU+XtbDvudyknYp
CMSLbGKxEKrya/dlt7LYm5ajvr5QIfxZ8WMzTclWUa7t+l/+/gR9xaHcL3liRSjUnh9y9jMfB6wL
fPaPBgOpkB2cV4zGbV2mnDfQtp2VHMZRoqR/PhpEkic00ac5PdQRGpVQMvyKuX6jccU3sae1IBat
Jl/mGkcSmL7PnvNHDaviBdg6XB5qMawP9GNgHToKJhk5Jb3mUU/x/+oF4d4xzjkydL5hpedxv5tb
YegTZWg8GBeoE2u06kXJpQmLL6S+NINaKdJGUvSuy86KQfQk0eo6PiB1TPJim/zWIhSD/djvrPJz
TAJLLzIKKxi0LgJWlH1XLwboQzOlhJ8tTDbQWDFt0AEveff4qyGoWHTbGtI0T3qpeb2fxpEPLM3I
Caemfkj/oiimXQL4DPmakfspWd6DpzWuCe9U1e5lpTPU7tHHQg8HJpLa3HuK+6pKer3QcmHx2/18
vcxvvKV/DPqvw1qHoZpMBLWP3eBCKiqiKPeJfWUGOzDpfcWUfCUnmOFLqeP+1A8ypiOlR6b81qmZ
OUR9BUAS8PqXO0YRQ4VVc8BMO0hC2/3AOHUKfgDxgdnsegMOebiH7yKYXCO08W5pIEWGnMfBa9hp
hoI+3zq/kNjOp9WGlgJ0Xe6Y6TAzu139Suh+uBKOLGoP0KDG/I2CEU5XiGN/x9YXYv385lBP4NMT
HZpmglhknZ8Jw8n4sjgzp6NMMjGKaX7JSTP1wlzjMmGEY3w7GwOdnWQ2Yig0HmlQGEVNvOFTY1+1
EM7vdf97KHstWLQVZQ75zhl6UuGQX7senms2rFgjdsD59VHaWhP8wtGcXFecvq4dXZ2P3/FUDxDS
rPrp7UeH4Pa2B5p5OAdh0qoN2G244bSSRSClZCz5TvIwxr/syKHcP4QNhY4oRyCGllCHhpmtq2rq
tHGMInz4rd1z+B0mIoibC+q6ac81iB5ftE9GJ6MWClHPDhh1itrD+Uv8TcokD69u5UoCTfCbquNB
nCgwPtQV7BPCPL+fD0T8eYVqV+FCokxLoSvV5c6LiPKgaODAzt008vQi4ysPabOcuvMoQ3KyBmIb
6/GTd+4LfBwAd0FQsACnxeSb3wtmexDSGXGIx6qvi/qDHDiMiPJtGZ8atxQ/AxxZaRYyPukxvnCu
ZhX4DGD5zGdJYWMz3xAFZ7s+EEpPgAyV2bObFA0nMtJsvHU79kgHbjSiZC0S2gpuBXzyZVPybBK+
0qi9GTho9OMFJgvgcAhJoPWb3ZazCt6Vq1mwGa8cop8rvKTuhhxnFCws9NI1bLLGQLJkAfT/MG9U
mKIFPUhTDvBb81MdIEQDI5drPpCtDUAQx0TgIjgIlcdbxIxrEUSo4uJk+QjOofTNnHKG+tsYRTc6
tx2VEzO087AGk3mHvpr6fAqTnTCHfTq8qaBW3pC7Lfq35IxljW0bNHP4MRWEQ0045yoi1avpb/RP
jE+z1VQRwnoGZOr8FCiEwN0XebcEkzf/pgJET9FgchCFwKRWjPxWSBmzRV67uxUzJ9I/d1H7k1rB
J5ggUosMBLgF9jPgUM+bCjg1skuQE5ZTaBt0eE84HtT1L6eaVYQjWlPvONwan6sT5wKMgGyzVu/g
yan4n3pawYh6oLLnmqgk2tN6BdFBJhgbqz0PiP2XwAvRSHkw3vyF7+Uh7czKKlsV3VNnoTaacE5j
ApRCHfIEr/6k45DKYSjsecKivQASRwvXGSi5e8BwKmNRrIkI3m6Z61v7QADg1iodLxLSYC+7EXCd
4Z064DKtB0bVhIu1g9HbrziIzvmewbz9/rGY3EbD42G3EotNheAW745ZFbbytkMPDJkPq4Q7bQwA
Ypm3hzwxyYAJ57SVfLWx2o6Ep/OpQhUXD4sFQ87J9P740FTM8HdbmdFVhpWYQRncZtwpULHcbmOd
JauLxeazsszIEen5k3JOLdipBMh1Gp5w8rbjWj09yQTTSOYOxTMuqubeTMJGeNzcklpzVwW3OGTn
bEmHby8nVCi+hJ28FJM4PZYfYlYPCVEMDUNjPOxM55MV6kYV1hVjp7zi0Kn8zPip8B20pt0pRhg8
/GHDfqqKJkKQGD8m3kBNObmmXxuk5meJZnSIKZJ4ezx79IS7BukyrsRw1izY+wE/+d6KIHHsV9f6
UvsotEYZZ8e/iaAcMk7hAlW5xoah3I1XyvZPUO/NgnNjdYiWIOmQO3OSX2FgjcgmEMAfkLA+DABP
9ZbFj+ymPZgPtRfDF6CLJN1j76XSzyCy/rTF+h8lrd7UxrBhHMyTw0ytaXtNS669Uku+0jF3FNG0
SFwt5polqD0hCRwoua8KO4R/HKx7ZsOeDJrDWcZabU1c2vi73yDvtmQPA+XzYOCr7cmZIDypfp3W
klhTq2sURxQoLfl+KFevPpjekvaaZitTGeWkUu9IWjPw+1qQVi/e+3Al4UjQEYCuvXjKddAqGYzq
+/VsK7V7OZRgsXpK+L1D+GAZhTcTk7xGYylTziVHVnqE4tji8Vr+wskTW3SHTFKTQ4MyyFazupo3
FTz+BdacWkxFgeHafRXl3HBiZLCPgddOnB6U0Vd9wV7+c/9XIv4DP0psn+SbnEU7h4kJOKQNI5v4
HwhbA2t45j23fm+yhxjCFF3KbMRMzNbiC+TcrMnIf+f4jDHV5YXNqUyp1MQXuZfArprLSQEYIH/7
6y/WuqF/l3EjE0EwjNvkEHTLRmGi2FAxM1dtA1RCEXIg10sWTFajw18li3sgKKPiidqvREyShjYt
efriNwI6PoFEB7mMNyS6VFUYbeP6uaA1NU3U+tLpoUcH/FSDGuu+44AqfKaA6cC9691VrIXxx4Ue
X/dtTPkjb3hLbnIowvXe06HG4zYujWqCC3slXEpJ9j3b9Fub0elfF2s8EviU1uy+8KwOuMLg1haI
koIKC9mFvIIPNwnJE57ZK3eWXEGizcYaoX3KkA/xWRdP+Ek0wqigRmbnlEBb6qR5P3uE5LRcZCV9
jSgegCnjUAUhKi6VKW/OPcqGZxRtCbAc1DC6F6YJPZ3wzaKwZqTlweeNQ/JAUUFOQacC+o5I1TVa
YBUoGw5++2gZU1q6FuA+z9M15I+Fwpz0tnBNwDM2WRh2wNGUh9mrTrL3kva18+Bp/X4Z6gew3/Pc
7fe/vKccdOWQeWa2O06/wWGTecnWuZR5ci5TpMKZ3nP+Z+RuG0dgbTo9A7hSpjLyU8c2G90LRk4I
QlT3rAwVuQD6zYgtCzfZn71DFHMqJSB1ov447ifTv0MTEW2naPlhua+meCuwCqPAnZByUUsEuAGj
gVvbo012vclMGfp0NCzy3nny3J5UyLkwYU1HLohIFoBBj1NW0aETyxEX+DwsDCIzWRX1I1nR/fgB
NFgI5fiqix48//S3GvBpF0l9o4Fe5baFZvj9wRRtGNIvB+fna6inKcfdzAO0F+0oDqziI6ZoNzMr
5GNVxADmTsctuVSqwLP8b3hQMjIqs+/r8lErFMgJBE+9zITA9zvq9yd0DEfZEf8NiJUBFmM4//Z2
jYh8XnsxaN6wmuxPeQMt7lfLmo486gmwkGQKa8Ic0+i3ivmO3+8h80vBBFnQudVnDEEiye5zOr70
oUSQ02/w4O4qiTcIxIgEa/oaYey4zlsINVAL90K02NHvQUS7qkm8d92hxlWYpAlIvWOHsV0JkOy6
wL7pJdi4c1gD/bM69F+IEH6pdsqAGI+V1ps95u/REoJf1c4coWSvXoHtq5ya9RsztjArKrG6ZtTt
Tt3tJiVoewnyxLf2H9zM4kMfTXpQOO1qp+OL11rSrUyxyheOWsYDhAjxAyUJ3NxGYnjw3eHCsROU
Qnbxp9FMeqUjtuN7bHly/nfPvFPqry+OmvCr98cC8K3V0N1J874fufuHQ9S3NdFr+JtosXBZtDvt
bgVbm+F7gkPcPeh98IPb2kSmM1vwbp+nJT58XbS2j6EoaIzNizuvQ1vIBnrkTAzRUw9/VAPQf1t9
APNl4kdArpIDkLu7YclCVvdU0jW8dKmlzF/6SiaAw9hZyz+eok/J00a2Vh8KddzoqI9Bqeh+xNmw
CP84k4SItDFlgKe/dwWfar0KmTY3zPx45ePwVK2qs0yvsc9yeJYSsbA0/TTYf8f/jYeUILgP2kv0
2340q/Lp8TrT0JdOCTpMJRFLAgUKrpnVSU6u3XB6MUgv/jZJLCeicaViMq8fSeWIxD8pPdvKrL07
UXwfdu/rcO0dMzSyrqPOx/zoThux8s6wpR+zmfg7CwU5mxFAlZ3aCTcxG/mI2fAaEP9LMTS1SWpi
zbciH6pUj0KVaMGeiQvvobiZ+y6dB0Sa/ieLmffKMqjhsM0hzGlWRKEk2RR3jXT0pC5IpipdneEK
l19Nbt2cwJnSLuK4c1y6ZiKVVdpep8nXt1ilIX/pGKrbF67tAZ0NrqAGcqMl4fUFqfcEPZgyaeNk
Sj4mZQq43Jdb5DrjaaEf41eLxPYM5kIOZPkHZ52N2kIE52DFexwUNmrWAaDcOD1EfaK+V0IW8nJu
aoqHO2LPvmY4l9xiJF0WUVRtFMGJMZtuMDYWOetm9Se6hifdQl0M7SpFya2AEpAqdF/gM2A3MDSX
J2LRIZ3JXyfPGib3yPcqIAfMY/0EHN9X0y7chX84n/IZrWAmv99tHKj83vjTMPMsYTrP1ue79AOr
yIe9SUU2NiJ91Q7rsNpCYaWRR/ZzNcNchXDXdbnwQkQIU++bXS1HxN0i5VsyD78mIwzTq8uYB7uv
G43/3iSGkCvnzEO2wXcb6HK+sENCqgsgWdrda7Sy1fVvJPPfYeLCwft4DMiYUM0WaPZwZvBuLWSs
wR43aPKHjA0JMVmZu9b4aDnb1BF6YZa0V1ZHCu8JcLw25iRBTs7I4oe+QmlhQ6KJP4UabNonTWhq
Z6KI8mtOSPGbqFCO6nNaifEDhXLHOrB0jjquezokjfkXeVOcIaELEpeCbgU+YX+Y4Y7R0VyGn0M9
tw5HLlm/Fc3k6TwrA7Ch93auo0isX0e/ojHjoZlcs9LH3SIu5tQvmUZkO+xxaA7LlLnNPl46Dliv
pKIIsg2Npwkox49Mq+whQ1hNk4EaOXRblDMSXaPRp/9VT4P8BxHmHNi0NyJS1rCSQfAfqBS25MCz
AOccZfmv65alTt3qixMRCizVkqHTA6L0//HPCoqYqFcw19i52hqdeApdwt2iAUlvOdqD9WXIAtdC
VUJG6kAs+HEEqfdqZ0MfWvkZtwoyrc5RLFBgZHPLBwYApkOmdBVjvDqWqxKaFoE7cmi0W/7MC4PO
ubxiS8omBX+HAPqHazhO+N6CSqXX+wozba/hbeC1zNG/ooQfXbmrAyqd4ND+75fuYmqdHz6BN7E2
l9sCO2lyiEVgwC19pHgP3TnX8E5B4ixWv2Rzh/Ag914pnnKFa93l9yMWyKqgbfVeXxPNFCEvZhD+
KAhgZ9m9FXe/fOK6E/VFnDqk5Oq9ZNxuJN4mB9EiLUBIUhHvlwLDVQg2NETuMplpeLn7KjS14r5o
niNcOnhxr7y+L3skHy9ZuUMsZKx0DSwOkfhCEPJwJEkH0LbDBZfNNLXegX0nAvt1Mv+3DEBl7bYS
dWQ9R+25J9tPdY8ffBHYTtoOmNgUAIeEVgFNWDuYlMP5yXjXmDDhWWryoiRJ07mKIEcJYdmUVWn/
YhjqqHj4FHOUuC2AEl5ma41tcgoshimTR85rHP+rrzwRcIV0Hzjizrcr8M6FCc66PKHBG6Pu53GT
lAlW1DNOwBz/qepuRhcZyeBWsVLRAUokPQRLpa/cKz0ImF5RHRNOp/su17qRzgaVVVAQAKnHCEZJ
wspYIhnOpfKAVWD5hmAge8IXKqMeq084tiKBmEMV9wQ2sL9Ss5FAu5kVADlIRJRVi56MprYSUQOo
Xmp52e+d99hRsFsH1rmi1lR0TFPjxMCD6sJS6vcFtZyfbmNQDwo2Lae5hSOmNZvil08DqFkrkUi5
X4a23epQe7hmMaoJ0yTWXVfdPGqmNBqi/73FAu0wKWHQCrx/41QO8IzMIE+MRDPIiXNAu52sQqZ/
iagPdMpiDA6tGr0A06mSgRaCpBth+h7Qkez/JU6/GMooscH3y4XvuqACV4WD5MyCuU1cLEsgIsVp
AZnOyoCllPVGUtJrzfxj0XHz0BXmLOqtwxoLpl1I8lPVS9YbXG38wIj10PIbmL+KdUQvkz18tf3A
DuNmyz3FV576kFgRt4aiDo0Bndux9VinraHHc6/lzDN0W+Rsr/QXtsV4PdV6Kgv4tQG2cnNbSOn+
Z3nN6I18zQTHYHcu64E/F0lCvWwvAYDpekhg95dnFTDQvCKMiM3ReWu4DLxcyCvgc4uv1sIS+mrh
KyGSDXXA/PY7RfcmlnFMI+SOz2cnnY6hNQU9+Hs2wD9rDp30bFV63f6ZadAFmWU3jPCe/r5dBvMw
RoHxvchv6I1Cd2cy1VgZNueFKuK9+KfmZtltdYTaje1AHCfQHx/LiujoBiEqJGeMOBk6uV1vkz5v
HHrJV9+IkrCIRnEQWan8DhNdgJ3c/g+AlNDTqMpZ+/FrghfxP4oDW3A6GBVZTx9bxUVSl81hDnyE
SANh2G79oe+pZ9pPyJNCtLt10ZcqkfmvWHgVUs0R07CkDj57RD11DZW0zOLPpTEXOasJY61PtRSZ
oApQDnKlZtTn812dw+XdPkMdAbiQXMtPKWqYKRjCQiAKVPXmJjTjyzcI2p4XNuRJZ8N0T6owJqRC
+XH5wnFbi2lIMg0GWthtLyFQC3hRW5uQk40ulf5PSsHx1EMBEVvbWXDpeBrJP5J8G+wt4460CJ4p
4E+36vSmT+4z9xgEE9J30epSrqwEFoj05p41o07LYMPNlApm0SrqKC6clFszojveX0Y2GqWoNce2
DlTAP+N+C/0+FdbVCpcSLBZqOD4zl5bcsTQs2pBtO1dNAPNz6BG7KpV1JbRvTKY8m+9kw4gGiMvt
ibNutW0YyCFh0vgWsm8rSMeRXFQA0a1Dorw5e6EZfWDLDYqbAe9zzxFmQe+7lNFGHRWk9wuNFuJ1
WimphiBOvDiNR0Skp8GR/U/ZCrj02hgZmAL2iA+S9pd7VCPJgCU8WA5jWLLFpu38bB3o7Pnys9ui
baoxC2LAwPTWQc9/kxU2B5KwloWVkKdYoCwXQBf0tFNZLHLCO9qHVMYoSeyF80IK7XLDt0ea51gU
DzEbB+Szh5spwII9kDpEEpDehlVT3SSTpss17cNNpCB6b8DfglWckHlimfuhNhpsEhMtbGb+AnpZ
5Marp7QbnwcGkLKF0IBlqkwes8bZ0pN+NOkhBNOSV62FGDastCXRcGBTuP0MdT0vwAbyZAtgDPUa
IN95COF4Z3eS1V//ai9rqQihVDpaG3p9T7ghRh2ylDBDauBi7BYA12T/MSNF5c4TyOD87gknsp55
4J+tBjg0pIEOsLxiF8PgE2Oe63M5sbZiscPfk097WfseOFi+rWPatO1mJZK5L4JPrt90xCRWYUby
yFOVYEAa3b2pQUaXEdEX0IPuFBHq/VOfVH+NIBlkXWRhIHg1KhQjePb6JlevLcrgT9xC7na8h3JE
K/WyLo8fgrGwmVvagdhVudCzEKxslttS9qvnQEVSXgU3zUFk5NKNlzU1UeaV15FB9rx9uGTOph/N
42FZO5WkLGSenMqNEXom4g+UCZoCZ4zf9rXjKmZwYo5wSBQbd3iWJb+znV80uo5Xd4g+Tdk0He1c
9B441dJD0SW/jo7gKePYBmSAarLgz6HuFhLdpxxksE/eGs0AAJqkamuSe/x01uVII1YjgoJ5M4Kv
j6PCrNqNMTecacDE76GXxQOg3Mcrkj2HGqK+pbGUEFFH4dpOpNzY4r7NYFQSbzqYYLb00jUWdiN7
q+rGCM+zCUTzDNst95So+2WnK4d5wfkXJHgB67FD9uxRpOkNUFARZt+7d74QflUdUQE0m8E6fQ1d
AbjACd/fSTkAWPpMiI13n5VU2UD7PdUPFoEmmXrZ7TpbVe1hhIQ1QgAbS5qQytc9LezCfvGy/g6K
Z7qXfkZZP5y/mAjKyw/7qMVCx37urBtN0/lY+zafBNR6kPKT52uALVoqQGJcae1lU9toDcaN3EsG
EZr3mqSDeWUu107wr519v8rWVJQQyk/4RICfp5Q5gtLaN8lgIxYjTaIUi/XPm2brQHVtRPjL7dN2
oQqij85OGDzk45Hm7u1KfvlyELtx+SyzRsmWdHbO3H82A13PiBlLyOeT6SbogJdSgyfIP2dtOBQK
+CjTTDFCq28sKH7PR9eSE+Buy4p08DF5KgQUwgHIiREUUzISmMIv2E6qDXgA3KEG2GgBFJGqNdos
VMFaMBl358mRe9nOb8savMQQu5nhfb4efbiB7/t5eb2KYSDZCRShmSAS2ss9WotKQbh1ghHXWwHb
12m+3NG9aF8/yw6EPQsvSGjqOxb2lirILA6F342DNnOCEpIsiTqiicNCnVC7LHLV6KjsgO8pHfvd
Vsbu+tPDrT26WkumufykT8EDh9ThYJ0uBj73aXc/a/7GkSpt9TSGokjfnD8HuoVouf5ZZ2JTAIea
ZsYjHHLx2LDaj+KcZwoPx+N7cHxvEjwUwZKM65rElAYCadDKFktR87xXZBM7j7DRMVyPzCqbN3Fh
25jLHAAJZCGRwp9CxY7JB2b737+bu3zN+kfo8eA9Ickvu0ATKXeqdsAoc7U27FamsvDvZeTUUV2V
Ic2chM28Z7tFsXp/Diy9uTLCuQ9xRU1/L4/x6BVfNrmX5uVct1cq8ul9caCPDkk1ms6fcqCV2zc+
VohJKkqn+eGvsYxuABqt+3pKZ/fG0shJeM/9LmuPNYfc0S0GCqxS+uNsqRDZ+1iEA1PjMWOHe65U
ojwpnZF4R3Fk8SRbIQKI98sAE/4mI56guIfgLkV7qWX7IA6f+F+d9mu6hwGGa7wN1xIkP+RIN/x8
6mChLBir/3TpaCxmGfJkMBNG5qElHrEWZNgIvdiSMkEPSq3/UHqMH0aHFDj+Wn1w0P93F9oFnR9q
PpFReW+zn1TDDTyLJASKYw4DOsybipaYAIVOGjHQ70RhInpZb+y5DDnRHyVu3EmPA6W5iGz12qco
Vq87BkxNaDhni6S2i2Y62XFkk3PtutbF7Uq5XSCkgLkhpaM2TvYVqGQAEX1j22Xdz2HQOgYKhosw
swNqvf5HwyRMJ4TutQEnJMrNEmyR5vB5V+hp9dCVAxVooXlY8R+FALR/SAn3Cv0UtSMzxmYlZVwv
VTYBdVyic9FxQkYp1+mHybLvWQ36/lFGtHk/QQEkiZdPAwzhyAfRau5vApvBDNWtCJEOcwGqO0Cx
+LxYnxY0+hMwLOj58+eVIzLVJbojg/EU7A5t0SO3zbIoErkML0t2Hl5BVq5Y5mxH86sxWUBD6G19
M8M36Z4KbqVhDgRNSVWq2r5P6xZ7pNThemHv+31THS3KJG+i2ncdiow06EF1B4qwba3KU8242f31
D///ax572GVsXsZv4GHtL4e/l3Ssmi+bOUnkcFPveyK7ixKnRDTa9OmcRNe//iPa9esM+CslwbW3
h7PHfWJS0Ip0urrU+TBQj5n6+E0Xc5nEGfJQ5Icr9voyJuRZWtlUcZOq1kuFxhUqWBmXa8CDwKrn
VPGXGssVyM8x7wY5Fuwdn9cXGkqKdE61El07eVA2KkMiIB5PQAx/QaKJQD8WRiQLIaivT+MiNCBZ
Qgm06uh9Wfzzn811S5U/Rh54NEdC9hq3Pp7aj5FiLufe8EDZSCBet/VWURv2KwRu5bPvRDaJuVd3
O1vRWxU1PKjqNFvsmiOjnzp3Qc484++U2sOSgQ3YOP5OOYwghpb5OS44+HsSnmX3pDArzlp+Ywcq
hS0aDqjeM92hLt/ZP9+T23K49uAS/Y8IkMmHFnDvqJFDDZEwJTOjT3hyLaRCnEH4DKMlhjlB0Nhi
01GtB35NuUo3vg/nPoKOVuNmNquN42c6kP5XqY1WmMK85nvGH7tj26MYHW/mIjSZeBuvahGWEp02
t212FSW0Lp6fXvGevltm3FhiwO+HDNOlCSNbWI9vt8sC8m59CzeHucG4wtV3BF5F3Y3a6cTm2PXm
Hoe9x2HvdQUeHMUfIKEtvXeM7Ta6mK+WuYFlM7cRiDwmIny+95EFgqFwavMPjkdvBq8MJY9NONp4
GGxgRSoZ5i6yCMGw321XK0pfeY6mtQz3hk3KO8ogJqNg9ZTQz7IZdl4FtwlDoweQhf0s/xzcow8U
9QfzvjGVA3LsNncbOEWnWJSzgUWux1D+TyNlwtsAYHKuuaEbVAq5Ea1CZU96KT/eQC0ORhMK/A6y
JM20iCQr520m+ZkkO1UI+7qZifKlLGF16LuaEpAd73yx1ncBXDzX91dhT6cKfjggKfjNQeWAkVTm
l0ZrohzqcciYI2CNPuO7Y5BsMD8+cAYHWcFzEyUmU9Z4l/9v7vuZ9ht/Xm9JTVcKutaU8D8hemxo
6AwvXY6FvHyZkIeJPTNJapjMzVshKmgf49N4EzodiH1LjBjPKBAHch7hFxGgXrVg++1+oS8GjsAL
GvFa3twf6TaIF08QriO8Kdk0ELW23G8uzzKHq6IWWugfgpDjmIzuZ2JluyYJGilKHBI2IsVEq2g5
uVgzhu1ycvyle4CwDlbYF0WJuws8YQjbSnEUvjoINah0uzNfJoXYKssUu1IBJKkwIEZNa8Z3eQ0A
VkN/wydBSwvNdx2QqNJH+Dkd1ge8kceXM7201kpkhfj/jyfrcHFrFpYogSvi7c+kiwu98WYcO25b
U17rGGaJwbVq8pxs68HzEtGsWAe3CWYBo0Jf8D4p1MdgFP8kF/8EyjH6CFYNMYB7t3ZE+yZPYj3P
x41DPLHuwlu+18qElppD6cr0EAMmn+AiB3bhOKQGPkhu7fiDZgaF9Rsby7gIGshJpa8G45/9caoZ
ZBrdlaKl/86KZSADPC0Kib9cLDnboHFFo1pRGpzaBsK+0otP354LHucJgcmSrebTgG1i62QbVA7o
/EjIaijs/LkoRTXp+G4m0eKlrgqWpZkiJeurbGaTgDNHItk2BiCqHbrxj1DzPmfCCskfC7u/sk2k
K0bqA+67eDverTV2NwQbzCE27VGcFlvr0Wv35fG+OdJAAULcA6CktXO/mM6wY+fqd3IN9dqtKrta
pV4AcvNDnI0gNWIR94J/xLe7t+hAW7LjwmUBzz5ocMQBrgREPN4JweTCPhYcBpsDnc3OLxoWlh6C
VlRG5YSoPTlhS4BAxIE5Tw6h+Gn0aRQu4aVMDQMdrvVMDJdxBW1TrdZ/clIwhkCCbox7kyzC7Jrn
aPkcCZafq2EYLyQFNJGpfHaszY32BL2Yqv8gPdAna0NTzeYeyhb5cdptOOdWKE1uFY3lVEcypKAj
6vrRKN2REYDut1VllKAQSv0YK4QGBpLUuEnxPqbx53NRvaCWnE+f4kcy8Bnbbr28BkON3ghDoOBJ
Ntzk7WKqWvmnbyKev3M2bjWNX86QRAKbq58sbHwhuxK2Y1XJdlYGhJJEBDseTnMOSTJz5tv7C+vB
Grnab7kfLGC6gO6jtUrsVsy5ysBJLs5GwliEPM3hTu1/RRLJdDbwdFB/1/EAXl1pEeBXyhaKk9lk
oXsYckUCyy0OEAyud6mCUHG3qOS15+bfSfpuBOOQql7Kd01XNAt3LoMbUf10qXk3XvF7uSY23mEH
PgnCxUQ0TN4oSotbgacjYJMW6jKOFIRSH9uYOLHOygPbiigX0w5qcjwcxObWnkjTBBACXBJl88NW
WDyxF4id8TJEV2KCRrGgTekob8so/KBmEF1roUnKMS2WCcuQehfVQ5rREDLdj+BdKLsCfIMie8vU
s+aAAx+MPUft99CRaqtdo0vkEquPXK5sqnFplrQr3Xstjqu4yaUPeaGTL2dEBnW7kT6zhwyOuKdn
sKjhomS2PGqq4VIOcdpa8hfg7odugQAToI2hqQlmtAm4DVtzTXHa4DPlUBbdMRFGcSQGupHQRHOt
eP3As1H82sZPXc+MMpg7ZYGK7l0t9c8wby2OpwZAHMJZlztWNA2C1CTTUfPqilpTwfPb2bJdz1UU
b7tpg6KURgpk5YdiQ+MiPCSvJ3Ls1Mt81MHn40kcSQaky7AkWKuhGnx2X66P48+toESl/O9tkW1e
8vIeKyf1WPzH3sdrMLVeGl6j4Bjb4oO/PIEv/nLaUAsfC0jbnZN4MBTHWGqRcOxcMOtycOl1f2aZ
mC2kPXsAFKjlzXExmMQ4QYFatL1VzYCH+SJJ+8Nwi5HD8lWik1GSvHZOQsYQkza3E4fCRxcHdkgS
5x4HK5JQaeXyVSE9FhJeAC1IXvx/2pguwHn4nwHYvqQ6YGf6noj4HJ7UL44TkOBsmmpESjRxlKD4
dAPBb+HSN8I/48VylJiwpCs4Inx4VEVhbnVQ3u0JPzYykV41N3EhHtBPNwd7OlBn5huHvExvyu4v
ySkbSqoIqQRgt7TJXHTghpCmTTS1ZI8IbHUqQsT3dtSIe6easGZTLjxZ0SGxXfHFl8SGgSO7NQUr
Bf/cbr3U5ZmiCO3M2WOm3TZUZa0CDhcOEjbiz9IYFYFJB6rdxnyW067NSGs8Zpa2uBFRN6XYelCD
DKUATC6uIHpbVutzuz/++3zaobPqDHA7pilW/0bUeE1QVIy2Tu+fF8S/OX2rpMq+aA59uI1mQg1a
ZZ74JlnrTptB/4XW/vhUAPETlLkfK2YBCSkF0dvueB9Sl5X7Gj3ByYmCE69/vCtp55sfOh8dRiTD
PXD5aEiZBm7KGcYmC/YNfntiyo3HOEmen5V9RPT3+2gmbMefz5b7pmloCZE6bbNnGBrhwJgkOI44
4yu9xjm2CmFWOMhzV0/1F+cPjV5oPtSsTSPi3AU68HmzllDjSs9/Ow3axHuCcSlAXR4qfLKFudz7
KJdWzQMr+rQ2SdqEzbWGu69btuFKc1sxPT6EBF7m1RBEdjrKpxcb7rzQEoxwAYQll+iMHdDdN+on
AJNs4pz+yQDA8O271ayj7REPoaFonx2cJEnuAeZHwiOIdqMP8UUGVFUX1wFyFSE3W8v2g+nHQcLJ
lkJzHguSHWXocw6xDsJQ3WfLfgGQ1RJydvXr4ehuGUAXVkwQkp4RxlDB/M2XxYjDe/5cOOEqeImW
hP4aOKulYon7l42v/y1qqDmZXs9dwfncphHookRt0kcrumhrAgXlhU80Tq7/s690coMXTueLdJUq
+vUwEjV8zqWDfaQyXNyRy23H5xwap9GfJMcuyOU+MZXcEVu+0MeIzjJqAn28hw/sJx4hrvKuGRD9
cKn1lFaUvFbZh6oiEEQyqe+FXeHj3D8BRO9iZtA7PkKcD0LfbdfuShd7J6xZC7KTO0lf5Dse5Epc
SD+6Y4UHkYuXrCxkOWu8G8gDkYhLu4u1COy4+tfqR1LlyFZZc6pxkhOHvLmFIRWXCnpBUF6Wf9Rh
4RmjmT+6N1ZIHGTtY2a26KprwKvKxCnWTG8GHcbtQKnwNKd/xLqPCB7TenS4UFZtMg8jejmFyZtL
AkXfz3PBfcfGbtyPHz6tGo2cuB7sOhojfEHiidOhpDjSZ1hlkO824/8AI/1KNZSmz+30h56AVFJy
gIvvNx4Ftu8Nd6l8qhhuXp1XY6yRIjrK3DsR3URwn7kl/t3d9O7c0YPMGIg/fIFccvF71y2mlko5
AbIo6Tbu0dmV2cUL9FRZVEtxredY2bSdActPclAcCDwXWOX9WjoW2NlyBLisPql8Wj5/6CO2XcNi
unZ2sXj0JiKOuOpXKCKtrvUpcKD7t8zdiyaOnX2KOvlBR6K+0pS8MzGxYpzaymRd0Yinp0opxijP
u8cpP9YCWfiSWXTu7KGf7jBneaunjQCZUbtEuWfBcfePdwKDN6OJGYmeAyCPkuKG8E39jBjlzGpK
qT1C/i79bDojadZ0e1sUu4Du9MolOYS7Ig1SvSJXXh+VRpXaBz1gkN97FKQDs3MuVVb/g/8+Q2hg
09yEDsjUQOWz0TPROz9llQXnFt2UodfA8rgBc5xxS8EAVn9Ujv0v1dZYJ1A3hkI7mp0VgCiMByr0
Dln87bZw8aJafDXzeJcbGAJE6RGICrbo8LJAZpRTyFMPgykfN9tkTqwDBnnCDOpltpYsgC6vL6s9
8ga6c4mAd2GxJKsrNLGrHegHKBiiurqNXddOGgitibkprdXSypOtrV7n6zVsDyknGyl5U1bWSAKR
Ye9kMX1mxyZHVNb3/iTRjpXGke8WOushXY6LmlHVOPbI5yEpcBoUQgOpc9Vc75C9oDDyRXOj8JaG
La3Jh9fZeTRH48Me6+xNWKkp7xXM/9GmDO1cuuzwEtTQJsruQrbcUwjvsFmtfoe8x1dCG67aVFtT
WaOlJ6gUIzO5sB1VgtkNZad07chL8sk3I12Z6elneGPmGONjEIZR8+8TDFngjwNnl935zr7xMI9R
JRt7+3tCJF3k99A5rKdmTmJQIQVqU8pM2hYSt4ptSUi2YHCZH7E+0t/8w/2O8VEP/T0XEX1JXu+p
rhrcLnYuuUfrAuXGSLt4RHIgiQfgfOT9kfgWHM3tEYbdAzD4bnoUk6VOzKPT5jvbyVQo1U1MueqJ
ul2ThR7W8W6flh8Nv2jfafprrU1gqzJRT6Eh8omTJq2Po+Ikr2sFKugqabWf3WT1MoRDy1I9VKoe
Pl2RjSYIm582F/xBOJfGUlnPIgbe8B38WD10OHSxvK5nQguPvJbkt4/W/tnATgTrFogIzomcebVu
Uil84Hygf/bJmL73j89Uvzn+Z08cjfvwE9ABhFKpqn02QGosmpnI9D31Gs/plNDBKY/WhEBaCos5
AQUu+GTCrGSx22MDyMqTR90o1m/er+ii33Rf0t5Mf7FoPEOVNAyCVBQF5siwebwZZMFR6CrMrrZl
0U6NdLUGVe03TzOO0ir1hDJgD7qR2CRmcX/AKFa8POX4UO0+GjvyxRsDbk16t//lqWFcMVE0KdAt
OS8ppG/TjvV/V+8Hl61CGaCP8gTlgoeiquStEtNp8j379IJgu61kPAhi65UvmcPIVveWL6ReqJmZ
qTs3f2r1Sh51uEc7PpySQryZvTtbJCfInpJ2TuI3epVRHQIo20/tIRJRF3eY3ohqQdEKf8uf+3fF
n1hM1cJQIKQEbtQEcXX/mzE05RgcHR4pGprDVW82XZk6u472IR3JNEVV+bWG7TJL/xzeW/4+JByd
/Ewtz9hzq/8qBrJ5Tidn5QhDYvGuPC2Ppz3ljQx2UeiMpcYDEJrJmRQBl5EFsQH+Us36GFhkrbpm
7N7/Y8+PXMqUsSDnKig7e3kpQaES2DkBkN4rBVvD+HP7bxGCenlkUaPjtESFIAFxH4EJSk1214ZM
fH90neW+YwjG06u0zcHLUV8Le//HdDemG95RS0UvGT/dzmA/upD8PeNxJMvHHz917Dd+9FupYmhc
B1y6q5MGc+3sZklZ3acvboZe/7N/5B1CZOBjZfQjBgmA8TeVD5ZZM7xDeacMC1sIUOmguDxe6Ow2
sWGMJ1D6UaD0s1gqu1OWXepuvMIr1mDArH+mGC2HNvxcwN2Xmc+wvml43axE6DfsESOke4ksrzOG
/2mnFFBw6t0PBpFktNXBAaa8Otn65i3l2eGr4G1qy1Ynjiu6n8Gmcfa+nsnEw/n8E/VrVLvIfLIT
B8nzsUDX2O0OwbUBieULscfniyXS94h0m+0dN/DGXAUXGDak6AGGAj5Q4GZPJoZfzVUbh4qZS8Il
nJ2Lmn45EI7NwkSz7w3So3ZSxMZe6BJZ8ppx//qytjzWeEwqvby270/FTReO+d6y2x46Hw67M9jT
Xer3ITVjWAsxI0V83DZWnALvrOyEWypLWCh7pKedj9m9RZrSBJgadEo22NYSUoSf+8no8oWq5TmU
UfSTWmARAUk/f9OoRHG9Vb22y1eDOJAri8dw+BFA/QCOGCF+gq0wUZ4RJ1EuDmt/ZkWD+S4uP/za
Cr8UhdLusLslRiHEaYY3akx8fcYXcR+nMlpIJjLBmWmEtz5nTSjWem9VbCCa/Ki4dNQ7RHpjYC9X
SlYse5HivrC/mVl4brOGBLyBjcsblZxbskFQylyqMtpnRBCJdZycl8nx9QIjwYdLxAKutv758ffH
e7QsuWLH8fuUwoMSqjtqVrRb+RLcAMAonoYYf8yEsbDTMgRhHY9H5Kdv7rACxEPriL2zGajuzSQB
ubSTxDROtAFlTzRw8wRiTrRq5dzrrozFwgl0rPpR2Zl1SJHIP1FLdzrI69oFt6SInAucv2hoP+qF
kLehrz6qcHSqg23lhDXJUm2SGKLc1jGe7jvoY7b6Y4qzpu0ssVEz2+EUrQPqTEHW+f5ZLqtJ3DYK
ZX/C96NylLFsxKjEdPjV/MadpevqdIA6HNSGuNrGReNKOp4xsZlZVjW0yoJCLOIO5u43vAeFYkO0
bmg5n9mC2q9C7CLE3DlymZLItc0Ys3OyTeyBHLKVqjKU0rQrMX3vuMvDxPsmvKeSvZKcGfCMnZe/
kXH+bxCH7o+zc+38DqtDem2IRHYsdV0RQLtnF1/9dU9nr2DogQS7us7nITnbPQPj4R6iZePpngwE
FUIpaZci3uBjedM3TdJ9HSsYP5klih0kIxNoZ5YS/8hXTbpC+Zn75KIJD/+IahqkoUGUdz9VQotw
+jdZjdNtGgeGB/nLnKPGR4hF1c1xtuDobrxMjszXVujfJ97LzBZabgE/66c7WVUBI0B9FPzBTW+2
okt0wpT/alIL4VafQxPeYpS5SVCGvlnB0DB4Zs5GB8slZK1xCNIg03kLxrRRbJlQ50oXwElOK+mE
QjjfrGUv8NYcQAWBI5l0cjLa5kXFyji7CfyRpnHgLcimHpPAHGI677n+4Z1GUa0wNjUpJO2SpHzj
EDEY14q+4tPRFLnzjBX5MJUO06GG6aD8ILFAKoOykWr6IefskpZvd1kXRVijxCkJS5p2U4JMaizn
WM6Vzi7F2WJrpXobXlghGChqP8ZQmI9JJ5nGsZHlM+/SvvxaxX7jd815VQi00EA35+0d+V1JEifj
fmz9zzpmE/9P+4e2tsO6ohhYyACvQlJ3uPCna60RQYGSkffxjtEzpXTBElLSssbgzY98gzjKR87t
ETeyOoigqIKc+yFuVxXqx9ME0rumPYscObw9L/xOCHPJF+NVwydz83tEHlzxikBCLjX4RdCirmkG
s6jQvGK5jk39h/rl2krVPKSR1qJ+3TL4QK/CIF0Xczh4jBRsvHqqhzpGGbcJbXrHg8kd+Mih8pbk
1c6bs9Jg5ZFg+gCNbp157Z4TDYjBMJoF/Vy/0DZ0FVWwg4mA0eWgHZqy+VorffDOEx4840kPMmZG
0Guhe3mpUgxGYH/g7pYxvpFVaeZd/TJbZyzznX5fzZ0/R15t43fZM3skZr62KiU5MTeUdNbgQJzX
Yf+IUFzGN2NXwFJ+zbh2AJhe7VU3NIvk+haNRXBkxIPXCxDgUvdMvbq5w+w/EBgBmPw7zNYWdmtF
ECdfH5ncOyJdUxchk3YQkUOReMCLLePx4RfzfzrfKufKsv0CwzqHt4CKW3oi8VYeVzSSK7WC+vSx
7NZLdeWgFwX4v3lnQeuERMQRaUmmZqtoOo4C2s92WRwvhKPAiQ/SwGnHGgIhdgdkQbdyQjBLts8Z
iW0H1h5WCkkebrziRsl6IHapr5mqNErlqx7FrOti35C1By0E9HGmbvPU6/UvaTxSI6EGusT2jU48
2EHpi7dKJjHBI7l1rOPoi1uRdUs49BA2eRHWS6C9zU/c/mQuuFRDcP5kNB6F3l6nLF5cUhgKEI0J
zsLLuWCbm3zDlELSW0HacV4gH29jzjGfRawA+UbcsGp3Q4Bjfx/HXSWhk4KmerNuwwFYErE70QNZ
JkQ9TbxIqq3EpkYcww0hpynGtG+TQLb4mGFh48TpheVaohbcsmxF8Ze8ED85y64G+wL4/T9kmAJ8
GFkJ2n8Fa0wywdJfPO4xd8YniqqXDqWmaeL3i5663EBPnHSjpH7wGWG++ArOBGbaAv7/tgS2moJ/
hoqx5IVyz4e6u4AgFqGTz6fGnTnPXA0WZPNEmI5IECa3jxH72wyB5/wr2FjxAsnEBe/x61arbWk7
492zn9DS0ss5SbVaa1VXAEOm4Dj2usTFceUkepVPWrVixk1cpDDZoyU0yOY/xQ6rYw8Ddqe+GOY3
xjTy+FoVCY6fEAWWPiLIMqE/6s02NpuyXOeMRzz8b6kl9QcyAN/AxPOx0b/j2TpdycZydKt9Pxc+
8l5cSv/sC2oVG3O9mUrV43WtbFSbjeX+T6bJcle3zxh9ymteW5L1O+9lz+ILNrMqamT1bJ3GXpT6
2ji8zk14Sj1RVfsT5339eA7cCkGG3OMEY14I2+L1gR/DGbZeD5NoOe2RcJjjT45cmhBptu4lOQa0
QdKQ1d7HFry8ZRs5Ic0jyp23q/m8DteDqBk0KZc4I+F6kDnpnr3kkiwutgFbH7jO+MCe+x7G9FFv
T7292dsPJIOYUMz32kJlwPVSAGjO2m98Rn7rZ6kuGF6vuOzRLpncqetOE4nj7Af7H89zhxV3uT5u
W92rx4lsyGQAO51Ro3cpoQNntOZ1/e3lhrOKDkDe24G9a748C7y85zcgUNHkpiVLOxJG1rnrIjlJ
FdLaVVH+09l4q0Rp15v8u3fHQeVVFsdovQM2+3nUaJtT9QUKwgcF8S6febToyA9/FKk/oCOf+Nha
uCHywAg9or4Ii/8/NTjqQ2bdi3ehX/gLZFmS4sANgWl8uctqQXeE8jKI1n7VJCQ242mOVLj4Vjrh
gm/WWUdG5CZMZS3Pm8EfSWfNp+NouSyWsgHZaDtgFDMzAx6qUNEq/E/fD+f/MK7LRL/z7BhPxL5/
kkcmHf8CVhBZxcCeK35+m0R0gDP5nBKtXzk2XpuGYj7rkXyloQARwCjrY/0dbkaXD9YtaZYCOP34
HCWG32KZeyVASIFwGi2OSErFzTak9n1t1IrsEtR+QaUAK4XOEZtJKK0r3RFW+doLABwOmW4uwijV
AF18EkfweDTy3GOhKC8BNcLXvF9zDLeczrNAWc/Tehdhjkhlkh5O/9PhlntdSPKW7xdHmO5iwDZL
D4RHO5IcQ5lTLk5icPBSRRR2kwUAv2OpceOwNZ9MR09C4RZswUOjw17is+1dKx5EnzFI6b/GIUBH
nFX0Jfa57dNRls7Tsxi3V/FV94g0eM145jUxwvpM3j1MaGURDMudfCPZUP43+wZrRzFmCZsJkR0v
GO+nwpz+jBpzQEoCqDS+9bTbQ1nQVvKDkcaaz+x28BAZ3dBzkrcbafnyFGDGMrvsslE/pjUu3YFk
fzypEfI22hgvB46/erQIBv89brUo2KYeBIgGhXuaBAA9EPXya0MZHaCBNlIXacdaYmovlDuutLkx
yPOiTt0ssf63mwqm2+utPlyA4Jtw6dq4dQ5qCJVALt7tLY3BtfTfqJXulc6FstCq/YstWk26kxxJ
zL2yjY/OCRLhcb8q7FCBQ1ObId6mDQqisa4YWDC1fBD3tZ6cXwmuo9BNNbUJCSTSSQC5rsN+ERRA
mzNXT5TwExhG+p5T/r2BQM7RwKCbHF9mfLbrVBg6aWdLoqRJj0TQQaPHTqo5LOj1RFnBXzgWMr1X
uBTc3jDmp74eyvBCogSS4QuJNhDt1t5jF72mprKM0goZZHUmkMuxe8JjmcNw9m8L0zpWIgTuR1ED
ATG+ngLi7kbz+O2sHTjuhIxaaVkYfxurKlHnE/bFw0DRhlcnewTwviMUEGm5ezluHzVg5wBD4SjY
PaTih9Dyb+WU+GwAS6y2l95gnr3e/Dlm7aU2MEPQP5X0d0l8beptJGpkseBWMqHeCMxrIMTvyXkz
MWpnkZfWAN3xmgcUrR4oxIRnLCf8Elam7f/acl/reWfTFlacs0OumZF+xwVl9XmzslcHb+Y8zs9S
0Kp/EVEmDFnm52QFdZtwd8TrtXRQ6QzrufFC1kAL4+gK9CZZYWitSKzGVer7jQHQjOip5zLg2859
d2Q6s78sa9xvMHHx+eZ6PB9KiCQ8mKzjdS299fU5il2MsRvrriFBGyukjUPJqnLzvRX0+IiH6RbC
uheaB0ktzvjURDa6A1WyclSznJcSMaOe6BMxSY1DQAVMLAfgmbKtC+wmhPU1eIawGX2ZURICjTtT
kjbeJRsZhulHt1r28BzmqxgzKV53nIPwnb25Ypm9Vax2X98s//+fTYTzmSWzZjzQg+VNA72PggpJ
0YpQesllkU1cbUNR2ubQrKnxaaJyGCrPydmtlI2HR84KhMdZROnp1byoI7WMsRXktPintFx4QSMz
seV7FEAevSAM/cBJVyI14r7KuJkHZcpPDac6E5G4+ot7kNhO9FmAeP+j13pfaVHNYLMRSuep3crm
BD+93gQLz2sPy6Eu6D7InsA55BW2nmg/kqdh0Cxj7SPFyQW9govXVlOYOvKvhPGu3fx9RtYkCkdG
C9qSf+IzLwPhgaTj0NBKFwCnSLdmgx2FJOBUHSOgLg3cr/BWQxQXpCvzX1qoIJ62klJCD+YXD1Sg
UZxLR2hD8iacd594QjWtDjcR1LFnNz6QImlPqxVIt1I8F092+4vGfYXVhmvP8ACrvE5/5oFYgiKL
2agDLvaWpy8jBwcMKOUVmmXC5mdl8AHlLurd3FMMSLU03K0ci5GdmFuIUTQe86q+ErapzF5x9Loe
wMr6RuBJyelN8thfvwrQW1P+ElSmL57XgqsDH5crLw2Qr4HEKwEh5PmvsejeYxKpUd+5h/aBcvtN
whr12yo/qywSZa/oVvAmc8GvIQXrKglklkVAt9PYeGNuZ775DbckWGl6R1rmCJxtoOA8GA5qvjay
bhZ/Szo1DG8ed5kUBDIhJ1bP0XM+rNbs2nBoW5kaT1c8VHiLEt/0SpzyNxO5jBI+FUVORXxAyT79
GYyHrLLDEznZ4cPrjchQn4X3QINTxeK2A+qy8nIN23MG+Xa9PCYfujB9tXCY9EusGb/jgiPiz/dg
qMol6VShhu+mSWhob7hUZHiFbgEA1EwMvtJlXfQLoS0RuGRjlydth36Hq6ebKWsDEiFOP/mrso00
2/lk4mx1E4wa9/lAZgKIKI+HoChfvVTZyrH7QZfrcW5xK+lK/u26bsvrKodvoJfIodR8JBVTQStl
Nr2zvd/ibNa/zjeHywm6t9mZHYX45TD3j3UE1V4BmU8QbPzYlbcO7jcTbiBDBHvf+BxzBrwF6HGd
VOqJDtSXcl62TUw3IUZMMP8Un6IS+WHpRASX9H/H/U7yPb46sYO0JCR8JR4oBogt4qduH3zszn18
gui+Ff8RzkzrTK7GhB2oXAhpxRmfu+jqDztzpc4VZqorTfxI8dSSUr7g0TrS2GUXV8WHBVu4nMeM
TrYLDkvV3pBzOVht3Ua9uGP7myhcA3dwuXVaTKONH4s/2/bHr2p4ZNO+b5rrYNmwllP69lbQccqv
8EZDwnJubHRp9XhwBUK9tcUzADu/zb08wlTuFF0IWgVqd9davMXTfrqN12rTjcDY9TO0gqi0QWy7
Pvakgf2kAWTJmwzTgTzh6D3zC36opIJWTU2G3YnjMMNidn5GVJyTaNM2g0yO6MK4ICn+gTa8o4K1
b4qzt/psPGQAye6KZNgjxs3ryO/F5ngYzR4uZ6kgNSWgx4Oo/hnoRWXl4j8VZSDk6App0ZfQoxOT
hHuOd+74s5VCZaTRMdF4qDOQfkzVp30tncHAmVApxz1/gon0ndl3OHnj5mA5qbLGOeVbbyMiCPkX
Wz7OT9mRf/cH5W8EeWrxW6DjChY3no8Zb3eXY2sXFVHt5yTFqXgtAQjaJoE0W6SnYBM3U9olF8sD
vrXhWDLU5AC99Q52RdGJ9AIAt7zHGWhkboHbRIDXDbthGQyI4zVNLiABEB0LuiPLlwT0NL9ej8R8
33JJ5zv2yBnYwiiKf2PuN69EbXcvOfAETgwJ88uYigTUgqEWDHx3Y8R22QLP48f0aPs4s+WJNGVy
NuvALu86WB8S0Jwn8iV+fpJb+rWm1nTODaJPbj1Qieb3BS7SKF1ZhhCZhicpAPfnfxhO+WKDCGNG
4+JfW4LoarnvOd7X42mrAZJlbVY7nye+PY4lSIoNc4H+g0Uz8NtcPfhLSbMGaTsG7zsoy60lNnQe
59wXeuHUbggC47pH7qEghP9JrzcWTBYPJGBOVhhNwcgzWLgbVtDDzT2v5Sos5u8N5XRsBQIG1sY2
0mx/HKL4AVrEtSh+cuMxQUEDmm039Vh3KemZEgwQqMtc1028BEY9sh4ktLOGz+oQidmjEFuEYDSA
Unab4tjiMtseamq4sJOdiJyRFtAkPakhqvb356ZsD117dF3OsXTiUwXlXer+VMb8BXZc84fVgXid
Arc/95FvvGTYoSPRab7UJXffDzYniiABe20mQegLEjrDhZmZlEwlC/iQHyRm/4WQ+IktCv9KuzNe
ORUDfMtbPQ6YBcPX4mqYXPkzFzrG8DERiG2A8yTBaUmGFnqgNzK8MYyyLeWb0LpJsdpbIsUe/0+G
i/HdElrs6Ql2i5260mAO27PJ8H7nqNX/+MaWiGKwhOZLvlYj9D2SbhC3QhB3i8Cb3VsyzHfy2UEI
e3qpz6x+PY/4J8SQrgpVCwW5RNzUCjc1GlmIJwaaTTnimoXuIOXmqlELyfdtmGzko3fdfoqipH7X
QrbXNSLMhUmz5MhEMJFTuNQu1RUIXm/Fu5G1YFwcC7Z5eKKElzb3lB0owDRsfhNqhIdjG8YeuS9K
aRVrRjnMZo9X++o8LBz3LyYoQw2mTiqc8MbMLdqKQ7dLfpGJEHRGT8klQtqP6E7Ac55EcvtdoUpr
2uW5FVZ6up1ZVY1BgFndD/6vP9vG4EK6x25wd/+2kKKTGHmsord2GRkVcQbYKEx2tTcbe027MbJP
r8L0LKeZeKwrBYbs+OoCZ5KP5wokh8KKROZbCaORncIUd7NM5EXE6/+dnOhAIF8htrgubE/9tPeo
eXTLGwHKMv/RzwzZHC864Qplu2YaUjcJYwo7sWnoC76n12XZO/y3ACSIDJNt+jMmoL7TdQPkyBIE
Nyv1c9Ku4MxwyEa9z0pDPdJu5NEX00FNPDnjVHoZHdH+0wmzrMho2Kr1A25KrKnacWiQrFyqWfVc
uhCmPDHiN2MO7gL+Fdlo+aPopR6c0WM+by+hS8tR3dqkEcxlOSwD9f9flGvakFAG8P4RWJsqGL4h
77kTHA0YQp4ez93eZcSFrP4Yqz4snSlXwb7OvucPB7YgeNnBiCnC7X5PzHxhP1tN2Fx+GFOuxTFO
mr4AOsEnMgkHOIViPen7pDWaT/jCa1q4eQbhIOeu1FDSt6KhiuxYAIwlVFXkbNfLJSZcCSgxqyNQ
WondH28m/YHg1LV9+MAIr2v2jmgWwTwXcBBOH6fvkp2K0uysBbiHci10ysng3l967AvJGlv5YYjG
Ug5NoHlUaAoc6p9aspBiAnQ7N2CiEsW4H+oR0OLq0LP+K372iNRRe+TJUjbMYLYnA+puEMiROCAY
N7qKqdTSG4nR4r9Yd6zN7ETL8lMlwFGTDQ+wLhDnIRRrs3B7ElDSrUR16OEniiIxpO8T4ngJZiHE
BW+8OEojzVpOUoj9yunXIrtXlmMHCI5RA1AGFas2ao0Ehm5cT17w4RnRZ6Hc560f6S4Rw/+HHJ9a
P/HskRWY5tWeQ0TLa4sS6muML3UISEg5qLkPgoOOBH4Gja9btHv6jOWVt5r5gMRk/l5w2HyeUV0h
jjL3GH0cCNAuxjv2s66m5mm3RhMyImlVoa4p8ypNxJf93ILcKHdCE4EYysLBjO5jnaNppj73yNSI
7WqyeMVL1O5uykHO6mGnYGGOahG6z1Bd/kf946UnOhi2nmmWFSBdWBy8sAaP2odlTqnFLVrHWk6V
BuRS4AM3adcrbFBx8s6Gka/hi5IXaepDKxma/RRu1ugVr1XCO9chjFGaheyacsbxRRXxOdKuq9Q8
4CF6BSORWx9UztzVffVL8qq78vx3+ZBw4QGfSaXCHVeeADtllHhqoMfm84zcmM0L9OiVPCcoJ2uG
9ENmW9bpuX87mUsaqnwVj5kG/Hx2Zy+6cC4q4WHev3gkZbhiB4Jqu/fNCvrS/7RIwl7CBh1/oVdz
qDOaQR8rpLp5eDoHPmGn6jYo4TlguupWNJFU1aYpTSUPBn5fqhY8GW8rtnCmPCWvILojtLs0qtPs
llyF1QoMRFdguGYl2ez3TRhEVrTmngit+14aBi3NoWJdFtAj/2hdGY2zkQ7rSKo13wldKP6mr+lN
DCQ8WuSU3Dee+SVbJhCEMLHLtb2uUjwHRmtXc4vAjQXGzF2cTsYLRLaxATK8fYcpP15IlF/qixqE
PIJlSpXOIbfnBgh0ErpTw6lGEbVrGH4rePgQkziiNLHuAsfcTdGbp4KzXosAJbSul4t+SA1mHmPq
N6MuiX/jr2JdQt7vEwOnHHPIw4diIwxhFwwcGOFHfC54nD9jf7hDYpm33Gj/PG7rt225LMRXcTpn
owj0U/U356URHH4chyP0OoEnBHHMOu3xvB8Cd25xO8oml8SWwdvfNdU4kSbwopAl0KMSM1J84bro
fya4ONCcrw7g2x4eFa1y91wBKTebwuEakK2juLDxhKwHRCrpoRylpzXplHZqPVld9V+3cxsh1U3S
701u/kvLrC8T3Q0mN34tF7R5m3+QiRvvrg1e1ncTR/J1Hg79xVJSODUIgpQYxzY19D8LlB6pejfv
rlGOsB/7ms31wwB840WM6k/l98l4ry6jB0BZczix/ZpItMFCcJlTnQkHTJ0LSjqpp8BjuZJaiTrQ
o7w/dBdAFSVfXCDW3eFOHHDa8xaNpASXADAPMkn0yZNRvl5XFQLWCF2vghkWQlJLUnuIzQ7l8xgF
UOVdGkRxIu2loazRz8o+ZNE5KzRcb40kBJLkl7YKrUO5m811wA1nprbM/MNeaYZSDoKXBxQ/ez66
GAyb4q+rNPpxjhiT9VrfGJRhN8b6+NPIe2jPlC6zMzk7wBIR40kKCwkvhuErUes1pVReyCtMvRFV
J07CvyQYdy3w3ZXyKVA36Ji6LP27gHqeTrCokSV1eXhOcKo7CrscLMzpnZbZ6pL06J/k3+VwaNX+
Yq0L6kXitZZlmmN6HAYxmynobG4VtaXbYvqBkkL0lsOcRMxse1CdKlra3k1OzLNxDt+wYhMdZrms
wqzqLW/GukFcmToeg8wItohHYnuEcctkhQ4MiV+mUHtuaLb1y7290p8ruGtaqnhODVJqX4zIVO6I
GSvW0EpFK4jBwE4ueNYqT+emtKw4+U+k+O3vIFwA3ceII2bSJIpJcTHz0deXyopVLWSj7L9CYElQ
ioAGddvO0/53DgpzEMeTid+/o0pS1nH+kbZsKzkCkELFgZfKD2lmnPeqUTneH+0dlx0x+oGxzQhw
tZlQIpEY/AAhgB0A022MGDIs8wGIcGVgRsD03kJRXjDmJMd63EinGX6odtyNVxCYWmaV3Uvbj6Ao
u7kScz5R+nrZ+7rSzvj2Ywc1Wl9WNY1MDJk4bbq1u7sfocMGD0Lzw48dk14LQhQe915BLkG25SIM
hJFNYO4zzrAJQ+Kqsq7Zta7slhVbRgmBdXLK3V3jQLznjMZPRwiVCw5iJ+gWAEHEzmKys9YL2CAH
U4eBSPHCCL6JaByfKzw91Km0/ie12ZIexOH0AT41q+T+KGvjjhqraVWjxmwC2jGS2KrqSwpTTT5+
mlChRzbhycuu6K4wLhJZRkWr0PCgSyMJm+7fM8krG7YfXrpwzpWu+GqTQuxcyzTq89fPqqoq6erS
fZBiKWXo7YqW2maAXlEFKSeu1HtVjpZx4PMTHlMhJ3jl2eaQMuBWz3rvwgiTkYlmWVE5wWvQ+BNa
7DiQJhulH/MHkE3eqf/axJQ2ccxJnmg8wgm1FfV4IgATT9BwpUfNTIUDt66Er5nDhQFRmtYjfwO9
YI+34m/itt8V5eL+GCfQye7NUwwphfUauApIneVHzHWKx7flfHFZwhBky++0jFKyuDCZWccoTC3Z
7f+tv6IthoGAPjOsczIFerFaw59PBTUhyq4fJrjl4KajUfDmyXe1643spu+evK/qA44qP2u6LdxX
I7D6y2PgfmXSHjhbQ4jLniBfJowCL1rmTbbJFciWfDBo+Vm8Fz2GOZ1ZZmRY0chEOLapZVnPFrCC
Yma2zJ5Owv6PWyA6O/yve1B+PmqEzj79sPrkvFlcwKlMXgp6M0XrDjn3x8hAAGJQZwkrxJOc2MHy
U/gbquyQi98Youc4kuoU1eeJCUUE7X+6XaAb86Jzvcdg1miDi65v2OG8Hum1ArRLsKl2GSLD+jYi
wQEr+NcwjXSmE2oHTfqDbDvcp1vJywFj8YO2adGgNlUWIHkPJm65U0J9QJ6wajFoQ0AwQCQUJmML
T72cn6HbnPtj3coQxhuCWUJKsaxOTu49fbeiISbadRtqrAPI6S1mJkrgjNetA8QXv+uevJOH3cUD
JQe9m85Jffu+VjwPD6GXFlAl2NC2O6YS718yqIALiNgy0ulhFrfHRmWL6CemHt+CV70mKEHgofK9
L9OeDGXXN3KqpLehHOCoLhyB8FPEJ1BpMJgBk5TqdSl9VnHPtn2GgAL7wBQ+RZwHDGBNWWzy1+Sj
B+v/u9zLgVoEMVaW8Y6PFCCMyFiWQzm6GFCNTH7EdeZz+xPmLRU4J4ibhUnjvhnVFIB9fNI/eOde
EjrhL1NTnVjh3KdUozvdu4qTxVp8zlk09QZA4TienyzWLvMX633jCW86t1ovBaJfaoQ/ThjGmwv8
UkS9Q0Z8sPYZed34mt7RToSR9pMR0bxxxhvOMav7hkPAieVBIhmgPls6gpLaZtd2VC+OhUvF3A+F
t0bWm2EM0Mad3izmVSg4gJZKHBzsQe5gYgAakXm9H0dkIb0d5z+45WLBgyPRXqxq+ttkRqMuulT8
ZS7Ona570oZHkHbSR1aOKddzUIXI3v1c0yA8AyvmDN3s4IQ6W82E1cGYiRLqyp/67H5ptPET1k3w
g9xg6+ZTEHuRT58At0W13r2P3UrcTiKfwLcpoqfvP12CmeRDv06v37+oQfhbnFIJCe4RbL6i1Kez
aVMYeTL3GK+PMN59fpNQMRhY4sprQeVjf2UjrYodLed5u+Yi6qINKZZREUaXEF/WNd8gZ/neTg+S
vU7hHBoz3uw/Oo/TrCVGsGT+GlU6m4GZOUdIROXnDfhvGty74A9PhUpV3Ot83To9XGMBiSRjw52W
mkpicqafqyLkP97RVPdOwdr1BH64lDx+zcP/TuWwFYritoNWZX6KY0Az6rzzzVpTE9O1odS1qy1P
Dsiy3G5UWZESEbccg3UJmFxBtwxAkFnzu66mo//lRR+X4s82HaKvljlDdYUl6Dzn608pSQbn7HSP
lGCAhI5xDFw7EEcAUztssC0F2fPHAodhGygnzxuiCvxNrs4Hr4G2hQKNjDUsB/I//wdNLgxwzxXU
CsoU+p6uYjn6/IRREslLAC+hL9dxohKDPT3VcJHXSY+qmCC1Rm3vNM9ChrTDWGYXoa4Opq1+QEjj
FR74DkZslpYPzN2ecsgQxIUkOr2o39EENOBfyooS7r10ukcHCW8KEA5hl8xaWR+xQYdBeIZLdblM
nGGPBd6HnzjiGxMulAZn1g9JgGqbQPPfRYjovS/wuRuMMp38Z15/rjUGKpuuOXvKvAaZyDWYG31W
IQSg1DgOGS6ZoVoIY04svO2MHxKCNeqtyiED4npb38yclssMVOOIKBJosvE4uDvqRtgRbFV0Jr4Y
N1IJmiu2Up+CKUa7Urx273LgncL2cTUixql7nAawg4EIPorKC/j6mREGuvl9PGd8b7jbHr3icqyX
1lPwHcnu7wc07lKRH2VXpPsagzRlVFveggEeHx616neG6p7VO5Y3Q/DJcd+L3/SQirUat5mDkM5k
IqbRVK8wVeYeOv2m91CifPxrrwFy0KMiFWMt/vGAZZH63VRdaFTvHqSDZjivSNwejHggX/rlsGVr
sTR9+1WouWRkrscTY+yUGCpipaTdZw0v7gl6EIx3pjCAvh30309dHG/k9870S2Me5jxLdm7kHDEV
u8AOYxtmhm3lB/6PEqN/Q0Kiriw+kjp6TiJBlvNoRPmn4YMiqQN/7I3Z3CWAfyobZA6BGeCp/YPA
gvqgjqUr5yKrXPl5ikCozrn9pL4p8NHKdmXsoUPQM3808LXF607APyrAkSTRnrxWrEhAOiY0tLhM
LlhlVtdQtrnQF0yPKh15ygYXEqJTs8f09YQ8m1mp4FvDZVirVpiQhrxJLwlk4t7GjqjClAZ48skE
4QzHM1RR+96D+xvPUKFdQUK7vOuwOjwPGl6alO+eKKk0ZeyvJam79MdODw8k0YAb/E6PCq6IGqLW
78/ez1alZklcEOT3bzb/EkwSnX1baGiMHK+cDFXHwM8MWONkoOqZB7l6c8GJTB6b6r1C3uJtYd+a
yadUNAFAeijAOAlg1Pz4DZWVH1+kbSWgl3ozZyiHXzabkgvxPXJy9k68rxTlNvRyQ57UBh7weVvr
PE2+KSfxwAer6xT8F39xCo5AwJg+ivhnPmYfrXDKSa7kcwkigX4TVCOCQ06TQ5Pw15Evv+t57wH8
4SLQ0U9RcrYJZKGGJZZS2b2FV0XfQAO4VUSJjXKUOVjHFtqP1Qx7ZyKwQH5F/ibDjEv/NSIui8AA
qnqupS9EDzCaGStseiwN74soEAdKklE3czdLL4EcpXMse+kDg8tp1OF+Ym87tfIdaqiqNdzSxsGa
eiUSrgYVDJksQVJ/DF/ER1qXxup0AcxCGynBlWKk43K1lY9Pf9PwRXX4EYxzBVXizi48CjHrJwd4
j4bOBaR6DmcSuZyprbIbitys5N2+NeBv5gdw+ofXUfWFw9aWhx1mcM+bg7VC7+tUuf8GH5LR9jzU
/55zTttmddOZW1N0VyLR67f0C1taOtDulIvWOzzpH61jalB78dZxgsKx3JDmPR0Ag2+amJidnsMr
Uoiamp2mJshYkRQxqtveEZo8q4bcH8w7ib9aliO7XQ1FyLchacZSq1b9dCPYautfT68q/wv0iX8f
DaDdoy6ZUiJpGxvFAKTEy62Zmq66Gexneehkvv0z6ch1UcHgd0Dhl1kxdbcq7yHoQFtEHbA8ETNy
G/Jiqp7xnslT7WIfw2xlWIikJAOgkPX7M+vrHqKVUIE7MMsMl1KvZlUdDLVWY8qV7JQchiQAqhhO
TnHidTEXadHHY+hKruCDXWVd0y2DRmrhBfhB+OOCyBBm/02/Tq+TX8pdmtGL17vStww0nQnH4Sdi
BsnGWeez5ni6FKAOZH+hBkqaBUE289IjDwQuG7IvaQW/kyfS+Sg2Rk6JH1LvL9BeRm6y/Rr+LIB9
rh2BiqrOJkQjeNeeI1CQsf6KIaFCaGN1avVNONHLVGHZCb8uCXhnbv1KRZbFXuR/fbQZU6tqS3bC
FGmEE0pgwsgqhETdyFihOARuCKqHNKjZUfka004Ed4+vuo+2X9p4IbYfZrAY3hyagHycjh9yrXnh
rk71TW7EcYdQ+e3Hkkwp3W0PdcTQB5OL7u3aHq2EmkzZuZoNFUGwuHC+aPzjczZvypdGl8tKzLZv
WjZJtv2ugr9lHDSr/qBSM3qiP7GBgbWXVo0lge3Xe5xOFcYb3FAqWw1GZNGGEEShLHe6JYfiHuNo
Aji4+M+TUuQWRTZIl+0gLCSVfJFbkZ+BduXOv9Pv3tzo3e884Qirm8WVJdF7EKwt3RGqs22CoFTt
LB96h/Ui4cZFXpPyzsLYUrzKM9nsP20TFN7r5dbzOj0aXIldCpPdyLtyTCW+hxaFYSUUzy0hNwd4
7Jv/Qo3P+VsnL8hEfdfkmiriW41caklPUBEtOxcPEwgqH/+sFDKXNx4QvHeYtOG9k+t68IxgDSeA
kyWmjXQKcrMcvxAeMMAKheeVopYyRh3fK1JY7lGiCdl8FzKEejIDYhvl9qtQqasWPXVVu5ZnX8pP
L07B/Otw0mYIiXz9KSQQDX5MKaqQJReGRsPBzkGtAHGqPZvlGDFbtw6P0uMAMC9efE4n3sOddIrF
QV8yqkjvPpuAIX71f+bltIqaLT8n7wMhIgi7LHwBhJJVLDe9rKLxImnxXnwN8Wl9ArWolBA7tn40
rcOrGTo708lVG5Q/qvf+5R0mcSuBc3QtFuFlsvOB+shM/0jdpwaYSTE9HG6wCeNKwOTbFTdpsZRu
tAUW7wwe+Bm0Cx3E0AM1RcliuLxyDoTk4HXILtD+5ucKlmnWbv7LT7Fy/yCxq6iMRO4Vi6wDliv0
DggZNO0P7i/HE+MXdsCBgt77g+GUa/cmoIiaQ4RDoRHGKh2fbAFhPXxwtRm1hnwJ3dTxp1/05eFB
H5tVkAX+d9NNokUJUvQr9Kv9KUWcmuspFmRTmH7LY+tisVuJPlSzEkO1qTrJJV8tTYWDy6fhRGWb
WgJ2+BSWmUjk0MZt51ribGqDMWvYLkcD+MuKt+MqZI744jJRAMT8Q0q6Ki7jaWelD3MKtSw1Hb0/
PHv6Nfkj2Cq59NMmKIRRPrYJ9XB3OYplCc/ypyXd+zNWtxCx/1yF0MxHQW0QHI6dxY0NQKkDFNDz
CR42PYL9vo3F6Ee+DpqgO3qTIIIjTaEe2ssxdTG0JynOF1DZuIoRvOFyWm6Ov17W22499D7EqVlB
CjRL7ZIhADVmq+x0DL5tLKm+GxDn67azVvt5VEoPKhwdiI9ZhEW5uxFHVDu6X+fV0FM/935pHTyf
zJwgWmv2lNd6wtZ9nEb75TaaOENrrb4WMaKkwtQMg0hVH4TwfzurBMBAlo4Ug2bmG6e2tUfvFn83
AZhN5VnzpklyQiBViJJS4nYPs5eR9bWFOcHtyUTE/ecjvivIRGNqtITI70wL8CvylKxA2DExiPSR
CyfP/QAJPW444LhFFgAPfh+B9aeJql2P+y2cNCaFsB3fXmKkT/uxBO50kS76KxleX/OzJAYjYyqS
f564yjEqXuwL8NsjaeS108BX6mT6FWM1OjVSY1j1CCawDxZLdJRO0vI2mRQD/p1TNP6KbDcmHkbB
u6IEtn9WTWZZ8u+1oH9q/Ru4zOc6CTMNsg9KNLbVFQiE8nWj1er0aZ3X7Oa8oD7UwPnMV6Mse61K
yqFNncLlnImZMfN/d+XnfA8DltRXueiyYBwO43qn6s6uvgvGCFFRbE2irZI3MW4HaH4oXc1L/E0h
uIkvVlhjgm5M4eL3KuAu1B4pG88DTJI2T8Hwi/KtZEgrsuz6F4EbFZh7dy9vi68jDsF5GzSSMncR
81tJ6GQ7CXYaxSLEm9NLT7bT7StyeXU+Y3rOa+oK42dJqIk6bRfGOvQw32IeOZJdL6HslkJlPM2r
T59T71RsxDB2KOnawoc76KuM5ttz4E/0R6+1tZ+7WmaAOfpyZT7rh4yXYsIXB6We+8SMNUGjiJ8B
E4MVmQCc44665STByyezYkV+s+kbn8noBHZa0PQd+ygfEIdjiqnjJtAcpfiFWBYhpF/yMuySO0Vr
aM7sYYdOcQSCqm8giZcooBbgThbO/0/vTVra+4yAe6xy3m69+IANZXN9/fyl4Q0fKfJCxPzXsT2q
KNSGv7p7Di/I33py4oJ8AuXldR9RYMdFfSH74CqIyxUBQXjDs/kR9iXi/ztgNhwLwRDS8svwh/Ra
7DZ26fGEsIDf6689DGWUx62yjhh7QgcJ//UnkVmGJB/i+yMacqYc9VReZSmsawJ5G9R/h9/19uJf
rwd6oB0MYNNrJ1ULI0RaSynl6iGPmfdYnjq9DnR4yY5u7b1UodlxdGScNTb6kU+fqTTySzhVRsBq
aKqnuMqvRgXvnoFt0kibd7SCnMdWipe3LsPo8D5xU8k+fPN7HQwFDS7lwBQoixb5lj8HVmTZ8Oec
S1sdunBMyGO9E6Skw55eez/uUVGggpFjtnGCi6oAmqzVveOckVMAP7JkS3f9F6yc2mamR2OEiYl6
zhFEEMwnc35M2O+8EHZgxeQXCyNTT/sIHnkdGRHXow2pKsCHEdwRAhGHk1Gv4Nk+qdHLkJTWNglL
rDaY6GCQD4pXFbDxh1QgI1VrjIzGNjQUDIVoYQSfBoug4NBFch3kNjmceIh2WWWRbvsamOFkxbJh
DiiO0dJZnMmzJZWFhIr0omPrePM0kq4qPNgV74w4ifMLeSvqpZui2Yk05CqfpyJS0+4iAWbQyTdH
KNAMBS4WRd/0T3lIGLKf0EA44BavmMJaw08HLclqmzUJikxZXvFWZGMaBcoJ8/ahEsAlESig44jO
UV7B9uhbSdQKYI4Cc01VoL8jhE6Z9bW6kTpnhtMyPD038heCTNzAQFjrwM+1oIGDuuG8TVr4gniw
aRNXT9qfxpaZbRshtA5CqV1KHfE9GfCvsP9A8SzxQh7+v5hn3sF3KOxnHv2PZJ1xz+gQeHeT4eYw
1BHmcnxazTIVq8+HZE8qbEq9OyP5WlUf54DreRH+5HMafc4FEADp3FOJ+1nd0w6c9Mq4KWJErNPS
EG5McblUEu9W2wYjAiEyXvpbhV/sbuFGIoieYeAXaaOoAdiZ1IO+ObB0XWlcGFllCNlYcwWJqbmZ
/TMLPj8/NNFOppudbWha88zLwjTAXuEfePb6XVCR2J6j50eWDnqR+J3DS/ljVc5czkbLVg2/sWWz
nwR4VxTMsdUIjZyPB3PQPvn9+HlOuuplwPZz3l9B8qSA3e2c8RH5lk82M2HT9gQwMrEvFNMdtXyo
hF1aygoGem4wPbZ0yiNH9uXzjrlFFn2B6SDp9WfyIbtJW/CJm8xbTRz009zSf47hh+lzfntw3Ywh
bTUKTiunXH6XaipcbcPToWk7PDL5x2Z7LvNSfQlV1lWEd8zHOtCghoujOLgUVtqtEQfLetGmXzaj
VJADJMBJLh8PU45aQd1z2poDcoDof4y6/96BIt6o1dlV6AJIixjMMwFFYWVkX0arj22rWycKtHTz
uzDjz1fk+G0oyN0+QVQI4klZSm9rwJWlMRs0Zv9SYuSbIf9UPoK0a8B91mLj2SZFasn+BUZW6hTi
CeRbDEPllPWQoTYOJS8tKcYF4JdPHtNgyXUaeVy8m1Sq8/RE4csY7GTmSUadkvtI9xxY64ZHLd3/
gbDgbLe+C2UVC9MAl8+F85Pcn0Ei3e4laQgJlclF9iWCKfVPa9WKpuBv2iHiansmQEppEMbLrkaA
yk9lQqOpYrPw5TdNmYscEsI9aIHaJaoRi5ApLAinX5cvkKOTBNxzSE7/TPZQFboH2ayTtkQgDv3w
COXWQMGP9qRJFYZQcbum4KLE5dEnm9Af6rxcp+2O3N5dxhMTK1v+CUgkLjIHxOoqPajB/7taBwhG
pMbhLaCn48g7qJiHnFKLRG9TBgQ0YFZDUPS+Cz8pnH0orv8P3c/PzdoCccSc7+1UcQjRSRdzt+em
CEkfjDk7rg0xOajTyOuFPcp6xp7yhFlJXZWR32oEvOwI2wXv/NwluI/NDMtsT664v84IlhfdvWxy
RFow+MpBsvZsKzcNLPtL+XVOJctJtPWyKSzFWJmRwXMGiuYbYNcwwfPdKtnPbwzPwwDJuRSymMPj
YDKnCczSskVM+cT5NG3nvyQrH3SVTfc587GRFuuo8R7Gl4r/+sjsgu5wuKWm+Li8WbCI9RnvkDIe
K62WbpnD2yweziK/ma4XWV+aCnTGRkIlgEE3Z0rYCj6YTo2kAJ7hYYWtBoqcXj0mA61C6LKdVviy
VmycZY+3KQBq4PuXWz8o/OP+SSfwdk+s/6smUkNEPOtVkb2+idQKSL0v82rAj8tTuX8t7FzVY10T
8hKftcpiDA7VcNbOWbeAgo5VE4JRYSvJjNQLqkAM1PIBorgoZhK6C87cPMralBY9JJ8jKFpbCtE1
SzM3+YjZ8mE4ffIQAd8o23XH8SsLv/TwOEU3JIjoDCUOjUlonVF/pFnutkSe0X7dj0RhoIesjfPV
m46by8zQ0Gp7vGJfr6akPmSmSh1/ZqLNsk9xvIV8VZjP2Pdgd6UgqVUEHe2p9Y9nDgfyq55d+0Pk
+4P0/0N+zsphIYSRjTi+JuPm9PQ1h/bpRiP+iB2lQXxKkmACIrGj+BEv+7+toUEZ9BEFdj35u6aq
IEjxKg68yq8bKhoyWnpnad8bj3zRhPyrWAjNrmOfUGEd03IEEOVry5fHIugIBisayOW/QoL2NYXG
CIy196a9N9IJS5qcgWGELvks4JLznDmxwv59NF9nHk5L7OZZvLUSEHUKwbFZZD11oJhEnXMBPL2M
ATHYKvchC9QH8FY6q8dxxcJ9cxCZFjBpKBFtBftdY6rYOOwdfTaI3b7l7eTcZogYQ7BLvAi6NQv0
aacVmrgeNnb76eQwy2EVveLr4P9zcPej+BBKXmoBsjwCpL6og0Kmle6tBVWJFHWLrRo7EIiLzvKD
eFr8RAmbNvs2+BQK/5gfArqVaYeJbArYc6HNvgpxhbXez7uyGnR/F5NNazd8rRMkiUTQ5OKoL+yG
3/SQq7JHsI/8US31NW0SO1VRrTNulHaACPt+1YQV3wgFAz/lSlgbFNiQvbT8oagjCWGIZyNElDUb
mHcEhz6/ZkEL+zDdzpgg6D9O3S2Qnx/aRGio0xonhMj0fHnGzWGVKOqsVg+mIV1P7XRBlIeXlFww
Yi07vCJwtzp1cktrBAf87a9IySGPJpgSKooQTMYfuXSilRfysDEqA82LApmx2McV5NleAqf10L6E
gfKiCLA3vnCi5L1P8n/QowF+bK/LNOElkoXtgMx++cPMU4vZeIrvUP+1aKJuW4vrPYxQNtF0b4e9
5aah0mKW+4qHldITVSCgy5xRkyjbqFGgpQWSpYHQRChFYajfcuVD/5qQgsXAnNIhUHJt+kAU3/Ob
8wvI73iIh9alcRLzqUczcU7V6mtRQSzaOIFDhssGsZOdcf98VHV7p8etucD0Vv/GXWCCJNuTjqE3
7V0ybfoRAMMoqT0yCGG47usxHh21IXjaoAjDmlh+A88bdjbo0h53qA8QbLPns5AljPvioRuv7spf
pvgh9HDZVE8mJHNzNnueUTMZ7q/nynBjT44J8E3Wm6InEtoUPHEJVpo8Ns5+B/5tetLn8ZKZKZYu
x9i05A/ExnKotrejiFm5s51BmorUpRX+ZMQXWETwEbFqo3nbqluwVG+fsTBCDRR2lbBq4WvtuZ+c
xQpcoq3e+yjy4A5yVZ8xR7g72sWKyFy7AkSiqKf8fl3oYnBdUt0Pdtc2O1vh515aA7nyXvZXLwFU
LA1vfSCfkn6bS+OEtdYsvSD/NHIOSKhh4pJksRTEn1yiifDSwsXztaLtMEr5fWol9VsGYHEPJX09
cZuEYHjAYFlRhQk8C9W9wPE0AKdxc0qy4b4R6rT2FUJBcYClsFZmIZXzlxoNfO74YPuIQZT4ZBk5
3L5xFjdz2fNjVGseLUio4zHBK/i4mDgv18J8JPWrafr4vYGadEeRzVYua9XOm/X+V24ONow4TDC5
MV6wWr35X8x+ZlgeBT+qZ3xxVl5OPffeP6P9Kn6CQrWyqevIW8oh44dq03q+vVD28tI+xZWMN9YM
0DVLL5u/++Yb4MUTa3WpnmBppm3snSvm8RqJtbgd5ftEIsie2Ub6bWKAH+ayyFY5wnFarzzGjxxC
NzXnAnQ4otYjEjgE9RlvqYOfGbJsmTdc83ZThUVinWiFuMsMDdLtTlxNPT3OIQl3sFI4WmSXqrNc
a1VRbUINXO0PDsiev98mSoL6ezhcSUW6uzcId1ZEkxY4MZ27BooMqltOA4SvoU+wpyHIJVxwY/T5
d7lMgxiH7L4g1xn0nMNp7UkKph37WG3T36ntHLwfreShfInR3YYFC6vtqB6374skB4zUgTlbwNON
wtLHxqePmF1KbhiL95lX5mQRxDZHy/lJSyvbcEMD7dFIg5rbtuDIHTu1pkr+ZdTKqbXXMR5+58kZ
BGazqiMQLP6Y4uvy23QiIHndRfDLRdcTfH/1JH+0+oJ8w8B0Gf5UQMI9OKL6XpU0PjtQ3IHBKbKH
eyTW0oAYmzzTR6FY9ofLOQo6u+e+qpIfequ+64X4apT6FfM6eypCBfnofCgR+8InWR+BBlEwZGDv
4DDVyEzh8Aj2KJV1NiqyGkYeY2UfnmkqNRj3nWFrLlqRLTZG9eouJBGwADJtcpdtdAla+LHEO19e
UAp+t4HPKtQjmi1XiSHukQlQRxxHIlq9q6dXoD8Zfv+LefhjGve5nUq+wcTNq3mx2yoQapDmMjSE
zvCT+Gq3Y4u7NDKmNCJRSOug1AAZZffyRS3+xTTXwj7qf166zYyef59orLj21Bq5E0kQ0VJr9R0c
OYKOzx7jAgWc7ISlAP3oKT3VgjvkIwFH4zAYYP3uOp+Y/5X4jw47HoiCh8IQW2HnHi5XHXMLo9MR
CXljaQrWgDlvdEMqFxn/piO614Udna2CRazSjW/BAyNZ2ZKpjrsQn9nl7NhF0S+byz+cr/eGXIgt
b91BeLCCm3wEJI6AXOx+G1C0HolLPdNWhNPhvJea4zLkOD5tzrkl6JHLuEk+9A22/VsCWL6AKUgs
G9sBXvr/molkYduMCO77PNqlgPcYQAuhaz0pOwOTT5MtHrJiX0wqqHj2kb6LS0aocAR2EXdQ1QNX
WszhDgbd8a5iQuZMHnHbkYVrNlljmKiQwWRrCKWEnV9Y+nBwmYLJanR3myNFP1IU8MyP58YeiRvf
bwGNVJQvpObyCoymhmxUymmdA179GsAfap90FDqqJWiRJO9P0/XfO/BQpdGsaF+BikFEJ9eKHKRo
8k9iH3Gr92M6OOSvqpUcFjtUzfW80SKZfMg3+ErYNSiSW62f9Ck0F5NENCF2zSX5OZPDT1RYJcca
H/1Wo7gLLTy6BdK2jFJp6YauSHxxMuikOMeQvQcqsJ5qTmqJCkFYy1S5bawcLe/2mex+XaeKBXaZ
Yl4TM0WTJZA+j8N/rHFUaEsNVSC0dJ1tTsBgXg1Dfa2nXoiW7oh7rkhb5jCAYMFBJsQtJPeF+hzk
HBmDy2boVibEUMLtC49pEsdRkt33EmUPsjplRiCbBcgzAAYRXzv/d/qQo5q45PJ4nxB1eN2v6Mu+
4AP8dzNKXay8ugSE1YhExoD6Nm6z5M0pVFAUmc3/tyZuA93PSAZllNTEE70g4eWC74WOn/ZpzM9Z
2FsDk7jeTuRWZ65CyJ3TbUnjjkIdmIzEKDuk5TakVscPc76l1s61EfY9fHgJLcZ7EUxemvVXcz5f
iLgEZTHqjq33ET/PkahAvCpCaWD5i6ytTHRZx7UNNe4xYMEbzy2H2b5wHgGXRo34+Du3xpuOLvSU
p5AEHkn3eS9yRMo7YEIyrY0fyIUZEdF/sbkK8/9SSaGzs7yjHdyiwVCYB7HydVWpaVWa/D+bhHC4
calt9j2o8rm9aMZjzqa59DforyRyNJOCceOoHuuBip6wrxyB53ff6UdRd3eZG6su1qtUEPpzMWHr
OUiC+IKBUcAn3Rmpd3WhD/HEZuYjexj1+Voz7KlAJLFi8GYdPnwe6bo/pBwWUqMuiX23piDI6kam
RXXUaG8CI2hFalTmKd6qoTvffqDqjOQS+/xVrxI/L5S55kHbXu1OrhLYC/f9pt7BjgO3YF6KXwJo
GeZM43pQwKpc7taiZfcDVPS3hxXIx4mznK/KMLnvWCBvJEwI2Wlzyb8o/8t8EK0K3stMp5OQJzL1
xE9Wrvo0qI+s2VGjMpfudQXH1V+tvx7YET9ooCbo6WQ658VEQg0nXQUL7WOsMRcBvYVk/R0wAdsH
wfis9eevcLFKkOBfJvhiXb11UVlvzO/JKt5z3bSvuCeK8zOf0IhGFNgdcuy3ATkWG95MqnDpjE0g
3V8WjYJA/Wn2+5QqRGqZg34WN22eReWLf61OHmf3CVHo2F5gmnwc/2ADIe+w4w1zeW54pAD8y6yu
ZtkXIfFyNINVn2XwPWpLtdL745CpTB6I1/1KVDhvcfq533mSbxxM21zkZo9FG2KVk2Eo1hy6dMYE
Qej62r1JdJis2R6dvA+h2egM+lK2rF+5UQvPK9CBiP5QzoSIfpRx28vymPyCKA9IixLslkBCSTYC
2fkpZ40kybxIVHvANQ1SVptoN3Jw65Yby6SBvZ+FhmMhLQ3TWHUAM7ARtjSiNSD3oHVmzm2QIh65
ZciVksPaYmpIfc2DDy/xlnOzlEHNyQR31yRZCog1FIPPjEeZRE+4B5HLdcn3wh78TDj1o+4xzt0N
dcxmn/xu82UZIrU4Ps89KiAtCn5hSphC3p+Oeif2/Mh9zlpyNUqXbGIKEE1seCMAsn3YKPKBRL8P
oJpHHXlzwJfIM5HgrxLd8nF616td8Gt7yIIn8Tmd0WxBWvhE9PCLDBXyM8x8hIa0OhHHBf17vkJQ
G4926EqSY6/3YJPSFMUEI9RM9k2mh52r911iIc/APMCQvNqeHOuh8gAGQWMcQWIh/SmGMlAYYPk0
UwiGjPukaq/BoED3ABzGWdjXQdPN/JZ14HJz6NnzNln4M7zVRUVqWNdKtQD67RGqGDhCy7z2MlGG
kJHizsHXyP310T3YCufu6sZcRayWbAIRf29al6TVGdELkdRHZ7DkEXXraNRMAD3fKTqEpSXJyAsj
LufFwcp3O9zqjlSWG+MLQAcegpKh5RtBuZANG3PHsRUo5X2zFnmB0L9DGQxmK/FZbxGThj2ndoeE
DMXlWqnqXhuEBMUPyoCczWKYftKIGqDTDjWOmmZWvHnPehCddaq4kY0cGF7cLOIRD9+ZG7MbqM9r
7ZSEMtIPQ+40A89hOJH+igFnQ7pZ0JBTni6I5GFeWeioDWmTWdrMEB9kaZ56fsqspBNTqTGUQPvp
R8TWP6jaUb3K/fNdVp9jVtI3W/v/sFr2tj+q/b6o9XDbWhkS3tD1hEk9tVgQtj0Tc163pJlPPxdq
so21wmLtFVimV/eNMN5ZLj57hZz5bKRxAiCy8me44hpoNLgFwwLYtDqs/bz1RKRhmEIENrnKQzvv
KSjVGeOXb0spcxkpMv0DRDEXu4G6f2FgzZlAxG4jS7BQUB4Dspwx/GDQgwkj/nw4/7yXFXWRKKBP
jtrWTr5OYwnm0yO04eaSEnQAB9yVErAthheYALfrFPI+PCOqs2OOPVhahBzfyF4cUz8147qgsq8U
1QGceIZAw+G8lGy++XYEv67Rayh1bK5SnIjEVy0X+uvB2a366Dk1I2LaRvl1Bgbg5L+z/iAomEgk
tOgESZpzmYdaaCD7HQAYooWOnMJRocj5+x79nJTAq6h3rIUpsU5qMOOWFe+G6/iHOlUUMa1SVVSg
7FXVsXfxZYtyLFK00wKBRDtZ46dsAqsmcHgZGT8/sLaBfvVcT7heKJ9JYtGSbBVKt7O6Sk4v0QCS
ukvgixcVFfdpaxF8We32tt1vkzFW3v+ePv6vfJupE23+2D3XvlAhmPn6qpd0Vm5yG5H1FlztxSvz
kB3HY3ehLdt3Z/AXc/XesMOD2ww+brIN2rbPLkwtu0UtJH8uCvxh/1zTv0vpcnPEvLY4wu41FYKm
ivoi0ykD/OYOC9pwnbZJ5DJo+4+rcuraqIXq9jzeNs5ddUqs0j4wjVpo0BZsHTMrjr6spRyn9w+3
8NeNWqFca7O9v0nAEz6N90A0v84173/sfHoQ8E1TxkmTPQtxwHgStswCupaQ6HUuqS1/pBL2fe6a
AmANrt6N/W6e65ZgLPFzHQBLkjzVr0/Ooj5JOv96CefEYKlANxbmQ9SjfjCDh2qUyGAqe4ND+tQy
KFxV5+NQYe1GtnCK5Ut+q0MjI/R/UQWKaydAievFL3FN7ywHXQT3qL8neWNek9dDuDxhJv+Daxdg
DmUxwJ36ezSC3edX9xMsyhv9ucqeDj5Frbj5D2zm/7fH6Hig7PfAqh1baX6RUIo6rZZgEU+DO+ii
19+5S7HYwc3vcJ5im4Su6Pz5q7za2QE8eebGXmhopvr3lctVuX4ZXQm9YVsOcuRdcGirGLyvvjSy
dgXCKj62/I4iPkKg+2/JohJ4pynRZsACAVpsezteFjfBJH6TPIIpvhwfzLaai7URd1HDEuv5WTpK
MzvYUww9GeHADfyhXGuT+rcuRCcLFXJh+csuGcV0AJ4wwmNdvC0XNkygU2rV8/Ukbzqh7Csjc+F5
OCfs4kyk4jnq1ryLovxBIlnFI82tA9XNOJtJIJr3pUNDnkrugC9fCfY0TMxZkO8sOmkCszhcg2Hh
duQewSQyLBhXSURQUdioVAw2RGbXqFmGF+G3ljkYZfzIAkXmFXdUYSTxVXu8HFt3kL1NdnjqpBfp
az2G6MJhPyw8TKG3pv6Bb7kKtCcjiHMPF0gCjNIPuItsL4KVDZqLb9yjudlvpnpr2tvr92ZiJF1B
8Esw+FLKLU+TuAw6VC9D2/8W2p9kHZRJpA5xQjUVTXc3FsiIfjajUrTxZNDc6v/U8Vqd/Ds0B4yZ
LOoaZxt1ZC6jCyKi/vVeA5uLwSVb1puvlLqhg+3Wn/V5v2agLKjhgtfhpXezoKwq8hZ8Hr+y4AsQ
SXj4QCBPXuaDh8mhG42lYZrzTe9A+9Zs+036/qYagY8ffkEm+4K6rpfjrh56YmIEoXOAQiG16zZy
89D/USL8WjmMMad/Yrt+9pcfrK5orwC9YiAXbOt1WpqezPWSvnPaBblxjlQJPNzCj6O1/qGkWJas
abxqgfPuz3CQK0pmdexClnn2ApoGPbCO6YZg6HdT7VlJY4HQtsf6n8i5I9QSFBePUVQUik0oQaZL
C2PQMGXmJ32RYGNc0AiUp9wbUB56ythFS/i+dves3ZyfndkCYG0f7fL4IcuSGF6Tc4mK11N/uBio
qXM0UlH1eSJ6gfl3Lw3wkGJBDF0vGjrPK/+/m+YmIwhHyQlQoAKHDRJEFe64maxMTrNaRqrbVqnH
PrdtCQBGtNyVNQMvThqbs+4BNam1krTVqs4+NC6Ld0ezujewp/kZeWteaCICZpFPjl13Y/eVAXS7
apOm5gs9IeVn7koqAAuY1YOPydLwRCtWpj9tsLJ9oPc2oKP+JgNmQpjmkHjWtDBwA2c/+4ffo3Ay
teySKMZOfGN5o7HC94JQOJbJ0EN9zZEtKA63fQBzx78+6T5D/IOLdTq3bes2ja/WkIMhuHnNaEi/
1EC5Kw0VEFPh1+vXbcJjvrvZTF1nt0B91KV9ycB8c5wl2QE2rsDoqaLqh4NVMYZ0JnIA9W9xPax+
fDaxZTSVNOOp26//eqAPJGKzKSqPFRce13KH05EJg3NqYo7gcnPBHYNOZ/tth+ynxLl7dPkILzcC
yvsYWJiAOwD4cScP2zyX/1i40uTHg7kO7oSQFnvN6Qe701uys7EnZhS7zloPjs3eEKJgo6IXK4nH
fc4Z3AOME0X86+4xk/LamzTzFe9mZE5/fYhyoRfWaU3y8pX4d8E/GEziDkShhuff8+YwBEnoaTGJ
o/KHnfJPW26mbcnUntqD4NKeKbSCBs5Pp89v0nTXkv0b4dccuRYNDOtdQ8q7hVe+T/driwNYmmXh
9MbSkUB53stB7Yd9bPPzdc/mXfMhKcKQXdBoS+ecJPBubuPq1RyUEtItAecaDbdL4W7tA+BAGm3T
9BoVS9E0fiN/OVYwsc6qs8yOeCTN8bPv9LHzqTI93fA4BYhNcFguLxM8J4h/J++L0rUVK7O+RV6P
DgbHmH44YKYhikNNx4ePNla93MCbPiHnCi+RpJATbEoUAnc5EgTGeykMTrpa118ubrcb7uxDmW+T
bKpF40YOSZ7loR5T055IIHNKOegC546yZnkyWQx+ceJaGrT4wZojU7PivAXswHBcNG0uZbNQnCkd
DehivMv4PYamK4+kt09t2B9rxq1FGgSIaCltZZ380PfxwGA5lftQO6GXrvrorAIFgjb7xd5tFj6t
zOuUuaRL1vrD0RzA5iYy7pTIDBgQQMHzeR1DkUnRDLWdtZfG4DS9Kw3eGBfaM9gceuQkCtyqO4+v
TkhOitskxupYkvnKhuJoVYBu1EaKSByCiIKFLgsTZXGn+AvQaiTQUuzauLRcLjf6S7bq9Hxm41MG
d3UyvX6KwS8Zn7QqD0gwizxu3N0zlLIYslIqtQLg7H7nDABw/e47eBiIhMAtZc2b4I/ZTGvBhEmA
3uupC3/vmM39mgUJA4TH825sPNYK7wT1cE332rhfwdfgOP2JCcFrixuqswhdMK7fTc6KwGJS6sXW
UbS0vw0Qy0A/zUuaj1fshGd/cCqO+jdi7BzXGsJolSuFvxXgBJPhfZMwBzM6uD6Tn7GE9piu6r4G
Ga3vZmMtQnaGtU6kmnoxK6I/mRMWrstkvD9vjUOHMLYHZmThHpE0n3uRbnay/DRCgUyJbHUpxzof
zqBP4ZHwKK8dThjlpdOis9ShgJTtNJypDZzO+3vp1RYV3sqEnDhcZSS9GKQfrOAGfdS0YJtdppTi
i9mB5i4kXPdtyC76pAvw+Z3RToCP0wg0pRq9mv8DGGubONbw29bWHbvYDSHvOOGlXjM7uhfqC3lg
BckpGIfvuIhq3S3XrNwhjmczfPBMAKBWDvxnoFWDs5/jxW1JfWQTGvufU14stOAfl04rh4gop6L6
HwhXE5g9u6SIzai4xhoVRoc5+Xx8sQHYUp9W89dHNXnhF7GuxdLnIRSncTRbHAmlVb55aTv8hvQ2
2BeD+xCfgKAws65cCrURrHiXAvxDe2PQ8DpjFDYppe6Jt6gEFOf5IeyGl0teXKybQLj5jfUtP1KX
l8ZXnP5tS8odXIXElh8KGykdIv9OU+KqUkM97//L9WRE+1DI9vyn+SIOMa7It2UDiudWTJZcZsFO
L5JH5VuKxmlUD1kB8hnQIaw/ABl1l6o98jnl77HK1jowYoVHQG+CSqlnv2wXh84YbqbEywhepn7u
1+YERbqdlvTvX6O6DtzgQDtcYfJxEkF0arq+/9As4fTkME/hfTcMNIlwsfz5VhbxSOmAs95hNLNC
2/k/PeXzKhKBQhKMjKMNik0beSuRKncN/c94QFRbInr3nKkH8/aozm4Y1cjqLO+nF4fe7Q0zoRmN
pxrllpBtaYGqBa0Lp2YNQd9yJH99DdjB+A2rcU1zQ5KAjuMkx8nAOTeY3n2wKksfMFqt4GZbZo04
b483Msd0aLTLiLLBXKJFkHhN5iU3csM25VG1XIkiyh7GWLPKa0/HSTMJP133KXveIL6fUAZpuxAw
rmGIfRb0zExsidOODPhXcaoPCLOsaX3ypf7Lms4JuOfStigV3P5G/YXBnJLTkgKzHs6zZD5nyXwv
dTpy+d1j6bNeiDay4sDRHyeUblPnHHaLXLXZfyv0lLzHYU+W2G6zWVdsNYOzus2Gd3sIYBBbO8re
CCdxpN1yxJ2VZ5xiP3dSIHFEmskcYHdy4u+yvRiQ0gBHG1hIGegAWIZh5iyt7SUSNzTAq2pIQ+m9
yrcUXp33ISUMEXtZcmOvFGTBea6H0aCIPgAFogeuH6YCXvyP8laTvArV8kXxjb8bFkTZgwKpXkm+
8EjvaDICRzx05hjuN0feYutNXX08doh/qk0MBJ3BvohJx53tmikRrpbGNjK6sVVI5mB3Ewsx2dzt
0zpDyH3FujZbhlrITahxxTH9VzOtK58v9s0vJsXRCzWM+GSvK0rFqEZkGjpm4UxGBqG6mzZF5XAa
lZVXtEmVAYEKDFPDn9m+0UG3xzmkv6ChirvaZnCT7tkh9pCkuxykhBLUJY7OwYGGVydgl80M4RKO
EPQoYgmN5TrntJIILFU1pGvWu4kloStKPpycN/qDWl03ykoV8mjwoS3Q3pKtr2eph5zTKJRWKAf8
qVMD2/RTuTlgL7F8+vRhg5GoiFGWA0b8qONVBeAl3h1sPCcM/r0ZvN4iQf7B3dPN02Sh60qd8O7f
prY7cu31AL1VP0QzDYwWZQwNQf7y3po+KDtOTAWBLR9ZZT1ve1AoB2qZsTEX1tyNihrHMkDg46RJ
/EXBT9LICzkQNqFH13CIqd3CHTUtLN3N5xlfq9gXuuepwpODH2w0C0zQcJZPTkknzDUpRQigvzrS
zvHLd2gnGa2V4hPplM2Hyte+kued9IZbpLdTQ5IsgUp2JGmcYFz127deKY+Vi38lHyvY4AmvHrP/
sxa/nVn9KyqcG+8Sw49MLmvqrjgR2fUpxCDCmhQH3dlzpJsuPY0dQwTE0L/sytf9adXjBNDSViIo
j3GxVzrEIZZhB/SLf/jEQcciOrDa5o7rMOWX9kUxi3d5Kbh/fgzRByW8Fl01hbNxKOH7AMfujxIP
qfGIP8WfQeOlLemczJr7GJzlnwlB0PlnO0iC2J8PLX7CLdveBaGDks1PRzDbE4zGnEaZqahriErk
DKq86MQ2EhEOUbP+nqwr0ZvijEcQH/w9rJznqO+h0zyaBJGHUkuj5aOSfj/dwEbwi+Lh04m5lAOS
z8ZsYRbcGtl9jCqG0EZ2RTSEsKHR1uFm+kULOh7rlBt1ye+fUqIHQq5UhH+793gcPzBhJfinr9Qq
SoNlikKSq/R0RiBW5il8/h/cdaQGwXUZQa1ml60CCoJf+y1uYYtt2juwZc0uKa9mnVOKTp94ckKh
+hxPL2tfVc8LFjc1MYQkqJ/uaxurVU6VgR1qFFGWZ3xXvYFOnkhMHyWX1M6pYLHqLRmgvpS8TiBx
mSdn3VTKkLjcEXXKbswOJ8zYXnJP+5cuT2vKCRbPtwyTVZYVOr/3X4Wiy3tJELoTVqPLWRCZruWP
AdRaKA42/Onkt7qwZrFYyn8VyKvGDKrVoHU8e5FIKxHJWbf/FoCeN2cM3Y+hIK4p+on6v208LSga
yO9JmFlFCZ5gqPJtFgafCJ85E6ns/AbsZMyQLvG4wa47NYZ8Fz+BWLSz9rOo84x+LrAi4gIvjqNE
Jc0sQQFL1EHhe4yF+nsDHaxCocV12RkiBht+dytUsInYwqZkU5lD6Dc0hsR4cf7aj79KB51hLEJJ
phMuKPY/eeD1Ph32T572XQaPr8lHo1nH6qzPoDXD4pQoaPIhtM5nY4VgcQa3a3n2rMgkbbyWUYqV
TnLo89F+pHyEAwj+PDeFlny3at5XO7fplIH5QgucZWqBT4fg21+KkZq0G1hLwsAZQVVOkKq/vkyb
TJ/HErfM7MuzOKuTnJRxrq1wVV8suq9CRp/Yh5f911l4SYgg0fzR64f1H2sTgu82+LOnNp4YxmxE
DMyjdmKSs2nWQSS03YETpjAYdCd/VJBuhwNDFdV86V19/HGdpqslVIX3Z7h16h6pGL88RYhPIPbZ
H+z3YSAF1udrHSng1HF0Rfm5gfWSHe3t0RX1DfHt+N36GGD46NicHustMaUVk5f9y30d0zSXJ81X
WXtWQsOSFRMwr8+Hs3yTQTcA10sGAzvZkYqQMH3cVRanf505PIMTRzVbdU2BB8C4g2ZsTOgie2lK
bxbBBwN4JSAUg7Pafl1lI0dWkNq5scxP8EdcGLHBJkLyOWy7N2FBTBHMdyVtVLhca7M2pzK5ZK4l
QOKhlMprjs03jnaB60JiDQJNnYa9ZjSgOxeKLwXW8Pa/2MPPiOeKXzA/3CUQYaDIvXmoUbSF/DPs
NkQ/eERz1hFbAlVxPKtiniBBsR81wZie9tStsUGnx84UiTYnq10WA/n5qeH8a5HAmMfn/0YXjFG7
twtMrgLHJR/sxmSVTC8MWIv4NyxznIMDum+UEEejk9XvCRQYc1IMI7fgxn0OLUOGKYOVNFuqVnWw
F9WDsUxpXJHjkB5ExZW2Vl3hbzYIho8nmYG0MLC1c1iioDi4/+mOBxnqx39GIZvA/Num2m03Yqrg
F+mAACRxbVpxGsxuAUnhNyAkuEkAnxJ21CEL4/ps0zzd1TgxT/6vq6YD6x6kHaGwqP0ABCmpe4Iv
Igg1lYGhvIPHT72pcFW8DLFkKlsHcXKEv9/xViV6mXE/dq+Zsso7ntchf+kP0AIoiTOTswtEOqRS
ly83jDlr/iF4frZec18+Jc0qj/z5Anb2qs3VbbygPMyNvpthw1noaMdqjFrvScgiXVSk0Tjl05B5
JpZdGLkz7nPphGW6OVT7zutPrUW3CeSPVjHcY6qd0AWxtGwTS/qqqzhFVPYYFJN5ZYLuK743DuG5
A47Im2NAS0Awn5Frnb7HqzqnbSEByB+d7c9yMRfRdqD/A3IwvaQf0/0TPZEiRU3QizGnQ1OD3st5
G3KsEYkdjg4FPdmHyfKM8horwVSpNOX7otAej4ogIkOFPeE2QwWsTxkGrla8Boq/Iyeb3bw7stRd
/vwyRJ87jyhQHxitonFMYKpSbnvcq7BxNwe34QIC+PfO305pUfzU5rFpw4R2TnVTVZAXAxuWEN2R
A4J4F4Mm4lJ7lDg8Jj7dgJtki9cNzq+hVtHCXlJRAXo1rAvzY0j7/OHD34RP4e8lk9Nb184sID/x
OHcGzhcd80fa1XI88TONuAZSDytzJik7Q69KNXZ8y5Lsjvjsl5BpJ4XVJLAAFN3+qU5kZ+6njalW
H3gZQXkvsJwU76ZL7xJOEWxq88RWU/mHL5A1Pn2sWKNd7VSxCcKrGfM8VcYJU9hRVyq7sMFTggod
tZELO4x3XFgSSFWJ3ltDc+KRIhIGqiflfFdraNos5LhvUpf4EiszlqivAPs0W9FcIfO8lqJrvTQS
9LKsoHgCiXjWyCuR41nC8hvSuICDBQC3lvrxlFJRTyjHmL7+k6M0j6asG1SdSqdppqRWXj2hFldS
wqBWBw2y857yD5N2mLmVS2B2vYl83iJ7RRDtJg54NGZ9pmut3YR+wjSSCpoAM/T6ksS+pLp3jEJ0
Ye/VfcTug7Us/PrkY0vqZrlVSMHgCtU7+/xG5nP31mMgoHeuZ4H3PqNEsrVztjXa9PPzZDyKVF+G
I5jQ1PvOPQv8LHWQZChhj7twTXqY9C1yNdMm/A1BhMrIU4ekSbjfIcBqTeiVIMRQPDM/fb5EImKR
qmhBAvggARPfsxREJ+TV/xS3SJmNERaC/J2b4B7FqIpXUidGrwlU/4fK481qrxnxxPGpQQe4xmtd
/1R1/Z4aUsetgOVssuRlx3LxudBJsjW1X3LWzorlOmtny57OBtNGFcTmftH1/YXKydrHLq5rmx4A
ZtZoh5lQHsKWgFB/hsRr9PzdVOUz3xyFIAm6Czpc56HwqqqyUjaBvwExXthu0HXOl8SxjGRvDU6Z
hg5lDHEDDPo6tag31sEkVLd0m5xRqny0Hup6eqvZj5ngxcfjjR8OjLdpLygVkLxcPQqYNhEr5CTg
wHlqWEWkiGE7lM/4OX5y4Y7oNgh6frTESGNfuVG34MFIhOVpMfXMkbPliQz0hPNNbvb8PGqo90gM
I+kY42N28Y2Iq4RO0LPt0HyZlg2ie1700eOZFOsf1yRutqov734Tgcyzz0q73L89Lras/N5GOfgo
Nw6Emmy6k7XwOTZ72i64wz/X5B35FptytZiy77oTBY/fyErp3gkbaJ4/rH317Qx8x+N98gMpQ2ST
hMW6VogQJ25by9a7xLpadbtCF3rSpibGyfQpxNGqFVD8C+mOzYetwiFYI0yHZdW2opee/dQawfTJ
p3G/mjqpmCmQn/JV8LQB/qGMXzHlj5AzMqZ7YzmlGlrs9zn+i5vqDWFIgM8JdygV24mgwZ/xWasx
gD7VfPSLaSlWRuDCHuLj6ftFExpwjwEKz83gmGzwHwDjf3K9koub4/ffu7XwBwwTqhu/LcI7N8G+
2gscCwufepL3RLUmt9hXooF2keCLpCZjcoeRkp4rWYc27bKGQdJxNbyI4tIxod5UBL7n1NNx8yg9
+tzY7oswvXigJAtnu46Njo19UGVmHAVHt7g+W631Ce3Tt2mlq0Bf9GvKqT/0lFnp8ZnziFFrpvvW
gWNJs04Z6wlcazLSaFsqqs7ZpOOKWQi1MpDSivtD1A196rRZsfo46lNp/6TzT3okd5l8P08KCdbX
R4DMojarr9hWare3w9UbeJMoeW3jntROy9IBkJWPFJiuZhvAflk6525anEu+nuWVpMKHD69/Md+W
CFoUs4b8dnH0Q5frCk0rzFlXWlfh5x/6ACt5A8UIQulTNKItUun6GQWNE649B4xz4gC64TZZR2L+
65S0JASu6SyOQp6i6pvnopBjwYrCg0uNkgqcnfLrYXDAeRZOPggnDkQqb1w1YBWXP/TaMa2qnFAZ
5z+P79C4qugiXvE+tCbjFHcbrrTbwF3+JXOMbZ7iAvdDmv9G9Dza08BqEW1uasE9JZLVMF32laiv
5uHoQyOEchh1zq7cuVAF2SCemTszPbkBHw6Topm+KUr1JEdbozNJkkEOC4TZ9pjBF/cGgrSRBrLX
jy7DLV/0Irsi46YDxFn0DP1nXn8wzTvAVwZhEDkQdrLjqHkAr60Rzlbs2qS9b5lD70HpHrt5IyYd
E7YUuCMjXAeJwIFirTeyVq2SCP2qGAX4Xpd9fiW+k1fMwG4NmmLH+ivs9ThmP3Vc8i7ouM8wWNE6
qHFYEqwMCE7UsAordfKgApT/IRxyvA2WiLBUeBJJSW+Wt5HBQoTNwXKCJIPHHkBJqpQjeBE0DsuS
WYFFFcUm/kujB2Nj99mbsE0sLJtQrtqUJBwE2nU2DIzQSsXVeM/RGXJZImVIdLPT4IkwGa9xDAsW
mAkDbceA34aPss721aAFeSlHq6i5vSe6A2SCWnSbtsCz2/b3beXMl7oeUNoYrIQ6c97dvHBM2gtf
EbGHLYLlYkKAQW1+7FnU2/2mZOwgma0klnW5hksxJZjRLv/qjxNqvF1wyuX01f4MV6I9tQqWrJih
wj0LNadzbbaqsGZg+/yTk7b8t9lczkLuY6/EOyHFQL0MFv/nbs7Vg6gMHjHvO5s22aTvpf3XRliv
7kHIf/G5cVxso5qnU2EkYKa6ExuKUAauPYtjOcE2WiK5j+AZITg04d3CBe7GqHAuGfYPxL/NgZIP
air0VF0GBvpLrZyJ3eB1TX6e29MJb7YqDdfWCNxFcjh0m6aKxYVimtwIvDBKSTqhRrIN0uoh3i3M
SwY17xTSkK25C4oewtE0x8Qfh8mXBGYkKsXRIQt3eTMxHhknyZE6Ho2sMoNc8kYTWN9UovfrMxGc
rUNViOfQxXDpWp5UUsjFxA249he9X0S1bI6ZeNqflTbcaSWEl8Pf+oAOJvlUplrPz/uTsRKxpK9b
L1QTl11LImc/jmqlfuveA/iEbf/VB+/muzbT0y8t1nrw0+eDynNBsY1igJ9oUWPUX6WGV1bvSjGL
Ylqiyd0YMQN/4Nr73ERSqyeDP/c83XRdYOA6FC2CM3SuRMlX5nwW9tHM0hde6+1XcSMT9SiRpHs6
ECWF0D1QLk+5dZzky6eIwFHWBfTyxXkfxCslxHvf7Ks7NFWjRUzwZDknpoJ3bDQO0awh73I8QVFG
aaVGTnZi0tkz/IgLDrcJJOnOEg/wIQCWyMDCdZCKNReET8dfExYdpzE3xxPZeWWEhOx5DoQfC8Cq
nXh8OCRcczwu12GRWHqBk3awX9yhGhYJPtUw+7adteOVh2OXs400J+wbbuONKYDxWNRzWczG6pJw
PU2NiWdsl3P1U4m4xJSX4qFJaXhtg6/x/bh3lYA+bjrW1wgZJ96ZxSsB9NfQCyVswBzNP9g+Gj8S
BbxiVx458lwSueHHtrTIkvXkFOPg1HEa8rQaz/4qM7D5gOwjjiIOnIVrLN3/yWhf+QWxwkAr7KbI
3Fu7Mem6nrUWFN5j7sk78yrExf6633MW/QpvrMpdWNMw4uPq5owVUVoRoC8MyDBNy7KAfA+HPwrl
GD2izSDafoGzRVbWQ2DcQ34lOANShjO3maIDR1bsQcsmMWUMPAABQOeSPoRk2B95tAK1RDyZqHZG
+uP3x1vF4hDJ55wjpp5N5uiuXafiA3GVN5mNGbXZ9+cCjelGNA1Ub1GsOgSj7QdFq91+RiH5GmV8
Lgu7zF+jURGmwaCEcFEgJJ91LQ4gMZDvHOfeGzfvgvSlkT86qy4hcLnuNfdLjGFcVWRqzqs9DPrk
hQG5FtL4ZjEjF3q3rYA7a5uN3chFsOnjNAjvPrxCk1lnM8NmpXx1LC2Hxyd5tJskolzHQu/JPJ6o
5UaRu0nJDysmcsGA/DfkQeWGujWZSXI3d8dIlMGxBQnIfP7dsZz6VJHCSqRfSoDf+AnrIzHki756
i+qgTh6ir7qKx6qF4vig/ZNJ9FimtOkdt0C5/OeCyhc16WpWpTG5NmO/GE9Pa4f5h+ROfYzp2nJ9
7e0colBNwtm8VQXgvUiKxWHYMN0M2tp2QBOzyAB5u2r7wGZnR2Q+nOZrr/dMf2uTN83MgKwoE/eF
E2o5xPa0uaSPBB33m2Kh1Kf4/rxvja5hrHB5PTP5P5Ni2/4HOkhqiVh9+tT5toD9P5q1ZxpAsp4N
YjUY2yMR7+EMo5WLn/OgZd/BQAfi9hNrpE8q3rf4wLpleBlvW8xKws1kUn4bnabEHsUfrJiKuSoK
EN8RxCGfBZEY5dYdUJnpEDMvY7DdLo2pvw4m+IkO/DR+NeTqUBCTfsRJy4gG1SNfsFJlVi5uigfw
4cHGDRvhr2OyPcQkFzVh6Rw7TOvQmrrnyDCV6OkYpxzEK5H7Zk4sK6BGEo/hsvyjtxxeKI7czQTX
nHu9bvzg/1jSXX74mT2Zx7doJZNrFkU2l+GQY7eAIdTufM49tbxddC1Z7E2Tm+NqFIFHIDqC81Ge
WvTsnx0TRN9uGaGyrDg8b9XgtaQimHIMHt6aZGB8NXpJruSoDaELirdAFx1B20bNUqZQXnpKcI9C
Zry+yjC+5sKFcniYjG5/RJDCbPFtBGZxANuRO6bjDPng3e9aXA84nvjVBE7PU27hidQXLS26otV7
+/zZtvrAcwnJKvsyB5AU9EF2vs+o0kkkLxjfnG818mnpAgWZkODuk4nO2J2jFJ3CZkM2XJ4OwQZb
XS4eE3ZeswP89arpaJ2r6mm0RzH7oHDrHr9NH0YgYAfNcNYAs6uV+Pn0t5gh28kbTz8YezQXpp6D
ajp0dA6+H8/L2fIeON2+FKNXUuKxFt6ragfLdQC0FEqQ770BCXIXEDhdbBVeVRGDoGpdtyvwI7ks
/vuE+YBTFMjp8OMF+PKSVmiQfWX45hrPPErXjSIoQhtp+cWFg2LiBp12ciWaDwM4fhr3zAD7lAXs
erfIX35OgMd2G+o3nxMXjcqAvHE8gaCKQgqFD1Vep631oy7Ib56O48yZLgQh718Z4pKTZMx0cKr2
49kKBjN0E3wugttux/Lr3G9KpzoPkbtdT0mGOkaYDNkqIRBA/VJMnDAx+WEGHMpJttFkNC+IWbwc
sy77Xdyz6F85NmJd1P/TpP26MWTUbNrYUAbM2X4iOHfDyjI+NpE/J7+b7X7lwlGrS0Th6dX7N6E9
VufleefZkAy9h16OSuTiZ05s2WKYxCM/8csjaPrO9YN7L0FI3DsIPLi6zQhNo2Ihx1oGTYE6BEeh
ivV1tjrYsu+OwnpF+0WtoQ3p21Ubk3JRPrhW2N+FvSBaswO98Fea2si/OHiidsBwvm6gq2fPE+OA
0C2bra6INDydgxU0L5CF1UReVIsVxHCwqM+bAJiCBMOw4g/eS5Ji5okJgSBGW+vi8hS2pdpbLEkm
i+l/iTa/MSH0qvBUxr3hoyBnqSOfZEAWcJXnPCyctwpo5xUmsjvV0Cv9BsZbfXQK+IzXwXu5mwPz
xYMOef4F84NyahTCabHxw1xlu12XIcGN8fpiwUruzx60eTtJsC4d7hJKB4aSW+WAly4BoqXmaIBZ
1bsy3PSnNw//y7/hbNuC/uG1mHWKye1guaUoLcUe9YOBL6Fm1u2JYmTiw64UobWkV4XAYe5W4AHI
g9cDrnlLpc9+U+o127I7k2WFhSf59ghYpw71yfK/YDOx+NUfM6hWIs1pcxHrBbXfjVJU8Abpfbwj
HptoFKkYIfN4UozC8nWYLdsZ3sp6tfcBvQgk/VLNRlQvXOJ3X8cy/RzGn6bcsVs8XI8mPufbvoFd
xO7aTNJi06yFS1LJwELLO5M3evhVtVlP9YxZ0sTjTzR0JTyqY3YrNBqD18RY/k0gtWvxUy9/3kZM
M4bav4S3TvXz0OmTU+okZcel7u7Hj0s3TQRr2kcPg7nDfbUQvdVqip1N9wZOA9HAVgHtt2WB98/i
xfibFKUvZCvQjzF17KYmzEFnhl9UEa3CdmJJIvJpAgkdi8xxPfHmvWnJvR9kVUtAgLCctrYKS0jW
yjYduyzpvcGzwXQyeUenBWc/kds4y+jMmNvuJw8jcVGpiEO6rm+eHHzDqM/i9TZ6P+69um37ecFo
PhhLeHpEJ2PDBNAy1clunOFBUTHZMabY56IgxLWCwWq4klhmjT1XlnT8281p25+oouH3MoHlfRVf
ZJIj79EheUxXEfVbAvXRyERlGRtvl2yR4qEdcG9EtcL5P/HDN6la651Aiu3UdgvSeaisFOlJCsHb
IjOuXolWEWOLs4c5W/mnbJkDdtDf1XSW2pDTcxCby+q4tiImdppDQpcHSRbI/u90A8qszQqZ5Z7V
4Ikgu4nEzfKtdLXKKRZLjudKD4/0QuBHnI0lIxAPRcOy+iXZ6AIVNRe9IQVjuHrOVTEd2NStzdtP
gR2nmKRFox2perMkbprejKdBzrk6cGOJDsZykJ2gLJlDUIElDmRSWxO/ihm/EpXNBhykYgBRf6ya
4yHTd90TeiTuMeQts1S98sM9SV2eG1FpuovNX62B6QkpXU2PQdNPVDASDeWp6RlzxTpHTNXF3zyk
IoSIpmasD21W68x/qhlJn62F6P+dG3APurYUxUFxjHjqYWhsf4n34ZltZWbbl8nabGuOZKuQsnGo
wCz7QTykEekAgvbbEJosTPCZeOjMFMOaebVOuxve2MYzJ5S7Lse8yjP/iR0O8Aqh62QKsf0f8QQw
dxcczd77mvxTEFaWHa6rFK8IptgC+jWqG9UmWAC7ZdK7VKVByYI4vPz35FNH5nNZecILG4M+/p9D
N7hSKBad4dY34/PCwEwEZ8XsdkUPWGTvntiXPIyCuUOGQq5AMS6dEm0klKSGhWGbEazA6u0jUdxr
rgF3bKwgzBx+Tx/EGHYylEdTLDwEFxELIH3KRWXBeAM3dEWSLqtB1I5QtT9nFGmvWwVDxtX+MeWf
CppEJdJ24uG14gwOid2OMzpRIn8Lb1HopZLjn6MpVQC2lXuflSiPYI4OMMAlYAn20XBzm+iQLTbH
Dq7Wkq5NIBsIXlmbJcHa8lHSdVW5UYet+JSPmehcS/NNWqdTXCPeQpxCqBFWYdnKJXgojvitGgpb
QqCd27dHE5z38EuOnCIDrHs/qaV3Mlr+o84QfcByQ9Pt5nFKlvkAAH2WhI9myS4CbjMlD2LxCInv
LznSCl+niHOCjjMB/KkfrtLfTYSMYL0qJVKXSWmDVwx47nsBFSX4V9MozEysMem/8p2t4pZW7fwJ
DjSKLKbxUFnT8bBGy3zRGxTFj0OfVXCAHVrWiN/x1EJLzaZ84+3Q7/oC1dfLOhhzuBQdXQ3F/6mG
chDq/7FMQMtzExcC7RMRRWI9LYEhtBpa+Rq2urP2h7NCx28feM/72V6r9FpBfqTmQNwsUzcmtcJo
bwiowjlmFSSsTgE/p7avWmANXj30Qs3LZLuzmmAEOsU54sh4UUGQeNQPVKD+80csN9jN5PRN4I/3
pdEfZHWVP+IvbKrGYJGTjBLmXUatp0cnQanPUs39kPZDSKZ3giCPcilIYxKrjfE+U5NzhJOfZm+x
LVxl+pIRZrxC8AKvnwRmwvMqIltZfQuCOq4c6yztD2qEcfYCa+UtNcPZKAMPWnD9tJR2RNH80shi
0/XOtP/HqmruIOqi9s6hjES1MgPri0E9abYP7Zf4BtQJv9PbHAY4SlcJopU788suJi5qtQ7aTKoI
/mlSI+gHATwCl7SRmNYtMaaxkLCONovJ8r5VyqO+cZ8SRs85/bziSAk3IyBTBvgHCQPpQedBvOTg
xBczKEDL8dB/1mDXxKV83NubwyBFkWoq9dmzxL6jGBtVrNRXUqs507EiueGwM8TbYQufsg35BBGk
Mn8kN2i89O62VOLsVZD4YPQjImSLSvoj8zQMHgir6PzdCOBeRMorI9/CBV3H5YGzRV+3wb7jQ/Ei
wR5vVu2l3SvfLktdOkTlW1c3OGpXcMCElSSnLQ+Ab4Vkce74d9KYPYxkOqanefkUZn6ZqzEs/z63
CGbFDHEqWWefsWX4EvUDjNnbPLt/T99YNHpSNfE9t+xSoV5lVVHNGxCIhu/PKZ/K9pB9VbDqYzc6
/HVkt6fUbPD4SS8jHvkYsY5JfW5WadqPwlpcBcT700BCgk41cmFaZO942Pz/l8OBmTj79MBaDKVa
477PV8+wCDsM3iv4uiSK8GCUdsIxgRkYfynt6714otMaEYuyaBetaTtfOmvT2gMS0VYS+/ea2C50
cL8kVv/RYG+gnYhXfbaELggN/j7oGq1Drj+MfsantWZD/RLQ0tjCBtqHVNeIJ2ljOxltsqSHRHAQ
DPCW7bFdI0+2f5kPgjxWNTZFcwAmirLwBfRLcaknkPvVJMOGNAb8O8U0Ko0MP5UP1FFliezYxLo5
mqALYjiJuzKEQXjiBwRiK/TuQ10PCy19HGIqU7ReKeldNOs4CiOnjXMmLHSjb2aHFBau9sv1mWKI
qtlmO6CS76NqIdDebAfUPylP75jVQRdgFWLi9HA5yt/WI1VXRV2xcSkLBafiiwgzelx0U57VgF9w
30RTus8ghiZyBJaTmv/Ak1RY/KT4+Z51zqrsNUCCsFT5mWmIIUfO4qJrh4yHxIS4p5DYvtG93GJV
qrWNeHhWfvHX5glXekm7Dpo6Zw6B7ms7nyYs+A2IYV+HspLKTPOj8HNtWFatHOvEP1Zccc98Yw/m
7WM4h8J1OQ5DHAAVgzKk0J398OMEGMfemqkE+PfYaRjl83TzqfxaNVdz0dxpiK4LgM9Gpjjgx4Dq
9J8DYtXKPT2rBwkjgNoCEG5kgLO/jnRzKMBTksBInK1OgwqQcIPTq42I2z2EoYMVXP4Zhxr6Q4qX
ixvVhadnXKjLpfuGv5HISkQfsWsFm0mcWmm66VyGHSBM3R58yAEE3SlSxR0lhWXZEHNA1KJSlsKy
+RzRhS2js7XN+crxgpWjxUbmYW3e2D+cuTI3xtARMH5JCyQlYH+igZ90W77Qd7+wJOy5CHnA7z8l
WtLjAwDI3szYdmEnNmO9gUZTnlrukVEFv6qHDoIAvBPwhIDhKBzlhtujMmaKS08Ha4PhCh3DHO8G
iDTIVtZK5IqhIZrNDVkR6iG8dC0mpLzB3t3dvS9/Kqq8fBNjkE+WgsP2k1pPSaQ1MNZMM8zHvrnq
ApXfdOAxXzXDwji8Tnv0NxdlLNLW0jkFcJoXXe4x/M24oOKmQDeuP3zYGMf0Ye9E39ttxH2BKzCS
CeMlf0mB98vTbSlrK1nBDP3l/h5dkvSwlfU4aStXDwUYSGEqudeBIKEPAQx+2PII21JMRDnHlqWD
YGuGukkCGEKhNDvvIeurTq12fG/0m1xP3zTJH9+y7SvGTDb/VKg2ZsrlzfotRY/0shGTKaobJGcx
7SjMqgMK4HznjQtjKm6g63Jsialn09bkVMW3FavYU25+nkCzXcXg1xWx2YqbE6osFQFibl4jrJdK
Avph2Qmf5fElbh0/QvgOSqUvBxuO/ZUpRGSCpLazZ/EJ7CZP3BxxZ4+Inmg3tXKGXMfVgw47FjvI
4/KYRQTXpIiue0cdQlDgofuAvoNXyxQbNrcX63iR293DVWRa2F4nOyTrxlZ6qi341IgVhk6AcC5V
7RDcQIWTox0NxcAC12d0zNRHKFHZAckE5lAj3z8xME8XtHgzFXL7jhuyGlSlHDztGhAfUvmYc1Vb
lAChZcFn4SiX0QmWe/IwAg4QWoxwJRuhkCpYB+8ol64/9ufmqhYGPiMPuFqYGKlNm64VRtm3NMkl
wyGKrAW7MO9ZVQklO3wIGc0ZgvhiTvn97gQ2l5HnjTyC7bL50FeLwLbGk47RZHnqKSfy4h2DAr8c
HIeC23LYPppDrzOTNpjCxHZNRFj4KNaM8U/BLSqmpKajbrLNsZ9FJcKyuxQpePJlWKIbWycVJODF
kwvd2dt2ePIywgJtp6V+wHz0Y3ybdpdIKlXEFX2lZTFMnkYdzkY1lM0pO3QYG0DPlnNmrKUF82Zf
/yqgGziBJIsaygyaNQ4C1Rkk7TquUc+WacfLU+QOxdlBGy3v2vvuSwUuvrV1EEi9G0yVlItWxVlD
A6uugRYGWaG/l0E0QfWZpKAJz0N1vdOawl1bzJjmFeFKrnJwCANh6MEFOL3wBPLcVfFRZ6yxvgyE
EtlFHjVMKYIdgWITORRep/0632GH/qSC9+SGb1VYsPZi76HGiS4oyOxU28/TTXcfyY1a6b3vRBdB
g4vXtoaIFqkziPdLiG4ho93hW0vDIyr4oaQ6lD2XFEEeRjanZKB4OwbTd/EuFczxdGuFQN6KreeW
1m2muFXIJkcz7QoKrABQXHWW5jcaw6MN9ZCFQVm6NbwhQbGHjEyUaDG8/+1Ay9Dv7J775W5cWxdm
b0K5a7LMOdwYJjcuR8r6SnjqN/awkTqEZdOj8kwo9TQlDDD9GI81Kk1hX+v22iNAH7AfShwJedyC
bm8h2jYJx+B+vFA8jgNuvUJg4v7Ko7VpM6O4QhTHkDzpfoCyRV0w90BNlgya+AsNjE9xhlp00iVx
R7YbC/AB3OR8uJQPv9M5VQh1G/kRzO5+c5JQVy+dk5diJeNdDtfq/u9rt41cJIM3BRmccy/yQ+BO
YmFphDLv8ybWSu1HZV4XakTPP2iBYI7DEeIGIjBaO6kaHjLh+klkkCTjFzNpaGIaJ+Id31KPV8wn
5O/isJ7aaLGnhCe+mIu+kxul/bjLUzkSpVh73iySqVcqdmfeowmPQqv72U46q/+ihdzc3kWPsvz8
bGPZgxgHOqZaHgH3A+vpzbsxRCODHjJQAmHXf8ghqFxwGZ25kkSgvRIkGNDFUWw4NXXkISKO3VSF
8XQUL5vOVNXGYY4GykXQRg4a7pV/+VzVkLS/obu8g8yL5g0FTib0IpZPcgPL0g+1hZTGrkTVJx8B
nfYO0XOxW1vQS2dmKQf+0T5AtMsk9K9oqxaBxHaDQKjjm2gAFrmDeDFDxCuBOhtSikJUzXN3yAfp
zhP/kjt+z5v+/7qtcAdENDT0hsCEp00y41Yuy8XAjAAFVIffSf5kcWB8m2Lfbv5cxAqmY8/73SnU
WW9oBakr/OT+HRgcFy/DBMPjFW/+3+oj4/bJ7MeiCXe020JFkNtPGnBaYjMCOntV/MunR/SWZggP
s3wJDGKeGz089Za6eyxfhe4zK+cDpcXcOTpdGrn+xjnDehdDgsPFDkulpBcpSXfCEPwzeCUgm55o
cKVPNtBTsOdycNKPm9y3v/GeIQAt3a12JvlcFsNWFUzHauT5cOXv2MYWjkgIqcCGH/jau1zx+UJ6
JAdlXzsSeD3O9d3sy/LDsBlxn1+20T8jGjY0Bmcs5F9nDNfHRaQkILiBXl0A+uF1CE2yWaP2Ctzv
NV5qxh2sySoEOxixXDIXrTg7UcFWflosJl2nNlY/v3ERVkw6UF6xsBjKKF5jpQvOf/VOYTskREfg
vLPWnEAcnhFr9z3YhTeZxVbngObdFYM7dhqYCJfT1A/lPFNjfk33m7HqSeF1Bo7TWBX49OCW63D4
etAug4WnwKJF6X2h8xV2wK0XOhyW+h23wLWHu9qPks9cqPNAFbNH+1W/pxUJvVzVBFAZ0TkdLtyX
GRCprGe5SnfoNf3Skzj3K4js3IoOEGjXP0xs7D6k6zbIusW4pAvfD0B5b38UakBGjdskzNXgCXNu
gnhtB0w7fSuCgHktbUpy8QeihO2GPYWLdQB5XOtSE2CHNoEChn68ft95YGEqeTnw367PyPFTJ5gj
7tJ8uPVnqtcHqi7ncsJBs1diUuG+0wHZBnOUvO/c4QvE1bt5v7O4Qib7quZpPPP02jXSlEu3eo3N
mrJhqs5D1cvYRLKmAXZWFBSs1GG4NUW7EQt5YzuazoP824/jvVHiKmfeSAtiqMZE9wYQKei5HnFQ
EIKRQAmQIxgrFYc5G1NSeAMVY/sei9vbusGB/uUuKgBSab8PxsXhk7ARD3fbji88L3paKm7ajTua
Osy0uwfCwnriKc6jv3NjTitkJvJxpYJYfRdGSNp8AWZ9o6bCyU+rNtNfRDfTfU1GLowdcuJgXv0J
iUFvyz1AqauY75z83fTMiSz6V82Q1CQE7QUe9Eh7Eo0ebmih2b54iDCfbJe31IDw7ycExaVuGIZa
uDpG8dRvzyBbVchk3Sa1DuV8C4Ouq6tpObd4UB1Kfi8zMOv2LT9/xuv29IMqmvVzDVCSkqBYGJzK
8JnUaWQoOc2li8B4+WyLiTM7wDH/NHsWupiR5s1oGrxpg3ZDYprXZuID0SV8kdKDTwyMREUX9wYk
BKnXTS91VYuAXl2hmzgsfC86Fom3cBDcs0mvdMM//n3LhcmsjImd9VLl+okVxik+2TxWWx83QC8v
SluonP3DE6SWC+82OzQwWoKsCpW6nNBHTVJLkd654rczvsQN2U9MH2yNOcu7a7x04KKoXAkh4Jec
60GJ2l8N8eMFbR0vysg3icPyHoXKtRu0dJMNxoC+uIcyG4mJvxfu4kLCQsNJG30EmZsOvq60VbyF
vNfnBb1bnwwOTcSzX50quAa6GlpAboY0YbuUTKxV8inGvRSU/Rn3BWBxsnYbunoRgkIVB4nssos6
857SnYX75xRpjjfdOxtrXRByJBryoVcRn2s8DfdemIR+0Ta8hgbyTqVZ7jSsW/0+J0+PzCYTainr
jsjnMg3msZtRl4w015nF14eJBq/eF9fjBlMhdaOYFwGXvZT9AOMH3RFI7ABgRWKiAdDn5sjLGyYx
uLMVkWdQ0PBQWuztUMt4rvd0wHlI05XmbvpOEXzcOa9zrBF1m0R26Om1qlHKa6pu1uQ8i/xYx6iZ
3UZnfn4L4WtmEi/mFh8XiDmLecG6JcTbtgRc0F0dzW1DLAeO/rComGceWMMAX7Gc8xd3GaF+OWmV
d7MKf3uy2DXF/j5Oa6bvBhv0VuJ6vtxus0ElfbXeiQsYPb6UvekqMjYlO2zFkuUk5ob9lJOr8uAr
S3UuPCAZvE3IALNk7Oo8OsLg5Yxi8i3brsqRRcU7UDhU3n//lvbGPXZn62rbK6CUSrSv4bntngbs
lr3TYmYISATGwlB2ut0BnWLCBjrxcgNi45CQRRsnGYhXa8jSEyxFoEMvAUmZdKraR9SxZcr3BVoD
tPvJ+HfQLkpxMn/gjAm9GLqrktuJvUKCpTdAeSrtRnSECylhnMVChYDdk+olNKZ7Y4ar7dbzK65k
ZuYGnGum41WnlfLBDo2tV8VKRnF3VjT/ufCYTLERY5u3RhzJyqw5njuPduyl3mYqqKrC1F1ZrgpY
VRh6TkF1SCfNeUeFJNSaxgoJVH7b+SNwE7R+i2TaXGOLemwt9kiNLPm8TPImnfmRnP/feA5jj/Kn
QKTFqYzORxHa5ATjYov8HXke/L2BLYV3su3YJR2hJWQK2RQeWNgnLf5jeV3mqmjEja3F0VJMErib
vq7wBV8yIoWVZ8QWC5F5XRAm+bk6dmSmeCR7aDiQIY78m20TUWYoIt0bKmyNHBIfYeM+zOh01yRm
f5Ls8w2/G1GDNhOemO5HGR6y99qNj9HC41HmHaYL8J5dTmmKCjm6O3M9Qpb+pQUbmQbX6+F9NeYI
AYGcpuwQ6pNR/AoFDRICWArppHtBpOGVGY7jCDDqaGfXIRxkcOfnCXEeNHvH2YY+0a9ppBCC4Pit
ThVgAfIWRCQqOkaPgtBOEl9PngyZvdeWRE8WYN+X9AV/yYAQv72+cg7flxjhvYtR6kbWVvIU9PIU
e7d9UtDOQSjHghezWowZrQ4v6/GFURPe+8HGRjZ3I7hCRc5+jc1Ff0eld1s5ac312NzV2cN/na9f
LodKoNw95AR9TfKDzj8tDNMJXJWa0bkIDKNFyt/5jkRY5wIcWh+/nPbmzsmHlnZwpbDGBgwi+30s
lnt+1F/Qtb3bRsGfYqoPODrrFIkkjyVz/hVo0KWI/xhcqIP5foTszhWY+gxMUalOnRgaT0BYxZgI
3uwv+LGdJzV5en5trmGIk1orEtE6kOTl84G/HCY9UyrxdRwbQLa8hYZrJ0ufmNxqrPAbKnUWj8Cs
IgrGH4fC14p0j0+cMVHIFhtQJnoY96/6dvivxMlB8rIMRnYq32rTEwega0is709yjz3EUD0R65S1
X9/kY8O7d2dBF3lj6qmc8CduE59c/7GYAXC6VkTctAtjGwII8tW7v4Exxj6mGF34x8k1dBholTYZ
2CXqMAkkIsiBiQ8yIrWcB0NzvJzg3SjdrHGKFH6ogopNYa8Uuf8u5eYU/SVNqMmgOLCXqeuZXCGS
XNIEQaN6MVzRKR6SWLD5JU5DGrrgrJ5aN+4YjXmeBYZYXHE/YgrUirY43aqiAfOqRngZq1mEr0MZ
zLBYk5yJg1lpmXLJXy68ucS/yaj2evxUiA+UNH78iCrp34rY/sA1furFTHIViVEhx1iGGXCA6sz1
+WhJRVki7PUwKw+mCgIK8pIwr/t1RzvKq8uRM1rvv3wPlgdca8aR9SHj2jsgkpk1GwyVqoXPKbP+
ZEFOXn5pCXEi67u/pPbzFjROqKHT3k59/ZzZFUBchA02WxQQQzP4po8Bmww+HpYDM3HrUffNbkdJ
ld6v/gbSUhI899K2rrpvkowWvO0Rh+nbq6dqmSluhZKpBXcUsxR0FSZ2/Fo+uKl9PPD3azx2dr4Q
+bcUaZ931QQ+MGuE+K8/oq7CL0KoXPrBX/DNA4uQcsyqMObY3mTBw9J54PBFnpd4odvNdsipGtS2
e19Q3SrmWhAqrbkTamcCcRJnljq7dIn8CNw8NurUOOng/Twfw1Xg5N6SzyabNtG6dXNsGU7x55zd
dFB79E8U5c+d2QVA1qLJey93PVqzZylp5ZVYRGmL/Ql9VKulONy/sv+r+NFEaR+JRsIsxA04eC0y
qU9Rf8UIUllZly3x9uYe/mYsTkOSPQrD5JmDFfJ5+OMgdN9heJ6LQR0AAe6SCmRBdvRlv5kp1Q4P
sEEvqCrUjy6N/u6IDWu41r1sCeksC1VF8UkU8Sg7NAs5UWch8rQ8E5CbE1Qeug0O/4fUdS77vs7J
1vshNFNH+zlvHevixv7vuhAbVa0uj5U6tUmPFQU8gJHgFduyk9yibAL9/vXmO0+eNyZAwlwVzz7/
rF3meH2ygz1mRmK3m3m4OOU8KkXTYZaXwa5rKb3t+DC5m3Uv8pUeaBh3j+gTSI7Wf/B3P6LzYWey
mrt7ENXNdf91ujIvBtD6fGMdW9L8sZ4QJzc9L7nLVlEDQ8C9D0WPC9WM/xBdcPegrS9t6pX6F+g7
LuPP2x1X1QfeE43wyCxHHJmAxqRwzZQHK9M6wMI0eAJR3Iz3JxncuQr74lixQ2QfIuGamaCe1Q+U
nbGEXDB1pTMg/QHwUjRkMOr/wRSv+G0p42j/x9dtM88uEtBXo0KyEZz64zThc2kHPB0T9/4Cnnr6
h1lWGQxSVpsu889h9QKAxj31RQIyhdeGjILqHOiiQKyZkzk2m+5NryAMTT6D3UT5UnvnOlHe5Md8
P6/SI6M+jirE5PgrSz/Jy0yAS1Dwj5Mv7JOIImoGhiuHGDttvQ9zT3gXwbH1TK15EhKnftFD4Cwk
SsdxLxo6sz/gbpqslhioyuWmrzbiFG6q6lSCgRdUT0YBVkDkbQYXDi0K7nbJ99u3P1dJs/WnHY6m
8X0WFJSsEunPHgYI+YoOYvhxoSArESWj9vVaNNJQqIMokn1RmHcw5OPhqO70Jc8QWCfjLXCZ04CB
jyDOHP4AvMFbeqmndxHP6Lzzdo4Ur722egh6ybAd55bc0HPM5xi4JLax29hgGj63Gv5o+XBT84+U
7LX9bsjdB8gkyy+mEaYUqWKLlvD8mK9krJS+zQx7TOd0EKg0TxaY8EmYjTjwDvyC0rSZ1lG5kgAL
PemD6b3Wq3+5GsAyfjEcsNdcQRPaInL7IH2zDepJALn2N+b8VeSFBV9gK/PVyAsjBilzdDX0wbv3
LCiVU6pcAXdel9g0EaU3G0nkoqn6y+Sj4Cfr59RNt0GlyyDM8MNDyC5Cnhdt99z7TdhjFWnnr7HV
hpJeQr9j8bB29jt6tHcLV9/Z9yLwfKi6tQ5lT1EJjW7LQdM6LbtiA07Be9H7Ei2d3maRt5siyyK7
oc2MJqIKtuSCir3xo3D1hg4hpDLJU8VEwn2S7fpH084sTMMjMsYgA6bb7I+B3nGavRytL7zCRqR4
PS5+nSzB4pvSREsqknNqwTy6GMguo5EPs608xJFxUha083bEANHFP5LUb9a4Vy8b1d+ihu7p7r18
R2T8wlTeGg7KRatCrDatR0MQPS79QhcOPo4ZoLqQii23IMAWyTl1KImTmIPKngDLllzC21EjhVpn
OTpCXC+CbIJX1jddzEE+WqkFtI8AGew/b8/6tNJe/m2g55DqFDUCXbHfzbL/Sa4iD33mN0+UDz9Y
frJ/khLOQgposbuBV40MqfEBToLu5i+ElqrOI86Np8C9CXhAJiJea8gmYgmVqwzsBCqVp9PJEwwx
SkjHNA80rGG+mBMfjZ9q4VoGGH9cJqlZHdtrGLhWxQ4gyrowjtR+x9utryiLJx4K0XOFqiqgCBXp
nA2/h6dXtft9bLWSKXGPUW5uwycPJl++KKWW2CplC87U4LXhWPNH6h2SvX4p3SEIJWTTbHGuLsZm
gWyWqDJq23b8gFCGFmvXTnqsz4R2ULJXDKMqXr8/YBanCd3J0axLOY/kf49kKIHiwAht4d2ov5De
+WJQHwcsE2GsMjVHspaTYvQsmjj+vF/c0f0PAI4cBpac/K+5HQyLF5cE+8Z0ces3grIJVDsTFGSx
g4LXhUDXltf2yozHJxjkgR4WUpJrTrp8eUlV3O5LyS4uggV+DUOhEjPHTC+CN//8nDvG7hG6Fqks
4egiJL/xPH6ay8XlpaAl1N53sWTZ+q8V85Y+CIUsxfXIjk3A8TRcpCG8saXUx9tsnn8/KUXS+7fT
FlEZsw9tJUEcvmEEEia+e523WwuccIa/RW2AWD88DBRm3sBRa2SDcxWCtv7jacBuy2jODDllPllE
/MNGnU2IKyts1Ah39MBfooSSfsFoNhcCmisvuRzJeqgOkbaDolzjjupatYtPQmVARS8jQFQ6qOH4
c40uJhGhsMgaB3U3EhQNvTra0BMwpPAR139ZNnLrKjlKm9dQRqaYKjoaT6RpqjZ+u3+9YC4nj3Ds
xkz0nljZv3M2Y65Khu6VDLEnMg8J0dbfonULTsLhmBKWvWaBGjYZQwdHCzX5ukqvQdHtQOpqN6ZN
J+Lxiktag9E/UMHo7AuqMs9JVRwTz4E3fNLpGaV07/EP8X3LuG+KAZ0UxxIQfAj/d1mwDTpEtyEX
6hA3NP8FhFpoylG6ozE2fRvSn0t2V3vmUwvGsQjAnOGFMJpq05dEggPXc//kl+SoubmUc+zPyBgt
b112xGzk+RlkeR4xn6IDir9y6hw9hxZgC/xOp9QlHsyNSt9GyqGigTarBzSoGsXH+tFL8++aoFId
hdSJOGeloB1B6yo9WOlcRqiXRk8aSY69vSA5FYERirYRmAp7fP7DOfisJwsZ+MOY2HOn8kZp4IH5
SALdNUwrpLDvMauNP0Tb8pjXWoeiekJkhh500uUk8A45aK6A4JCSqQCzUTS26GIKyMy6Qa9zKpbS
FLWZ9ug8YVfQzWWMywR4168Z3C7VMS6hdRcwYET11ZGe2rZtBp5g9z/Rxd4+m+QgEFrn1gStBh8w
m+ju9ZL4Tih/NzQSUuM+ys3rirCpc3oOsfMAE4f/z4fQ1pViN3VyEWzBmHfewujb64sGYNRNtrE2
9CJvFtCZwYflvSLvnPVf5gtNtBeEtput9BQ1mxaUiZgXt7c7eAMU3zBpnd2ugbyLroNseQ+19Qev
hVwXC0SJe3L8UFY36V0V/mjmF0/WOxHnjdEFzJxCXxYW9YjLG3a8NP9riUYdF7M8/bmIrJ3PzTV1
6VQulzezNqHwEvavSuUzxOKP6FfpuG8oAeuh51Mru4+TKYftdzwtwPv26rekbsYB30rcJgX3GaOx
9Zt9HHCzYo+qm+AhCyNbW2wuav3GM9GbOHdHgcKd5pC63nbTI2hX5y9KEfwgvCa42cvhV0wlBklw
nqVRDYmu5MlVcgWAVZyi1SZAJOFzOsMeReT3Fi9m9JrYe0oH9pb6S1l8JLNm9vKrWjWIl/XHNRGE
Ky6rS3t62A7BGHzSAwIgrgn+ygSCRtrQqYdvkGT+X4sn0Qwd0JnytN345Nr+KLzqHSZR1KeChNxq
DywFBvQ/8rHomzC5nReNSMFgKiEgHV/c3FL2Ts8wPBWbEL62X7ONBeA/RHkcYPXWQcgHYPvq/JQt
YlKmkr89b73fPf5UbJfcVf2Sdkl9gu6Vg/6gZUyZws5swQsAqqoogiEqvHB3IKgetR5VQ1hZYEWP
rtVg1F0zmPbAPedlSHtBwxqRhJHy3vDm3LIbobAQGaHc26MsXyp0Rfje+YQBHun01oGWmv1COqVP
VKbJMsF7MY5YTNVLFeQYhzJ4JbUwceSeXei31YZ2wv1PL93FupIaDxLjPyzOA3t5gtaJYdE8WDgW
6ywl+Xt/s7OsbCk4WDOntBjKcq8fhKOiJJKYkJe7Mk8yGEtKheanwgH/VUE+5YDfL0uIbgj1VK95
E7MgH6OKFUtHQU0gVzPjyiA3+bH4BWLC2rIucbxShCTXv+mqVwlquWGpk0f5kiUD6CQHGUOmwScf
vZ65EWEs2hElZlwTPxs34lfgTpu6xuQehQuXTTqbRiCBi2vl0EATHXNh1eGkER9kwKHzHxfzrDp3
UGbqnyd9lVCkztcWG7k0+C/8Pb3o4bdW9x4lkHL/ZIQtlOiNOTishYKOQ3kHinyufQJZhCdnSD+5
KLwieeQRbYv5di2GWcSBiXWXsL57PD9i1UNkgS2jdlm3OKkyuIk4IJ6sz4q0rDIGcSgwGEB8p1Li
QTGuvBFBltcu/tyv14TV3MNAASA4m2ZxaiOqgFL/oQHMeCLjWSLsjcE2r5CvpuHhebWo/T23LJgH
uNao4eLNsjw7Umjjpin9hmuFpAM+40gmbAYFCze5e2niU6ckVq+Bqj6hNhR4Xx5PPGNSuslU02N7
WrqHcRKQfjwPyoh+LQRXjrJOskMdcVM4xFvTBku9hFVaMy1tGkEGBEecbw0AgJGJYtl1a5dJA3Rn
5cFF6Dkj0sRbIyauHl0NMnEHIlVDl9Q/+C8Xh5w7wzOjZ1ftRXDQhMuXw8h6ZZpm7GwqtarwZd1J
/rG6Lfhy+4gj8Sw1I8qEQTukhH61OroCutNxrp00Cl+/HsjNu5B84GqyzYnxj7OwU8RP5xdn6lWG
WsxJDfSpqjaSMGKR9aENdneKBK4iHVpuo2MIh2Ubp3xXnrYQsurta1QjcUK9ehl6HHymGYy1OzPR
Fh+O9f1pPe19qHnsKb/9zPaZr2TdBxoGWW4ffT0nPH+69siYc0s/zr5d9rRudRPsQn/FBL1Ild/c
YOraGtA/ExMhkx0eTefLFAk4RzzS6PQHJ+F/+NkP2c+byiF3c6Xx/aI5TU4nuyPVKoVKzEGG91gR
NB4NpD+2soppWp/9sVtXpnVeel4MsGwk38Cs0Mb2mP/4N7VAKAe+h2fGeXv1llp4svVAd/hjrTyg
iRKaHKOqyhjhfBxhbB/tYfQoylWsl2z5fM+tzXF6pqYXlEY1j8wD1fF36Z66sja+Kv+3ghwBtExR
FavZbATWkwfrx5ASlEt8Fah7DdP8pUoElkzaZsEqDFylbwh0qId3dw4E3BnqLe/c0R0Kc6xLX+U9
BsqlawwEY7sL3+cb0aJ3A4NWOI57Vq7DcVzEotPoWXwaCd3r+PTm7id6lTS20SdkJP4pK4tJOiq5
I2Vw+rkxpB6GOYqJO9Ty/rdianioSGe/nnerybaOr/91Q48t+WXdk28b+qpseSUy9IddP9NvtxtF
LevwXRbrHuk2RKYQesT/8nKFa6zLS16QijXE1vb/MQyCfI35RBjdQFkWXdAECJx2mTUYxX5L7geS
8FLVA9/yKB3sZLPi+izY93K8txYi9PDTDMbjbOPDjTISR1OlEcLesY33VVUcMAWZv93ENJ1D68VS
aLdyJ1LDBSF0lRb2SGc0pTXeFgo/GrNWvy4A9B6/2Ll8j6tgtav55smHF0YF/mT81YM6P4cw0/Fa
sfqgAnPdA8Yz2QX1hGAcPF+ZRNQssE3yp7YLhK5uvuEoe59CjBqic0HsNi000q64VGf81Dik5tLy
f64gzqF9O5M1XxamR+UYCT0VB5rpoDx1FKgY4LaHmCPR5MWxhgtCNUPX6j6BRcfNGElPLv7gWzPR
jW17NGbCtT6HDucIjQtjBn4sqVfCv2iCb3Jh1IynV0EwILRmhOYLx0FccIN8JPOTkELXZpo1QNZD
hb2TiKdUtILgMQdj/LRHoBtZxaM8tEgqtSCcFpX5o/JDyK68SB6zN4N8Cs+qQHZY1UEvwXoEudcC
R55Y+wI80DjFKiK9NuJkDP6IGvWRetAY4PcicMitRb3Mp97AUXEEvFHZBDWcPbDN1+pYpStKx6Ls
Ww8stXR+LyrjgZ+4zyaOLc+sw9cC+kbMv2zRReomotbdfu3HzjPw0aqiHvifBphQtrTe6j3F55kt
lSmb9tsZTfZpmzSdATiniJSG8d/x2jEBfRoO3GdbTmYOhcuQq3LGslKOCHiO9gKeVcJwCPx47P5z
kexeVSN2JtWBALrjLtn+7RIX4ckecoSIVN+iSshDq6R2hvQevX8CnDUfJQqM/wEtr/PG0MzdFshR
6kVNOGdDljLbAVIpgLvKzUVGHT8XoqFvDUd7tnTFeMDJc/Wq05nut72HRpg5dwoqg6Y3az3z7Clp
IYU41qPX9F0RtgI614c4r94pxGOGFKEKvfhs4Lew7iPrvZS5AM79edIigGY+jXYLhU/GgNidIkLr
w20+KDOwCPfqVY6WI9gebjxq9gint0Qy41SS4N2LoYiptLhYOo9IHpJsam8yoOfWSKehZOLzEjJf
0/pA1nIiNnop5/urIFwM8QLLc9ldgjnHfPD02LoNevzK8KKpu0YXFJbZMGgRMOfvhw1bUFzgN/XT
AcEkUPJJA1hg9xpBHAJ+6pZVwjM2oAHS3pYyGlTEXIBHyV/NgjP9XvJJexMCw5UalBS0cunigw62
1IwTVaNtrMN6nW9wNMTr2a889rE5R+/YuS535tL2xAQ8JtDb3iF6RKM+s4uabVk8k30Z5brN271z
dPEWG4wSYVdjDyNsCD3dwpIhu4InYOgcVY655MFeCh5BwBGCbQpuK4tW984gRzunfdzmJTDFFytZ
V3uHPvhY3eBB8n+Pq5sRjBNrsc7WY9LsE/7LvVG8klb15XNSmofENPdnEXr9LYwoKvCDAK7hOxuX
TSAvIDmhGnc0fREhMtDrj3dCy6qKLIdm8RM1a+QYR/ZCn94kncSCGbZSaco69/GBYujMPzWYBqwU
ZfWGBYhWUBNKgQgyt47lulqtnAcXHhArfgMmih8+DD/gXw5v/BnmXnDoYupL4KJ+QczDrecUJ+5u
iQKvRLq+IdY6BU0W42iC7g0/4PxBWw30TGSGlnjefY41DdxBac3GObwJHEN1fBq/wtiJjE9rAcSt
NBtRj+4erjM92zNAfGAlBo8M4i1MlEXJatHA178U4lkFyTsO8LsXgFLrpbEG/DaAIeHTNQnr2wG1
aV8QBhZi81cYYxvE565eLJCBX+984spYo9FJMHTlJYiEYrpusWFDwdpquTxb/e2N2oxgZLRQzzX8
HlJYzEjRxUfpEaGPd/TAtOEAshRf25oMe/k6f3k7ANH2RoqDE2dXM3FT1MqLtjky/sEKW/PTkk5H
90hVsGFyKWa+k8XAcKW3dWYJXgjegHswQHEY0Ih79QnvW2v+BrVQMQNQbuBUauICSK0AHHITtZXm
Qc0OOiodKoKM4iO2OCqv1YyCeYPJqFKc0v8L4LUZ2jpFZz9Wy/HFYYTp96XGHhlbKQz6OFaz/qqM
y0LO0z+87DTrjEWDIUIs5UxlBuXVvfbFZXjRPbiLoIf4v3MXBQFWkigYLBJxw7rtkFMDx3WH0s1q
idNO6ulgn6MoaZDxV7WeyyrI6i+hPDg2kkCnewCWegw9ucxcN7jrFEMyI0BfNXcydjDGRIetfV1l
ftxgMTW7AkDRBz/Y87PO8uzWdmPAcDI0WzX1Qq3TvhDK7NR5DjPSYaRuLXqc2291bHx5IX2GTxBS
bYokTuNOg/GWOf/M8YbV2gqetqNTHlxthv0sc4pTxT4n55eZEkBJn95KMvOzU15A/bnfZRssKV2I
E0k/lBEPeFitQyW9jkTvlwS5NGVtufFt40kCUneiaNJPHjcRTI1+7eUQqhHLpQEpAQ/e6ngpfboC
u1FrlXloCN+D1uu1rJMCxHfE0Q1zz+t7SzgqnezNpCH0Nh+zBVqiAeH9H+c8c4RXDeUP7bHVhVL5
jpPbb8p5G0rNaKws3tbSxu3nssZG8khlAQ5X0aumOL902Mk5wTaSF8bxBvfbFW9awbeRqNWScANx
h9HVYVbvoJGikbZznVj1qACd/tOIS5Lkt0EaYAe7w7aGbg4bGZJCxW1qHC/YOcItGnQZdvROFWUy
2eiYrWXvGe+3AKpp9ru8obm9kiNYgtkZ2S/KLnuZxGxfdIHS2Pb5C7RTRNEQTsMu7mHHEMSfScoj
g4ZldNNhq8/A847emTxdRr4UhPzpVEzvOXXEHdP40FjJWi8O5AeAkFZJrkSqJqj299I8OhAyqA/9
MwXQYUu35R++PK1q3tHCX0PrVSEZf9u84HF4mgmai3r6SXPcI90n/9acy1gee6Ql+qj9cfQ8qhx7
s0kwKZdEHm5PR3LyNYJDVp+ZA8IgOUwhO0Eq56iZq09pLyW39M80KtgcpeoD5Erni6ruZAWq/HVm
bJ4sXhT3fPNih6+kKPBWR0ML+tor2RmWFn7BIBMTOrNl1qNRWebFgh0+GNL4roDDxUB4wZrKXmXC
Jay/DyqGlFhd/8Ujf8wg0Lcb+luJr9YAiFmpemCijtotO6uPKulLsmRG/Zj0WrfLaJ07wUwt6p1X
Kyphgk3w7XIOrqMAVD405xdmQJR7ryZUApJlm2Yvb4j+BqQX/b6W3svTTM8eyEPQpYJ32zHhZsSa
T+saSCPkApaka52SkKtfHfgA9kun+RtttEm0JmEf9D/c4fRZU/8rfJL0aiQgPBw+6u4mkrg179cF
Bfi1Squ57tF/IcKhAOhRLLJQv/dAmP/Afq2S04RWH+aMdtHahLzo9+FqzP8q3UsZGLSuitdZTyc+
dJT4e3REHzV54Opx7TExMI9LnZAxQ0DCvBnSlc72CYfdbZmQvuFUyoGdSOA/c8cFxIYVRzFpU/hh
dngvCgKOYBzUEbXAC1Vi4rio6YSNErF+vBadoyG/wK8EWmsSAfL9a0/hQI6ryuKGon06QUx8eYQX
3QEbJy4lkVe1JjrQCYs+85DS8H4rpJddaXMkdfwdYorvU+lTOY1WGSnt49E2zr2Nb9ddyX5w4YM1
EaYtO+OOBixjYjferIPG67aqZJFtppM229kGzk6eXQ3AL2nSD9r8JLLKYA62mAqszxadHDko9pIj
JkMKv5vYh7LmflZcRO9EkWQvdLA8yI/qhcX61UzlgPbE1AN0OPhc0S/Np9r8Ez0BdPp5gdolbZib
cg54dblM1EJf4PbrXkTNOQDYFLpSSNuuAwL5r6EMfr4BMl4QWyuIIOjPQyxc1lhoSI07/phulOzP
108fZ4WEQ3L2YBsIonfJl6rlsb45V+JJdBPMRi3yaCc6W/b59QM3DLeoNEOCjuX6+jNbj3zC74Nw
FcdwxmQ1VqofZcEAk7jsq54ek4IVid+c+pn1RVhV7cwiMYaPYQvUF0VUk+Cmhv5vx8n1IFogbYQd
1BfLvaNIaTOghJECPLI8ily/hJmi58TjgJY8YNXGi5+hFQPLbILVggMBeLd6PlExwjMt8v6XbOFC
d+h3ogCaSrW2Cbw2jsU33NO/8m25+5/rCIbcn76FfeuM/NOt4oBfRLvzpms8YVAmaQDJDgIcMQnM
e4GeZSstawNv3232jRs9+ujWb+al52OSgg1gU1CgIGEEc69QfdZ3XK4YBpeTULtazGJo6QtKHYK7
HlGRp+G570edUOY4kGkcQk08CHMoRAv53+5A7Er5rNFecFUPKIuIjluDn/bNziQlfTnthvAfIfbr
lb/R6YQb/Qaeo2yw4l0cEQ8WmkuiSpVVaL4uIU6T3hizx29B/Yl/FTa5pUJXN7natnMYM55xny3c
Kq2FLWZs3Q2dZOhH4LF0px2Xt1Jq6eoJBlSXRM+nVu1FeQgG+Eq2rE98Kdv9K7n1pZq8811ttNsY
1lAPCT8ErAtvjAaNQrjE3jB+C5T/Z+j6sVE8K9ZFm5wp0oy9sn1QwOPQerorsErtuiCDLR6t41jR
r4hVaTx4ujw/9EP5zBwL1HojWnfZivAzkB22Pf4iA969lPWOpTe7PeNdusTYN19Z8qhSehLwNdFu
D5CDjuQgaMXdtZDs1xG4dbXlqSW7fDspCchmxAL7MpSTQ92pcP/OyHNDZ8G7XJTp7bXmWTWRVKFm
aUVfN9B6ptai9wK7KM3yhCJDUEcbhmi0PIlA3xoZjWHHLvqpr6ZPBeyAIKLw7j7pq5w1olIOh7qA
qsaofF+jvdTFS4JspEHqVtrV4XnP/kLLI5kdyg8dyHfpho94zIp1bHGK4cehOWIHDIrBvaBKb20+
agkbhyNB34BVaDWcAtlf3uj/8nhVZ9r47bHdRdbZaJh0vRe8eqLZa7GiI4uT72vuUbgWB5QmAfp9
6QJu7jFxqE6xdJcF9FVjgbyfRfFa3iUO82Z7sXy2fNUik3cYmyzNpnLdtQtZaAr2JscB3qOkaxmD
3zfL4F9kGyWT3VgJY/NOHPuCLwdMH57uG8TLA0/9lQSRU7Km2lRb3FBvs3gI/2BGzskRF+ElULnW
WxZVOBDOm3Dck8jjQmA9wlXbYN9xIUXSJh76XN+rSFmdN+/zKqOg89Ap3ARoVZjxY28c2jXbXEBC
FDQ3hDg5pohG+NtIqoboCDx2sQnlQT8VVI3Q3FUDUK+a53llJeNG7edDjkqM7yunVMD8ChH3wFc1
aPQDlsfty7z20frM9Yy2+gb+tNSpZ54rxqYk+ejzSh9yIQ1gFzjAkMZmmI2157uby3RXVprV9U1Q
By+QQR50Wvo2duRwZZXo8eAIDkcHLLSZmtjH2R04rsf5QKSAR30xK3FdAv8bVI3FVnHwQ9kIS+82
4eJ7wRKvNGr0ejFeopHNoLyQ8W35qdMOHODC2Rhvrlia9pENg35oh9ivSF37zzNmnkz+eYeNEMQv
2Z+1otI7oA0un96+moFBT4ssJEeH/BBnG6AxjlwxSy3KHSVrr028fWMfG2uvShHcRcgTeeZFXR/Q
RELmCMIVVF4YsBYH/Rm4jbFRlLMEDjKSymGpWwxDIxc060AprQ2lb/EEirCFUgJqjakZSxuaDREq
Ft5ZssOuEem329za0dzseUQHa/c2HEDjSO+ucUYHpMfiDmmsawTU9y7xBI+ZsGsxvrIrRBzga+13
cLW3rCWEJCiSGuA0ieYT3u+3snHRVhfG4YNcM238xKmCl0MYSirNbQIbq38h1imFbuFL7SLdq994
WnyzIRYDCoPqu/qUOtS6LCEJf5VfLlBs2m5EajM9fHOeK7S2JpDFnFdqDhZnh4sGiVKXz9yLk6lJ
37stD0WqiecrrYQvyAVcSagsA0S5uQLKhSv7p/qV2PZa9T5vUL3NnjUlZ0DNtxa0QR1pxWUpO4E5
S51j/uw2DGYmhygo2/tWoGcZNWBMJrFbBQR7tOYGUDC3gCsJYbwRiYcNYscDBiDAGPxiu8gLV54p
PS/ah1RxKByS0OJfySsOHZkr5Rbdvy0bXtO75UCNCV7eMOBmGIFtIjB28VE9f+rPdH0bxG8RGWo6
SIG4HgYSfeI2/Yh3g25IZgPFDYzYJ+k/LACf+yB86spN7S0fDfK9+Fms8LCgBzyX+qWvslbE81kl
kOkZBn90iRVm1XPmuZDFHqOsrFHx0DlQGSPnOyp5IzaYvlBwHJwTCW638StUAd7CykpM78XKxJH0
i7vS9ZIedwsbw/zeLZc6yYGRCHXto6u5y25Gw/V+K1w4X6BY+aKycN60EyP5GYT4DvGDq4lHcG64
1H0PcaNujEofnZ81goBeo8szRFF7fuWE9IBh/xs42o+EBME0/XnRB4BJVLgEEKDxNrdsdZHp7D/q
CGd8K66NT/Qx1flxLa4gEZOgxCiqU4uP1JIJlFLhTWK24/YxWamWyFxPRfJsYdfrKSN/q9bnDxve
oR5I6QL8GsiPA6PxXn9Gk/U0yaGQmF+9SOH2SjRQn9rQAGvegkCILXEBIzF8ggAx9ig9+Pj5mfBe
O8GMvYQuubsR57ksEVJOXdmSoe4FjFrJsTutctG8/BcvV8xWQHwG0bQ5yVYgZzd5BzjAUNa6/VdG
8jVSNWwEChK/53CENYKOKp638gDGGrqaeb71SklkirT2iQnrIddv9U/uHHGde275pHGO4e7Wsj2K
40Q8DddtGobRfBkWKb9ftILyHk6lZDhjuy6qwbyAv7BuRtqtq1l1KsRXwHqSDOZuOWTU966DZ8Co
c4jjPqLZvrYrE4uo552SP+SiC1Td5LwCZn+8P0EKOHEl04GboE/H2BjPiFxw90whR68UrOpUNmve
wPUjcuIZi2Q6K/Uxz3c2j7V1vINGHqy4fhgY6cl7pRq7MaqPl9fxoeB6KtMTCGvu4rG7HffIp7Lk
2k3eTT7B35vGGFshLas37K7kJm1kbGYERQVisAh4U+cxctU/8CZsFNXvCJMST70wbGGmHMNlD+tn
aVJIwAwCga60iHudLcn5vAuAIEvEOXSOh+6Zqbywlbi5zov8vmqOW/UizEj8cW74UanAoV17uP4f
Hc4JvWS9lcEstYmYGuI333AP86bxFlOitugJtCSwg/T9/ffu/PtcU3N7kLAwqpVjdRhByN1K6OP9
JwAy3eNJzTjLAu9gFEcVDpVxSIl+Mmh5TqlLQh6k5e+VAEK+/O73PY7g0J+9Uj9JoqXZ0m8H0Uhv
ZzrMImri39TsXftC3xYBb2Jmy6AA7otlD1ks9pT56R7lIA/H14B8vPk+t04Uj2mWelxQkJY6Pysu
kH0HstSoC7k+gVRCN2klZQ/JkG24xXhb/H/eK5ppik6IaXPKwFwyfJb+NiVAfeGeSx42aFA+ID5a
4rJB5DKXJcAjMblZxjooi2a8cCiyZYwSQzPDuEMD/UXkKFZ03jRcfJwxNk1lcfHz9wKmO/+kJlrP
H/rpLqNT/UKrBVyAxu+9cPQ0uaPNqe9QS/4kBk2GxeRZ2xfTsdKB8gDscQbgVy0W1mWUlyeSUQHe
tYda9Xx605x3d8q2Cd4vcp+8O88ie5soci9X7LWpEEs3/NVbtnFVp4Bp//ScW9YCLAkAwPco7BUt
pRzX/A+Mk7hbEynTI2tXmBNWtBeDmoGXudiRvAJlBZdMzYEh9htV2rb2jxmbZCQ7B1shoaCpBFmU
SW3edcgOMCZ5O1O90qUNKOkYSzL9Q7v0mMTlrhoF/VjUM68hcJx9jvm+Wsmsk2NuwhI2upppRCIn
KTFxBQIxzUEG2UHVp8ZwcyVR0fD2QmOIdSvrIXBOVD5dXpxAgdU9PSGOGEEMQbT701XGcm137Zq9
91Lum7QMJKqlDK3Dl5qdq/IPF8lDuW4dIAImy6RwscP8DgVRNsSIP3N0zgggvXhZqNA0/S6pIme+
sQ4kseeFWowI1PenmC9aU8VKyXYnUQTTKLRrbnL97dQmwmGsfK05+JfqH/BU1Lxig9MDlVe/MVhi
YY+Y+EeLeYgylbjv/iCIQjlE3Ya7oj6KE3s0YpmJdL0hTKveIWG6On6mbU9SDVIX5F2Ed7ZqvnZY
+qu9+F0Ajpi4mmhUreTWCV8rNZZuPCRrPs9Ax2htihhLTTlSjY67mw/mnIzQ+/g0oqYD3/EZrhgh
ib9ZWJiNKrgwgSVHFWf5WderdJMxfuiSalrHTgDCSqbAOJQLaWNOmRczJZjbmlSop6cwbdPF9NhU
Tm7FkVqXc16op4kp0kSUB1kU+R9HClFGTkWjM+ioX3eVcOrFKcCMW3CNAx/PtvhR6SauzZBCfW6Y
MWWb8IRJvWuIZH749Djxnd2wNHmNZiKKH+KUb4TN0jR2/85AOZbJc9rrw8JMi6AQvfId2C4s78KN
srqsHhcTLWHb4szOV0QLS463BDxs3LxVOEb2QYn4KLeZeGvNYXixuZFxKzGwfu9uFDN6QY7+oWIo
akR5eJOZN4GidUVZQ6bmsaLdsyR5bI9fLWc17RuuYKTOzPe5z0GJwGQRJp8A/HVoMl34vQ7ggq3c
HrpyBmGc2fDLIM4FM0180s5/Lnb3tx+ZaKmsphhn3idi+WSg45plc/di0G/PvLhWyBSIk+weixNY
aMZcc0Vd7GZvVzWySlPk6PvukCj4N9SDRwp2zGu+Ok1hRT/E5RebcsYqMFqp4BrKeW4pZUk9wovG
rwivOPr3kacOsVc1gBywyKMzBlbwc+hKPVDPb0DgJvtfmo96adNksjQftO2rG2QfE2QqZDZvwVy4
mZ/brsgq5k4iFrUue3UtIa2e7rE0hVap3Md0MutCDir5CLNmJxYeGV9T5EHvj9PYDiJNVFR8ceYR
9GutKjMf+Nb1NLKON8BuUstXO0j/GAL/5INwb7Cpl5ewDNnPTb+DPRLpNqN95FPU1n7Xtn6978qh
LtHEzZC3qdJ63IJ/uOK6n2wbhgi04BxOMYoHbKTGImSHzzg1dqvL6uiGRocyt+Pvc4l9/UDReY+L
v1v8V/ph7SksQOTxl64/Jo9B0bJrd+zybdikwKRQjWXhxB8Uqyxpk26bFfpuwSbbfu7W9wggTekY
rPgJrJ76Cvo2EQ3xUSjkdq9sPXeJjHTDqxPpBeKx26rQ0fhckG1Rmv/KFipFKNnm0qynbMPNdtD8
dsJrHzL+yZXCln9Bpm4rko4jpLhrYXPGhPhF15vFyHhYeWYR67oyuOVgYnzO7F6BYNnQMiZFopFI
MWaaU2Tbh7i/wE2wHtCN6cROvlCrFaHG151pnOjUZa9q0AnZTxFUODuf2H64nHnZlr1Goc6Dbg4N
eo3ngnamGxNTrZpnN6XRLDSxgmy6QTfrO4Stt5LxR0aIs4+fD9tXGOtJRSpcWiqLAQ7QHTngrmU+
o9pn+vbZ1xHza8OJp/wTNteLDwrrHE6qAA6KeuYbid/8Tv0PCUQvpgM3rgwQbnxG1L8g91Kxogc7
uUg3FMRK9KD7f+lqMIRKUEphPnO7f4mcwcdA/DNs3MxdPdzmkqOCZiil7/px3u14ZBvoaIO6p8bS
tOTqY5qcx+YG44HBKSpyURn5j0iI88aY1xZaT2KQGClzLXJKd4Vqd9gbLpYebrLztRGVs1aXbGk4
XCRjTzgvI0XEDkTDJRtt5DZlmTCFZ8Hp1JyU69jTmQ7KHZoQtCbfYCbmUkRQdG0iAghndPpoFg+E
sDgoZegLfXVHxFPURBxX5trmTBLFXzdqqRHrHUxDv/Ix7yzSRSIhAawNn+4l2mKpmhf2S0MmsPYC
3UmEpCC5yIfqRwUJm0YpMR2O7KH3g1uAhqX46mcjGJb04paacrD57s4xtoxliuun3IlNqq82V4zn
9r+RWGtZBcR8UxtYQQAaE6WAxrssP7V1wf3EsPgnZ/uCvzKoCAHvkhmDcYfZVqHbSB8r6Qsa167q
iqpxFQRLD+1vaMMGO1C0OYTWSuDxF3EbeQiaAI1CJpmJFR5RAWe5MWeKTu5uUSVgszYdaQV8kiQA
r/cLSASKNNP6gt6T1++4UHoDkoGovmNVzbNQ0YMtyufOnZdN6/+8AAGukY7VoDuNTUj/HvmwopL1
CvXh8uMsFJT30O6CNypEWLSFdBWtVSxg3xOiWuv2TyGzOKpN66wgMkMSNjI452XCxzCKWPVdJxax
ViRmkNxJV2TLglfjQcCIVBUDj2gRuJXa0tpeTcKI+ru+PP0ShjiR6Z1KpiIe21++JHjxeZMNukTF
mGghys2d9MdplVbabKSuM0ZF4SwVIYgbewzAba9NT8q6oPthxRkTS0pbNMfJiXCe3t/JjKQHJXoG
UYyfHu03byLQzdyBPVtZDCJcDMG3OHtNIfaX/J5LgacJurADi0+hyTj4wq6D1wQsySUnn8EpnKnc
4vLUeC825gh03WIng2vMyeaBALPBkz2+jxoXMX/tF1b8+8oBSZDWZr5j8zj+ATn4VZ5IHCKbCc3E
CgmG/BA7zFsGf5YBx/z23eZCn3jIQFD7CphUI/Vi3HvL5UX/PA8Y1ot/1TaUDzktou3X9VgKCRLZ
DmdSHJq804GjKHNcQP+Hrd5acXIfkteXbmTLajoQ3lSqpfyP6UupwipnGvgHO9QQs1neSmZQr5Xz
fQ4oTNTR1u3OtDzeADfJFmWpxEmRuVOD1yFmGBpmUHpQj7bM8sY4sCrM62JYnMqwZoW3q4OOdvPL
FRml2q12SdubmEK9K4dTK1emvfabxb07jiZydiAxvvAkBom43ge/glYN2Fii1wz6tQJCBp7q0fT+
P0TD0zivcpYNnrSBE1++XYEEFLiu+oCNhP+pE53X999rEqDlgsn4QSInb4n55ADa0itjxVxCivOu
IGf5Zu0npLoKchwM60JOR1lF9V3wvgbxmeflrPydzWYIleQIHxvPvcldYmF4yJaET30GZVyF6y/U
EBJQD59wmEC9z5WyXKk411+a4u6E7IEmExs7NNI6NyimBypJVhdkgOEHcelSPAiiNiUJCrSCMj9c
Cxxa8mLKyaCfGbU1/WLJkH1Os2d73xhqnCWbkAsZHGhJChvzADPVkulztxXWdMZxbRgksReH73El
9qkXTWOwbaS7C4dZuzkaoQj9XYrsNY1xPCy90JBaQz6+snm0uRee0/0oEA1e869JL4kX4Cm4lEPR
XF3X0nP+axxnJf01bUMGpicdFNPkrR2XabKNVjDj5y9ScBgtNaOICU5SuMBQ901zUfwjPvCNWo4Y
Q42qfJZe0hm/f0nxRVJ0qjC/EIvI/YsnD6ITnlEbIinTSGtLu7NFK9LI7W541hBt6DwVnlkSBDsn
0RAnWaCAwwcNsR5PIGC4zKWt1fSlP6LTfNXnQx0I9Q4nrbVW+1DR/4JZ///nmV5sh05W//vtQUhQ
uli2BeXUu8eAU4R+Q0HXGrVO4rewG/aDWDl//sswDFUZ3U1uDiDDQkBwLcECLORQX9IRBuQEf+um
/dcYuHax8U1+Uoij97x7gOwkrV5lvTa7OvzAT4w/abOBhmZ5RxGjjb3mdXfm12J1darRXE7hBKvF
mgL44TJSG2974QQp7Hfdun0NRalEGo7PDSRlIzwbia0/p8ZGO7zLrKzrJf9qfQqQYcnGyejUhtuZ
ga3n0wksOsnWIIMLdV1sq0JmTuLfwdFkdvbjk5EGy9XUrU3qxEQYrbKIJjbseNp1VcJ/c2LW9EQu
AEGB62Sm0mnrzw9R3QU5VUMhzkneuTrNFDm+nSd65uBfKk5bvJBKvmJxD6kYW6rKqV+r5MmDqmu3
8OdMDyJ8mDmlz6YPAh/iQqZn20TYFekV2prbcI5jim/vp/Vris8zad5i5H0hgWyelpqo7Bo1/d+j
eXRLn04yiy6jJsyo5nyNxMo+ZW4wRWqIPSfPORNrf1/XVgDSaPQHm9At96THOn7sKegP8yVWNlua
9Fn41msnnelHaYGwiaWCfcRLeVCenGhZnuYdr1JSyCsjGW35tmiY+2Y7YUmvQJihmUzAr8/VPYr1
Poi21O3yZbCmMU5vfkR6pdZ1RXppGOQVv0xPfXpHPC3kfGga/iPvikQdp5yiJzoeVvtupcRo477/
R56mkUhMnXeporZ6C91xkYvZ7KVbc2EZiWW++qZDAfCY2PPzZJ4oniGRJPibsAUiMZmmasfMtnm8
xCwb2szkvelwHQjYN7r05Y04kuPN2rHDygF3AdsZ8jgEOWESaW8horG66vjhFuABTveEnZOgryeo
TpjXqzVZWX8hnEaT2xmNV5xvqTy76ix1t5vMPqDtYnMQxcaRJpW/KiI/gGuaY7p5Utts+rYTIACu
wfGXSFtELWHhJVBJQbSYQhoXnUQdijHvAU9NynleAck3FMpREAWd1wD3Pf66qL9GmsR0OYscNt34
TVbAy5wqC+9NCf4XPev05uHOjGfbDg1PH5U3pIGu8KwVseaACaR6nZqPrX8kJ8H3HAXtMqoeGTLZ
gghMSHCZJlWY0aQ+daa1z7hoWqS2j6dwZgYkPfTWK6uQChZN5CXtJDxzr/At0c14KMsihWqYraCy
oh9J9tpsg6QSfrXQ/Pzapsz/JMuHZWLZvzA6fslDGTT+C0dpmgrJSFOf+BCaVkxou5VShm/psjpe
+BU3RRrIl9ttl2T0Usiod69bsBuITMmkqyCnr4oOOUQIf/f26SoAsQOI6X9d4L7WNflOQ+GXEHHX
OJhaxd/hp4BJMsnkimw01uz6raV4DN950bOVCx6z3UX2dBBXCq8cOhmivRzptV9/t0sbWjoY+EiW
XL1rV6TDURwv72kkDPF2IKfBNc3kkUDeJ6ao7huLs7S14BciWJLTa5MwyidHgvjMVxLrpqhNd51x
/c2b8UmSa8l5GvVnKrj3CQ7NdVGYbe+29TLlOsZauFRay+S+dGlCvyp2MufZb2ACl8pTirTJRO3z
f5XOYIi0Ub5x3wgdjvIWK32bt91TrfmSDpl+HWJjLPXHS6VAyPoEzStXpXV12DrnxCnTWLsLCRf5
Rk15XmmMahmVksYs9rMMzvC9ZJwT1w808D0VztcmfPmmrENH8RTx1Gj4GmxFZ/vXnXE0PIUaaXbh
5EhpOjjYrmUniIixaJw++dKYLlc7mrq0x3vEvml7ubxDjl5wCIyP5KFCh5CEGfPxwFSpKqYu8lmv
9ykWjXrzw3TK10RKU+1+YEDwku/OrfbqVFnlJRI5faRH0JJcX+PqAcRxDAZhfU713YNTg676RRYv
/pItb3dgkMHOnfrgN3i1V9mFn8cpbHqtlHoTuRn9+sJz+WGsMargMWYGrmdXZ9Oqt85II2Gai3aV
7+gYs8xbslmJN2LClN6BmQSrpKMdpk+1Pv+lH6IPXHFDqzDGxFSKDc0+5ra7V5XgMvC8ErduVoaH
V2d+FEH7ckxVYkIel3KjYvONeaokwmzxxYxBvjOnqBn5mVyLr9Mn3DpY6FIIG7Ojqve9/gCUmP33
OjndRiXmECrETrCPrr+o18gTi9NHI2wdPqprhSyhnNq3B4ayozbWAFwYhfSpxfJ81q/Bq1BVVuGV
pHcvdhCufQiaAg5rkxE94qCSd5WuZmBObzsjNHFV4GWINJa/lvgt/+ybhKftdiEtzOum1UD/B9Vg
a31JL3TfwKe2lz9ICojPNQrgJil0riRVO+Dh9cDRXvIrWy/a/6gNpgghzq7ZdroYyeKL6jwCTmEH
53ycIb26Qg8kD3yIoLnxxJCcut41e2Rznj/s16LcAaM5lYe6nAwYlZF+MUAAopl0KH74lT1dp8l5
Va5u9MNDZq1l4IAxtGXgmbythxx2fkL8HGLPsKaFBmbL8qPAV8q9V9aLZe2gNYzaCNOX3GaEzHKs
ZVca8gPjDua4egi2pG1BMv/bn+spnBoxN4JBM1n78f5UreYVc9B9BXRoGB3dFMulFz9xdo7SOR6k
PUNL4Jj4Oqsl2pbFAYWF2GDwP5ZCkK2VGiSjH+KBWNaZd6cGDb+hD0wEfo4z3z//FKToH0GMzsTY
Q7wvEHForYALECSMedJRKUUMC2vxkdjJuCXAImNzDymoa+69dtoSSGhWYVO6fuuG5Z2Ah++5ufbD
rDbxcI8SVRkZRVljBnKTKSEFOiD8rrZ16c92gKu6tNYjzF8ufRCm6xcX0Qu4cuV8h0SxEvOMWYrS
COvDFSqTdQQnIFNZ1egkke9N3G7GoCzteXPIyAagu+u3f7iY4lI0kE7O7FSbB9+N9jh05zCDqhSi
McNF6Rc7tgdcMdMBQG5t9pTdZ6MKj43U+/o6c6ZoEz1U8Widh6HA9dd548Cg6xg11tuAnuHwDJIF
306auwvl1xPflq0xavXJ1CFTNwMZZJtN/tEKZSqhTQvOh26EWT3mM5m+ciIweXsW6D3Zs3Tkfbyk
4EIwLHfvsPp2SrFRkM9zUfYGYa/NzFJ54og/zUto7uNZQuYeEk/5dBCPtt1wvXFwU6bEEz3z8kUO
1XNfge3VnjvVrK5frYj+THC+50Af2xaiPx/1Kafxh44yBq53oDS9gsGbVzweIrKIWI+s9cMnQlQ8
WBAMgOzYpKTS3uzQ7trOPX29IPbevDWVVouePXJeZdld9W3fYuu/dfM9/ggsN3CtJp9Vy0HzmyA7
4l4qUI1zptu6xG18rEPH/uMZc0nxKqZEWeyDHdTV86GfE0pwf8GVNGCSdPoYRm8q2okXU/w9A/6d
EFFSKQvRpIW+Wp9CTyvQDx+0hfGoWUlF93NCZ24BNgksyk+qB/EhE+84G4XkBrOak9o+5j+7CkHM
9MdDTlcepN5XfST8hXWpcEXVySl8Gt3VZum2oBwSnm+IzRcB8M3+bHrzu1CSjCtFIPAfnM8Sox5c
9qKDMcaZIv59NMsNvIC7JOivUQJjtpsZGcQPovb17WGA1wmUMusarG3MwHFinX+UW55JvsABIDXG
G1DtTQlGhYIFEc/Keq98gu4y46vqwvjgRijKExyVIfvhS7ouszAvdqBR0NLAFaqq9lgmVxm+aTpZ
JqJzFbGkqwSJL2UZB37bLb3OM56F4FS9zrCSh0NkKTFhFiP7FLZ//YNVvjTMONJWzzC+GbiQ/nhz
rlFHmQeeyVjnrSOs3LwIXj1h98cQYS3ngS/j5zeELge/XUX1AOraO8j4tOwMc+yf2cfmEj6LWLeA
/Y2aDTzlzr2sBCUAaaKhBrob3+ynfFLQmeMHfxvt5eKBaM0Y0Cx4UJmsZvfztOYCGDlxUeeqICYv
dFO0meBJh2d6hgBA4FpxtRIJXazT+sD+RqxLCqIcaQ+C3fd37e4grptgxMzsyep8TRCzB3Ckyirl
elAqrc51Td9MOHDyIpDqGrXO3QIDqL8iQ7ssfiPMzsk1kGNGEOYq2ImZ5/r/Kii7Idws0MqELdE9
dkbuPmJ/d5Vdy0V8S8mpH8BcmuJSdHPbIZ0Ch9n96tOy6vr8q/gVLP6cd4hWRwLAZknJvEgoenbQ
1La9B4fq8Dw+wvFnc1NJZuYmJkVmzoYjLKumE9Au6D2Z8v9XPIbpt3lgf9SfMFAfKZ9osfpJIeFE
HVY02a3CYyUjqV/soLoFLz8xqffikWOM9Hz1TWsYJM7VFv4FlVTAKLUxEhe0g0Yg20690kDEiWwS
8RnLPfmiKrc4BpAGx3/ecZzYVcgkOMM7EWdRonmiScFBT6TS4ZxwZt/lzu4X52J8QAHRr6L+tfiV
A+aizoR3EpMnAabmZC7nwrrZF0IiXxAxemSXae8+Q3ZGtx9V4YA4yzjjOjPBe/rPrjcgY7v+iOqS
F0hT3I+ssdWJWX1/foAHcd2FWnbuSp2nKpORnx/7BIkJtWjE2QICzz5SDRzri9wKieQS5gtp+/uo
XiIELljwTQ3QySoiIRzRmU0BPahNBGlQKUXsxzGZxH2IfDIs5eIt19ibH7+fEvfbniSDzfAGv4AL
8rXBl+Fek7r1cln+vHRGczzErFP4ZjHCujlOvb+DifOG7A1qc1qEj+tgghq73Y6BfVsMNlRJhj0c
X1MwNJzW/GLHasWIqOLi2GRn9kHY/XOTkGZDCIahtwv+RGhujC2gP11ueboFYPc6qFNoEx31lxbA
9Pnvby8N4xx1HG4RxVQpjLJIIT0fFbQjrmHlo7KM6365I6VUfkjv/xLglZN0AEqdotOsTbH0CSV1
y8TkVwNpJQ5R3HkiCginY3N/7dRvlKapnR+0CRFX5xbTQz4YYenurLESLX7Odpbhflwl9TPbbkRM
6Sk4s+2DuXcXCGm+T2a1DWPHiW8to3Gfrx8amxbQ5zKeJ54ONWBVSgVgagrMLTx6hgSG4vpRuvKC
VZdauvFtXOSKFlqSFLzX4XJbyscDMLAVke9m5cK2fgqd+pBNQbhF1AzOFeYb7Dv0HydQiT2wR3pk
qjgT+mD508slRgPhSPRe+xq2nisPnIznHN4aScS/oN90iv/dYZe+s0vf1ARHBD74XhvAKiI1jejt
8chHCHCGRdFHRzJSDakUywM/1dX/43G4ZYG1jz96DWmDd0t66pph/bLu4BE2KnbDN8oNdPlcQpvH
LmNAw/XiQYEuc/SApOErpTZDpXparAicgmjJnDyhp6Aa7PuvC/iq8m202vgJyUnGkbQsKaCR5EOZ
CT+it3vd0DBN/KIixrjZGGkyRlEYjphldSP3MShw7N5gpqvFGvwuKLcklVRTLPoLU9/WQctw7WME
0drpujkjh5FtpIZacuoQhQgyAP3FIMDsbz/y3tiN6BYljHGdepX3kRXTyw7tr9y2L7BvqZtGrcvd
FQIP2HzclsKtviZ3pp5qOfzItRepVJihAQBr9y3GD8HBzMdN4OAWd6xMKIz4TCqh+KjMkxfZHfl2
m+ave1/XRWPt7mE+he4p4G9AaMb8J/7jZ6wcTDq++A/jeu11koHX53JeYzImWEu6LzX0fylSvFnc
w1tQxxz5SCKObE2Ll/Ptk+69r1X6gxYYiTtsv/N+krCZNRMm1V6PhV7xxwnTZ/P5PhG4FhPjEuZ4
vVQHkS8IKLhTBDZrRE10eaAaLl5AL1MtDTCz4KgmRFa6QKsfAYUdIYDrgm+lKMjlC73nVstBtoQb
n/sOi8AlgWyVKtez1HwWrDoA3PUMar3zW1v5hlRyugFuo4IEGX+FWu2iEDxE5B8BQqcBvzFvZ4mc
m+AlHo2ijMqzcr7vnOehVgEgOZIiNhMoqj4dkEHdhg3wog1RwP3BqdgoC0I8w/l3URB9+01KtGC8
o096mngULGSl7gCqPxgPBmuL1hRYyXFQLkuoLa6Y4XgcwfDGxpm4gmJD4G6rJOQCK+L3E5VF2QwS
zWE42kcz/9pJr9ob6dwdmewGpUhmBBLbTOriZIBxLYEuKwFGB9TR0DErfNufkVlBgONEFPWPKwSC
sXu+8uyiZAzJcTw+85lK/r2WvzAIxUq57CxpdIv2DCZYTy3UeguPaavQitkb8DoHRUTUgmuhq0Rm
eQaOHEy6Eiy/76yL5FwMnhfVtBZEfNbRnW5Y1bDYMws66JE1BEcw4ONVgI1dzMPI02iyjwXhc1FS
DYwH+L+2GZpNxguuHOFrliOKQlBsP7qX35n3aEFSSFXzHtpofNpQdX0HBACCTBHDr3KgEogeePAz
5z5GPIDTfycJvKN4V2zGr27MV+ys2m1rjev/HLlMYOewaeFs87vxMQVG+WfGbCrgulOBXUUyjoNL
xy9ivW5kFdWi9ofPoNDvCSYQU9fjktfmWwjjSn6o/UaSpja/uixP0vSHywjD7qexxfizr+G3HJ0a
lNkbK/RkSiN/vOLR1iz3TrHuEPApU/0BTXzhoAoqaml01cNKUY5jE/6t4krPZ+0s65wAB5ZqNBFq
Qu4S8jfmOh8xf7TT6k4NZh+2Zaghwd4xAJMHUmSLpTV6lOn5BWa1Zp8TzCqa4dl4EIqpYT+lI7Z+
mtwRhfBA7DF983YJ5YZdy+LsIsUZEgO21fEEqXjSn73DdbVX4h/+Ctr2WgnYUqsZw10JnKu3WXmn
F/MviUoBB8Jh1ffyfrfhijtyIKrI/tYWN5OQ7fUN9qIU4AFRCmu4bud+3+c1d40bh/BBU7NBOCOG
NNv6JlWc2xsHa57ssRNSnC+B8dYsoqxoXvUJR0/HH9an3kJcVVNBJJnJKgFNU0etXQK/T2YY9si+
CrZfY6zQhM6BAIlEiDT3/OCPA7HFttDokj09Vhj2mxQdN/O2625RbRpdaH+YaJqAteSew+L98sNY
8zGUmL67fDNLYGqaOeLqvfAYQmN+/ez06kcol/iKZpIaZUyCtYJ7CU0FlNkDxIF+/lABcsXrNUUi
dOnpOfJJoK/VmUfjcQoczmPubICWoLzmZ6EtU/25CqhlER7gmerrM6+NpYPfSKuTrp7XRfLgdMCE
hr8vvnYWcaIwRF0Sbb+fkajnkBixtaCpT5pFB9ZiXe34f6/0RAMWqHnDNP3IkYVrGhrYy/T2vJ39
D7I6OnNorGyMpXIsAmu87SkmyQcnm3s0S0bkmxGUvH41UU8pBuWLS++idaiDRPXllg1+Phh2rbw9
XeI/Eafqj8rTmtIRDaPluNWRHOZriNt0hvj4777KJVmM8l6iUiVimXrErGdyJ0pnG2AQ/CH2gU5H
/ABw5RkcKtJrLvrBuoMQ91CepEEI1nUaebj4kLboxoQhWa6hRxUlMe4tFB0AbQQv+yYJ1/MD5+p0
jQAgAwDEUpHPYBYUhbn/eOpbHEHpfoMObUaS5FwV25+2bkKCZ5+ECy5i4mr7Otqcfwc9Ti2Q8GNt
QU63NtWDsw+Xv5xhyHLbTvxiQWe3Dn9uTDTnz4sqKnuQRoh+G9V/SU2k8hly/Sl3Z1vqeTmnfMLH
UtQPSCT23cKW4qVObB2H92IG25WzAtyjAgcLkyd8UPrmOYUGapSlvVhB5z7K3ADRN1fhdx9CkrrP
v+/9nVrLjUFJXcD3GXC4YoCNni03uGYUVGD+RbrX5zaDxrnoxLPMqPj+YlJ/Dz7WoEg2BWeWqXa5
Qky4YKIYSPGzFetCSAQsStTMFDcYo2DYRsOEdliZZFglYJkdAHi0JFY+s7hapCVzx2zVwxig2rX5
7ebHzNwOfyhEVcwWbV2IWERsg+flk/RhC2UOWHTMeqvDmLlJFCYzEEi6yPxxcYyZS8jykoR0sewm
+i/oxhFGQ6hOmexyC69zLNJAbDlKKuUg+L0wYdYSS4cvA3BPs1MMKVj++8w7qawZN43WzjdN0bgy
iTbTYaVq3vdZrYpjwkfL2ao7g8nLRBKm2V5sZVosLL2Nu4GRKtr4mqDf66Q50DC4+U0XKo96zPmw
KJfZZrsE/fwCBWbO18fe/0rTGprBcohoZe1YC9IO7qy/BFB50Itr/OVbtjmEOMkkswCA+EUkjQiT
qNMeDxmUxL/4s4vFVjluEvA+aHhFmdFg7Z3PEtMlXmLn2N5gCyogUpuBOkQOMXpIhSFLDpDIwbvi
5x7pa0HbuCh56dEn3jhnezOUL0VYWRyA3WKtfaslmQi3ACaMnlpPkjs1dAKeFntjN4TkIEUMb98v
odmGCrJMROOBtzP0PzwPHBqOCxwsafjdqzygW0lRV4Ku9NLgaipujRb6N4IzmWNsVXNyJQFJ46Ta
Z/n29/2SYHEN7qsYhjrMLxs1EtIRw42yCJ+mN8Z6UJUgqs1dnjSyyHiy21pLk8L3F/N9ValuPkbp
5BLMuoquyzNyreUuCluLyRMqIOIIwS/l7xetfSt7IrV9Ds9o935wXqQXha+6+sDhb5/9CSBRSCof
ql2MVUHcaQpyR0Ml3k/wNxjS09pFNGU3ke3+L1GnoX0TZuDliHwIzo8HLFcitzZk9iEhF69vjwQv
UeJnHVKG9uGJ6bzovCLJde0ziv/e5GM5Cq8dA3UwmgLSQOI+NqjWgtWfgXR4G3z6+dyrxSn5tHA9
u4XwAqMw75N8TlEDfb1nxR669oWI09zug+DBjdm5xuqJjuAWI6xAkfLhpWSEna0da//W0jGeA0v6
j4v84ZeqzyDMkYAOqGF0hSAwWkUSIUImkaLhGEl9Hf3DHG+Jh5rHFqyy3Grx3FN97mxZaVNXOuvB
PRkg5U/aXATKum4u5RQlDqCiKlnOzmHa9pbOS8P+2/T85l5Tp+PniDQB95K81qwwtHxmoqL3ZZIK
2d9uHdbxuyRb3CTQImWWY6uM891+KiI2jWaalMLax6mVAf9qgrSRp7+AqEQm1NI79N1jn0N3KXMB
7egaSPk6ggChfMXjzwEdWcYRAwPw0ffr+jLMWggdXv3joVidhaAXeJ+jQExsFs9CWaXrlI1yzsc+
lcebRyusodK9c6pw2o3QBd5ZTUcwFbcdeZlPwjjjPU5Wa3d2V/LMBIWVD3Cmd/xFiSN6vovXTQXN
AfNMod4Ip3nMLm5/FMUUH1fx7gArBlxkLE/hhZo+zmQMNm6aVmPAxRfNbkNV/Z5kNaBMB4DMlT4z
ICv2Wr4alqr7Hm8TuI2xwkqo1ExfqbEk6z//V9xQ+rXPcZCm0Tvn0TiuPFfuTrpRXrUOxZ79pht2
+c2HV8URoQK3o/oAnwNco0tFS7LpsI/29UrSEYHJO6i9XnHxaNY5T7iI41qU8lcn4XZpmwfzEtvW
3WzORzpNcXEaf+ICR+U0rnLVSUH+wkFdjiBQtDV7iGgKURKfoedti6zki+nQO7tdfo9zPYImVSg6
7NYdFu6pTcG8YnJJN5b4fXce9r5+LsdkwGrITPboGGvlhu8OTPcLM8VNlRR2rzmc+YT0g/gVbWUU
b5Dh+vhhbMXdW/EgcdkzRV4k6JZ7bGkY9oHcTla2WY0CdtDNa56RmY/SEkJyhH8xWWq8p2nu7O2A
AJdUGqqHzegH13ItzTmndl7C50zxuIfblwuVbzYmzM1nBFM17dDa91dauR8goCyIVrC1jJvWlPA1
ScMshPW4SfldBvEqcsBKFmuWfugQC25vnpjnxXqb2/+qd4zBvngYuXNoZs2KCdCyaHQYL2H+pwVa
c/uTyPrnkueo+uwpj2uB6hHiJOeSsPyCYxjsemSA1gcRN0m70JoLIzEz8b4hVuVTuGasnHLIyKWm
aeZIW6Ih/R19pMkaPijwVwIVMhdhykPOyjrDEWHyloPOJMY65X2FAammLGn218mccd1tiaWnldKA
X2yIoJJrNamjSz3MiqtEYp3foS9OwGCAVKDyywuJ1NlR/fiMNuUneG+0FWFIxtgEImEEpG9POLyB
noM/KO3DeP6WPmXYWf48LQkdi1Hpga0EaAc9UTuBJHc+1/LWWQYAEXOPoJPGVXh0iQILVLxuCmBT
+moALQ/uzd+ZHmvFR/qXt5QhDulLPDbWiCE/7IxiDbs+1TZyWxjshoyIWJQUroXfIT+EXT9E9tfr
kVZvXNmxRjVrts8qSIOCx4ImAVMJH/0qA6iBXpfuFg31W5qojLGVUx48G9hYwy0Mnha5sEPiL82W
dXv2roxKrXUsuncv4aR4W2F/HKISN/hEnrhwXWns/EszskKeU8LFKSzZJ3KHwZ2u1OX1lRRxhssZ
SxHFFGl7CBL/TdsPLFC1zXJHWwTmHLNO1sYQkzbU3YbxCeq66wyDenDKEGc0Dg4Fyoll5Bdli3Ff
6ExyeogMnqjkdZxvXCFNrsWrqa/FefRqIXQQrWIEIhFYPMbH/3FP5CAZ3asctWGQq3Q0OoVuVkPT
MtdFDTvu4BV1H6QZs3Y+V+yKJa6skXyp1Roz6njePC2khQt9SPnvYSYRnzWTz1n6l7PZZFbW/Asn
LFGpGHsFbEncR9+rXHi8vxpjM3okJpZZbhbC27BX9QnQBLzdl7jVBIpa1kQCkgTxQRWR6wd+zHuU
f5BnssI493R14DAQ07tbUDfNfH9uH6Um5W3mAHwNKMD0Ook4ePPiv2QQjSxmXHyYF+l7Udd1OCS3
tGPgK4ibCR522ZUuhRmMFUZIg2z+cL7Ruf68gPFTqJpiboU29MzL9kFK6ubOo12LPtpyF4mVL9wJ
8a/quIC92VCoX6gptSUiYYKygl1Zz81OVYvukTr79+7dyZHfVEprdvgPKkr/0hs9kfhMAHsm6KUN
H4WfLmQsgDb0LS0hFsnup2R96ZTDD8EW1zxBu+xw2mDrrStaPk4glK/PnR6AW8pUZ06aoX2KKViC
hlw7WWEkkb62na82c1ouQ9DVLhyZauMudNkEeDaymunhkDrzwDT703C1cU/HtY6dugd9hd726hUI
ludJpQuuugfxYJN3KcGLdjCFYovEH1awUbFbU1f7a9BSQ8bsvZSDjGDzenjmfp/HVl7zUmrbxQam
1oYoZDBllZenbg54CP/QEJHpEmJdPhbgVNTJcXc78+W0ro7IJYR6yqnQfMJBifLQ4G70mkoxCPpG
BHfw/XOtXt8N+0tu/Wk2o3VYmSJiLkJkz55LFpOlaQkw0JZ2PyouatSAV5sgBTK5zk01zVo+NCKQ
pgMHfhKpgjz7awRp7GJnSAERAKuGfbUgQ83qDRXWfCa7vXx3IjQQq2ZiVL2hqmMjkt4ACZwGORbs
HcsSwT/gKR+hIsy8yvOje9TlooS3e5L3zOmD41bHNRI6FYel81iKdBfPqmdk8gjWDmn70lJkXOBF
W1AFad4yp2ZiGlWtda0cyHqOhpVkFx54YObatvP4I53BWzZxD6OkPJneeaLml3NWm4ofQKOayNAd
7ex8fD2jr7vHNk+1hKeL9zjxKnR3PY7vznok8jdhdtjHZnr3W0Q/Hh6f7jkZebdkM+B4lJEDK4U4
xkPatFtmENTvui2iMC9ZEVBwscVYsm/wNOhmkEfqOnmw7McbTvFkGpdkNs2LfndwjmHqetkSRRv0
09n+uef1a7B/at8420PMp/ByVVPu+ILuU6AKzpBQvNOieDarLgmfN7x2g0tqqdhtSpdRDYSoZEH2
3NTuEhjxOiKG4zWfWIUkbWB2ugSqMdcb/3q1EPYRbOY1opXPM+cDBmiOBamBbGhxKcD5wnyTPEyv
fwIHNv4kGeKjbss9FYaUYuGqQrqbqKbgExb+BQ+x1JAAKmYIQa5sMJ0X3oyxwZJZP9HqSkytpegg
l8U7D3WcOUNyPcUn3U/qiBmpf9uuukdNr22tv/9PbSFsPGoafl4XGny+SIyx72NkKezmFcZa7x+i
PZdHYt2EkRNLd0j9BRTWfzirC0Vv9ecE71qHQZaY7QxtqIwkXmwfGomFNJT+HzMz98L0rYB8F6MG
WYNqfZeDF+lPUZ3NZPGnly0GlH7y05cybCc7UT/X6PeTNWd+QzeINE9fo2jc1uj5jXRul8yj8PL5
bEHs+spIisjEbXVRG6NsWysvv4RMf1vQakP+BxFrBjhH6p3hM6emjD744nPDe/AAgDlDpCWrvnlv
SrZxACk0G7o4XK+7FgFGNuAGYRG9xdZjia+10eX2AzCtBY54lhCFSVOXah2Zwbt7BPdHja+AqZVO
uiOnTYIjoMSlQIyr7OtVZwyJmE++bCo5Qvrj3Q4oz6RsGjnMs4gFJ/YM+X6L5PvQwwWEkama/2AH
y8wQ1u5BuQNeoU9XfSzC3GLvb9rM4KvbABNyCWPI/s/OFsJ1sJS7brcP2dNZsen7Yu/+svZz2pAW
mXEk2mudRWsrtyYkli0DiUfBQNHXN4diemVbg/POtZhUi2Mfrzby0J2CwwCaRnMjZzBNHil2alZE
MYcQOVtzh75QNrgYnGRjhszdXk58nhPpjd+txGc7YHfyN8sfP8Pr12z9dVOteFCXEQ2sEATy9Ao2
CMm5sTllIlL7EzlhP+NQj0XybgTLyaG0insi8c2JDcjD4ZSuvS+QY439f6r/r+WtEo/H7lvl7W9W
pG4sm7PdNxWOMep9NjK2hVhuHhIcCmCRfooufCGNEUkYUpF7UyNjAAgbnnQgUa4djX6Hxwjg0Pcr
rXsVuhPfjIUqTkwOBpFnQnocM8C5dUW+4oG+U+Sy6xgHc8eou+8IlCgW4SRcx4YuyLCYea2wTK6X
uKbP9hDPc8+hpODwMljGRA7WF55zKEtEZhCftGxb2CXN8/c5JGxRVEOncpqLdYeWXFL8/8sdIP4q
wIhPWDDlywMzuKMFQt6aEuFSfyOff3l85H3mS4Gp6LfBeHyh0rkRDuhNQKGVjCTQLUutKiS4ptBG
SMwqj8d1bdDpDl8URI67AQ8SkDBKrXoUqwHe+9vzpEZVTAycX1tl5xB0V0Wlf9rYbGCs/3qsZ4tu
xbh+E/ECmxlXzL5B1ilnv8nLny5V86LdgBc6Bza8ogVqvpcKcs6NGtYj8p7yZ7o2iK84EQbbeoJW
Dcmnhf0O5s3bB4V5m5owDK+Go7f0d+rGTjyz+wpAPxVJkU4ehVgjg7EN1aG8avMPcfptV++xh7DU
u70af0RKb1JtbvI29TGPfIfUUYcLk/7rQB3Dg6h15KE6S2K/sc/sla1Uk5TvE15b4h79YJu66LP1
80qqGQ8VRfXwA2fv0Cd8grXCtEox2cY1kQYWh/FDGleyltXemv4e0xedCGwZckV3Zn3KjL6EFvx1
H2M806lwfpSwmjYncVxlQAPL5jB6FwZJmNnGHAsBbS5gmAUD1LzVFUFYqmnLIJkabLjUja7xqB3T
7TRmPnLgpDEmDbeEIVt7J0EuggjJhrwOS4rbK7hPTDVFKmf3g9df6c2z2szitBBfBBmcsY8ccbDq
N02CDqfO3fL1vmCTYyOIiTUCgeLu2gjjlqQAzs7UN8o5zn/Kg7daUbtp2w/pMZ/6ybbcUqYw+0u6
ZC3TAiJd8Gw83GZhQzNnjE+OoashbR34zLXp1y13deZ4H1tzZAcFWIzIUQDbD+aLHeZ3q3Z2tG8z
RVhXtoIFDpjDTruW9Xc+owQD8U3HYy1mi/pQa462UkljEINRYaRFn/1+0U7UaqtzTA9rt6nSsCMx
HawjFFRbq/2SOUH3v10NjMKWw3egJJfuJ4BYa9c+wwGBjGU778AZVxXRt6fSxWNnJX8rfeNgchwZ
Z/v3y+3PrlB7pTO2tGe6+2LuAmtue5zMNKN/pIexkf7RdLl8cie+O1VlS7D6DU1MPNaFb2CRUm+/
AxFfAlbG7p146Sj3NBCuo6q1DwGeFLCREDHmvBCIxrzwGFQSOaFsC1VVV9t2Isz73FsPCJg8i+Z4
ZZLcjaVpCrJBKLtzHPIaxjpKllz063d6orLTvXSAT9llYrzHNfCOzO7cw5o2zqNYvgLgXTCtW0l/
BNCrWOgfGi0QwaPinCucCvGypjR0ru8P89mY2IMQdIx6TSRLLnrqze2Q4HLrY3r7l3S2coJuFbEw
9kIYLcPFxoHl1Hmop4GN/2eHpLz74LDpyqGi3R49zPzpcHUiCVuWQTkNEJ+9lU6fEVltPoynif+1
v74EFDgQ7wgSX4Rq3pu52rPTfd3VEueeuVdDT7ljQ2DN+eArhvpSyMUwzFjoBF2uEPQro9n9EJ8q
1usTmwaiy0eX/kahEEShIiv1Xne74oABvbN5LjLMYh4kkwBQgdTtJXoboIcAHDTR8mXLbkSH4cEX
/zZvY+vUzRpPYrsgfJWA9ckI/2ANpwyXzkzXE+d8qPRvGzqH7G1AM+oGvWFXHtRxMsaoqdlBXzQz
FfylCXHlm2VS+QbDnuRXXkqT0KTdLEGPglgZVnaw9eb6qGMS7+GU2WdYL7YUt5PRqq++nLWOhJ6P
FUOsWpAt8HDU9herIDWYzyVmjFoxY9FUXxk2DjDipXDQc7rUyWgSZtGfCxzIlbVxNt/Me32lgndo
NcuIwP2eNTfJBxFE9gExXRhkiXpBpDWbUv23X7wpdYtZ2+cJ1oEEqTYxaPtxCS6B4mwZxDlqba2Q
FjFsy3OhZaPZfUuVJ1YS9Ym4SN/CNNNZdchcGG4fKUQp/SSo+EeBfWwF4qxYKiKI8EYHGhRQv1au
+offnjQiHf2pORGzRL7cA2JD29sQur0+SvHVg+3vT6M3OoRmT/0ssfWewB+SiecoLgIk40bwJpbS
nJ+PYDDA9YblUmOUu9dWbOvlulyumJa9zEOA/+bEECAFu0SZyffNKSDbuxH6mBnqSDsI5CVYrySY
QamOIMZxuq91KdwppOipb07i59EBMzUzkYQE1dK1wvnZC3jN7vTncoKLzhEcO74vfdHc8bWVXOXt
CfjLiBn5DgILbBQIsy8IFnFzKfgimvaUHwEU5sSW8sllu4Xwbo9Xc/mcGTrc1nv7zlZB72STeuIp
YCpvPCBPz5REeeWXuCpbVmklvYMxpJuUOCDWSiyTwWsx6nFmlkrI+B7GinmDkiLzsEmVea8qaKUe
WP4GiqrxAwOBOWyIqOp/nXy4hGdHopX6FOxrx6encpMllDNUIs17zBFyCDx9WgwWE5DherIMCK7C
YawB0VSZnvyfzfj2xnW1mW6JJZecVg5zrE2kqqKjjWGE9h62UFVRjIgU5X4nwutyjY1Won6qXGbz
kWWmWW3Z4nFvvQbsTtXmSWuwHl6VaMl/tsghUQB/DIhV6Pcf+tHHj01SU/Hi+Z/9OfoU+YzUmm2P
X4cNXTlgHvM1k4VkLY9RgVDI/6twm8nZT6xmJWY1X7LIBzQtc+rtxQ0c4M7Kwpqw3Mdc+7GRoVOW
FNJZ45lI+40/Gw5u15iEMADgBwWdbMyvV8I0bNOs6m9D6+XMTfBhtQCPTt9fL8r0q4bbI3vabos6
/gmLoP4lMOkrKyXemT36APM3aQ2T6hLXv0b19akIyGJgduafgKJrklz6B93EcCOVdM+ZfMCk8AxN
sE2WdcibyLLQPYOdkWws3K35nSdALta0EH4BDu+3vUm1uOHXVzH9gk3UVb4Tbb7v8+9PFHz1nEFH
1sjrhAnWfuZNjdQI0TU0OUvLZ+khb7wMpFVS6iC1txF5P7FfIUSWKOwsqBFImLmbxB0c+JEfs7b/
eF0ReXFo9jwkqEeyIQrXh+0DZNKinQY/KG+AKPWuyny0DuVusuQuM8GC9ss0utGi4fv1QqKZEwmA
gPZ2VsfW7yAjmZxHvFy/z647dg5IaPb2o1tRlPEyVd8jAs7/JbYPuS9Mmzxv4KuAgtIDuK7VIhMY
SZzSJepPEdYwwUwnRr70zvolmn6zAU2HVLJFmhfb+Xx5cn2ClT0h9Io/sie6bg5zAwyR16cD1noE
h7E5NzA96XeERNP7IXOacPyTy8EMXNRxRIPC319qbrWFKP2byy2hFe4X37vupaU63TDcCP7RBef8
3Kv2DL8U7+rjLB2SY3kkJTfMNt8rbD+dcSJKaXMFyN+PoqaHa0sMVHw1Xc9/9nRsFAcZ1nM6Fax9
kopfcXeTVSWI7hYHhmicZyrXpFL7DACevegUeQKoeGrmPmIew/hvc8m7m8bJWLMaOYcoAGe4DrzD
Qx5hIjPm8Ln5wUpi87qUSfJgAQEFKducaU5GM5ctLcqbnikkZ1ln9Mvjv1O+NoBumOtQd8lswm58
q6J1f5EJlZ4BaC/Dffi+rqbRZNbdhI02Bs1/NX5PdyA7dlJOncxRKOl5pALVp/zeBEd8FazkOh5G
Uvx9H1PH+vpJLDUOtwu3TkT8ZxT12e3bHWiBC/COgi70EVj2MOWfA/0DT0UW2G5rVwaS9POXaikp
JMUDWJ2KZJAKsvBUV5nkA+h+x3eVXLyxWjLW1YFIhQx3tRSSsjP+aiIjNR00CKZZDEboi9PFhga4
mUXaizL7oCpoRnBgYdo4NoarYiDn6asKYFrZQd2VlKNCoe6+Dx6zCVB7DYaIrbW71WO57qc2tkhl
gVEjWnkQQYTLO3Gfi+ONYB4bwcEZnDM0NolYAVCZU3mBnn3SBCqBDFW6nzyWfbyjVzgYDKcUKEfD
I9iDPi3ko5g+JQjQpGKLD3HvSnmgIhdUHZvreXxE2ZMgUM/FFQHk+PFza4cRhAXutZ+sNkOyTHII
UnothlAnbaQ1Rfl47CkYjo3POFe6RMsZlB203Wzln+uc3qWDnpV8RGOI5oq+n7uU7a/Q+vYqAIuF
OArow7fxKb7Srd7JjRI7NyVwMD73TAaTbFdGauOHrwOQUr+bL93fwlf6orVHqc0BBUKxseI1XL5w
9OLwJq53AdQGWgJ0NcTGVfI5D8bHCrYAFyf1e2AMsKZsAF3dkVkFpGfNFsNROCR6Lf4lZs49DSp7
FAtTmMiIHiVgsHKiYg4l/P0w1Pxt9Ntrc1rttk226XisSeWUWEfZXKp2HqX1zKrTIYIo+XWs1RFn
SObNEX1a9p/ArmmGMS5CB0UR+OgOOCyq9paRA/B5pNIlrybtHgQERFdp+ilYfDt7uBe8CGGBRzJW
MZm3TPtD5TgsqPPnDxuBnsXmED2BrcQwyGBJZX2ho7r8yg2Js+FvodHfPIU7jCRLIZJyxlGa3MQK
6gp3P6vA8FCLYtHMmSjCR+8A35mk6yONE1M/GZM2td3t4JK9NDjdT2X920ZtWM3oChIj0D1eSwIN
e8B2wDZxPGjAm3SsNsSxALAMcDpFIus445yufqn76N/aQ/FxlXLILpRhm+h58gbGrXwVio8wRJj1
Fak3jNh0SlUiMuN++k0Gc6IAPclThciOMLpCctya633zaOdrt5XDyY8YYnRtNqzu6VQzMjn0hGUj
rfJaP0jbm2OLleTecpfX30GdshdF3xI8dy+YptGRFqdF1E743IV0aJaBY6WaarBh3NBIgVnYEc6s
K94O2CU8+p9l1CKYSso+E27Zo4rcuCzMDRy+Vca1cByPxn1MpE9qD88kpH4AclRthBQFtJACikmp
9Mgklhs8ifXkVaozvH6ctEpuz6tTlbBmpdcBBAt/k49kqyYNbGXb7Y7CnM3g7TFJk3WcZDH0CxbA
nBkQiD9wwKBq/DLJ44jMEvoR+0lBR/lePztkwyNGjQi3SgHygTYkOWIyOsHDL/MSics3V6dIKP2p
5m4S2XdKPOMaRShUpyiQaY9/2qpiewi/t9bEZooHrfw7J4B3BSdVd31z70s/mQQmjtoY/70jy8MQ
3+MbWPPFpNJPsC7y14KztkwIEY03uPnYLvpv331gqb5RrtBS4mFlVBH9CUS0AXBo8PF2NrKpAMvL
UuaBxQ1M+VglZx2E+1H3+3GFOK47USuicMIqpgYYAy5D1DmxJZZAqBlUXb7ojhUpSUU0Iu6NNI9f
E5KTzJWHWiDFl82JjIppBk0nV/Bnu+l/D91fB9xIiyrAz+BvO/dmBFv0Ae5uH8yY4apa1DvkDyoH
s5wygrToRinUNZ5jiZLHpR2OEcYLE6eNNJ1TgOKVPLSG/I/yA3ZZGigdvONd+AUbXjyYKadIPHI5
L1x349Ie1PEsZ+wvlio0ahD1i4+p+DnLz5Gdv22QYngFpMCq+ag93kODqsoPYqXfGFP5oZaUujCV
ZPQb8dvY6cqc4AjtbFnFpOsv0Ph8Xrg+K+S86h+m74RQQtP9nAd1OQ2zdqKMaZlHcBlvBRxFIpz5
thNZXMSZOea/Oek/SuDLAWtelVGR3+ddZZGI8FUQCJywnXrke/61tXbNOcdy7Eu68btsJUVzQ0Yp
cnU1iadC+MRDgRpHdV/zd/qDzoJYb6Ig+EbMKLibFHvc5tWwiwQ5JLDSVTOgnJzZzIPKzsC4YLAT
HMzFki5tSSeBJDqdKy2QVJkxjPE624QesgBwgUvu3y9D2a+kfvURKXKi3MtAEuYvr53ChWixzcQv
BR0z7ini4whMc3othfrt6tpGrDKCtUQQ0J05UcNylaQoL8Xp2peSRlbyXz83w1aDaK287RwWpPFx
C5W4FKbHBqLaFouzlpXqFLlOkscV12ln8nWLS4s8sJfab0ErO1lJ7okRq3BD6Sf09FlSudm2UuV2
/St7WG6bQG4SDKKCYunbdsuvko5aB++/tJK8m4jj5eM/1K3vXPC39Yxoz/ZtJ/DuF94z4bmroHdR
iGcYf9lK5TpCr5uZkkKXv0Pvncuyxg81ukUcUnDyw7fXAT3irdp9vKGnImri2kCpOEtzbr9I0yxQ
4pwepAzFIo5600V3G7EkBc4gsRzCxpqH4uBMyXRozAMurzQMBqal1oe2puwWblgz837m/iZXevva
e/vFT72cg1bczoB92f27dwijjHiv4E2DOY9osA6jkHjZUY52QJpEwfNRGCmt94WNXa4ElRYBZV0W
Rcj/pA7qYPeu2QWIPnf2bFOVPYb4EHI0gaISIELEHdUV2KcvCdPuwGTotCOt74jBu0AfxFcVBgHZ
IUAuyfcHg/W6MW0Lvqta9b3tW0lrPi6PfVMK7NB3LF+dFrNlf7dFakbDrxQCjMNAcaTKHxmN2i60
CT3Z1e8EEa4KJuV8cSUz/tnxcLOY0Iyl/hak7KxRYsrOc4vj9F+S0S6HoSac/cEXoNCDPhRSZdgs
IgEKwjDeSKOihI/88vbthEWe2mzQ7CnHFl6UGObUs7fgLoASc7lTCvhTogO7nV7fkUpuZ2IWvDVa
rffcmXGgV9GnjsOJanzNHyugipmxQ3cWZg+9VPiiQersANNEO6XgxwVkefOJ+9nIlnnup+DSVG78
yO9XsEEhiAqoQbhxFwUriZFhV4hKur65gOfa88fQ/asymaFOU5Qgy06aZruqZLfUYpyQ+t5KfIuD
d4gNFW/vKUMnlKYFjCwAAHqanvhpudx5jgwzCO6wHZugMcaVi9NEPewf7iLi2/qA8P2AIeEUFvL3
lOQ/qsnda3WLy2qEhB+enVvbtWqyuvcWPUWVKY1Wc7uJQ7T+v0JZHyOOF7OHcgL9VE6bTrsBIKJ7
4KPLIdiIj5EK7Hn5GwBfqqIKCZo1frm08vu5B2Se0MipV8S3TEnmUp07yD/paZRJdfeUa8ahfNk5
iNavFCjJENY1IKA/kt5czYNRg9Ywz5vltnCq6YF6bfW5ccjPQjllzpohRT+twul652LKbo66g8VA
0mv+M0yfs1Y481XqbqyvCWDOfK9/q3rz4TALSlmkev6wMIx9lbRFHYqf8yRyar1JMXZSsG68wQqj
UoMjQqOULnDrNRLft32mMFLSNKBf3P7xp11xKdC0xXdJP2xFOuSwLo0i04A68UAwXWm+u7GxypRN
90YQPP5HNu0h15vOgJA0Dka28RvEKDqMLjtRXg6Wo6QJFkVRvQ13JAUeFS0YhbOKowXNRlIY6Ca5
2Tt9g4672Jz98AjnIdJurAw1PWpnKPSnjPMQjmNtFLz0U8STnGw1q3SV4qR2wo/Ykl+RiBgwnmVs
2YR/PzDg+yQvunuES9509z9UsfY/3Vy0OImEiyBNJewe4xpta9OcW8uLkqo1T8kuXBJ7BpM6O1YA
ANDLBox2RLIVwl+8SPubTuNw2A6Q+9nSBt+tSqsnZeR4wokVI7mVKSs/0+fmkQYOjzv3dhC87Dzt
RhGTNIE0PCvFhP1luGvHqjTRXTR84AGsbS2fM0NtRCXl/TSiD75aHSdZeGF41uL3ninkuHDG6/gr
A//pvllWIx2Tjr/T1TzJaXr1FQjaTZ8gbCmvPspnKK9VFY65EJqTgXZ0vNVMfx2WkQ8ULhMMvjU0
m75eNFMRdSnWnPtujodyVtJzmEHkuZyC1e7HRtfK3+MU26q1COPFPljCzi6PZ7nWPPv3ArcM3IzB
8Q4aDTcc/yofOr3S659aWqLADCLHVbiu/PeZIfEVRAwe4Qsg73S218TDcL0a020IKN69SN0DsRW4
0SYdIdXBYy3kFSvlJz9Y+EVnG1ayIeQ+JJjQauK8f3814Sn9/AwfK5EgYg+KmZ+L93c5ATpaaXol
34E+u9z3pz3XeMhOAME2HO502aIzb9fzK7siqlotJPVX68bIsaNC2VHUCuOI09wniTVOjDVHzjR0
R9Jvj6ZcfpNnSgOUHR0HRXURnxQd/pGtRXwVxOa3OrRUR53SSGNhRvHGwPrceE4h+7v9Es5cYEl6
B0eMa4Z1MBhQA+TJWPMXROCUFHc4o24awWdEEFILC9tEgNBNqMDAEXadjG/rSKOo+pJ6Gogmstmt
arcwPfPUL0pOYQgTQynfuPpi7OaVM7U8SzPqs0hwZ4TpWLky+hsggp4H4QEegKzeVi8erjW6ySEB
oCn76Ve6jDheIrFVCuIa30gP0fk7dfuvF1GXXLEZSdPJDe5ONcPtaljR1V7TiXo+HNZW/LxBq83H
11a3TkXJ2/Nm8hzPJYjllFfXCGSTcn788Zop68gh9TPyE4Om7C4boNKkv/8yDIPhNfHllYpZftQU
6ef6dONSQ0xJxQzoN+pTv8yT6F0BPm+7PZ6MhY+pA7tiNXMwGNJ6UlpMXxytW+Ea0ipAQYNlJfdQ
UBx7sYTFI4hj+Q55lN2MBHBdkyIBL3odvTXm2/CtUV2tk8dvpnOillYpKfZ7hih/NvSIZcGI+Pqp
K3px6/An+o6Fw4Ge3VrWg6vGqSGelej1Jvo8zijPgtssLF22gj1loSWs+/G6Vk1XG1OUYYXvN532
sv6Yf+Ck+bEdFoU2htp5zrNo8b3yckFl1OkShTNKiE0D1Wcvv2ecmeuBPaTPl528idisdE+EpHbl
mw5KCo4JZzcqbwhwEaVSp0H5YslpzNBhkirqmWnTm15l4yGPHr7E/RFxKrT2EBOx7KJcN0pUg/no
rAyJe//RAx8R7lkMt+nuu7PX3/6l3lnxYeiXZwXoaqjIC1c2/G0nMALGRxfWmcOE2GZTKoXTkjED
Xs0GU1IWZYLRHr1UGg5I8R3lobRLPW5BMHhGhuEqOCPbss5nfcbZEtfzawBqvpodYAe/zXZ2/4bz
3ma6YXKGMb5VQOf4hW1BF35NkIyQW0vVaZQLPx3MmDrdr/+jQWJZ5ITmCuJ1+YciS4xYGyLGWhQh
zTnKyrAzS5LugX0iCKVrVGZfQzUSILX7lOSWX++7QaxrUQc/EpwfRrxhyKrXdWUOUczi+dyENr2Z
zvEbuszaxiE7o7g/l6okpuoBKegqY6QjZF0FaeDBx12pIea1lPfVQ0/nQOVDF3CVNmQvtiqfasxI
z6bIO0UjBqd4le4+PtCmlndRnIXxKlqP+dI2oIi+0mTkl4pFtWffnfW2/AqekvFLHwL2tuLrkC9u
k9TfxWDxqEa82kT5uklirAQ99mbWr0BPvkKMe6o2ag9i/wA47TEWiGZ588k6kWwUs1I/w1zW7EIV
XemI5hnBH4LMrrCUE2KJtEV98m7XHCspqK+Qfaq21dpAVV4b0SiZaxDgupWXd6sE/h5gAy74C9HQ
bRTTjqlcZqb80GSEOzsgUg8O+8OSqbW4Yai7S9HcNSgmvc42oSuiEc26CAa6ei6N/6efCz/aLWub
auELJP7r16NU2dHCB5L5+5fNe0Yk6pYbwKsSzBTEmNhUboOLyXC57cbJgRo92KKVSjZOfJ8SGStG
qd3/veDK6h/pYBhQDGUdmIWxZnvvIH0EjL2TRDvlLoN6yqVRfZp4js6RbUlM1OpdEnpnQoDZ/Dua
ZVsR0+SD1FYB0xBX4j9B/1VyPU0E9qEq35mIBJN2geMDgv3bv1owiHVS8d4OwbNUSwOx9GUvhZXt
QPu8mnWFzsoPNR4PANxUKrbaIDX3rp5/CmvNRAcNdEa9PrCQkMHhYSVg4Lw7wwTGEat/tNn2LL/I
kzFhcukRXyIdM83LCgvxRd7JJWfABkXKF+Rzd4B41KmX8xx0WQbZM/7eC86EUtZQqgRI/aEYJXQM
vK1vjISJ12BfmKPF+Lnf2IiIKaYNqW+otVduPhzjPMXmU49Xabm5wl1hwamLAaS+x5R7yA3++7x8
MFijxyDasFSb7h/zdlWugyJ2Rc/izQV59Y1ibFBz/5CjfqOc43AvuKpyJl33tmiexiZyVqbC6+uY
n8NgEU3B6XA74sDXKEnvWne+7qOs0Lh7cWaXGOHM1O/eMF6mqBVIohnUPEGlHMGhwJr3d9XIpE7r
OEaynJ3E9fLhJgNan+msRt8uKgScFGDA9gvKFspB8SLzOs1IKFM8DMbyqri/YII1P7TazdZOGuiV
ec+jAA3UQLyU6eKOIFpAu0FJNpGw+wrAKKm1VwFZbAS4ac3aghUc2fqIq5ZwsHauH/YlU1vlDqDo
m3+fvmhnB7nmgSgKO6TJTulzcNPmEtaELFxABMq+68ryQpqi/xroLT0Qld9WDl1RJtmR9FcjJO46
hw514Lq335hMkNWCpHZhzUnxeYq+69acyzPaAvNYX89MUqRyCpanre8QAwyV8qIaJuaE1v7nHMsU
DQubdjVwbEDlyZV4mg44yZPLTkf2kRKjtFgBrn10Mmte/gFQ4Z6UWJDyXU7E7eR5FV2vOQkWvSGx
hyfgglYCnRfXl59Brez/Krb+dFuocyXmXHWI/FhpaIlEhI64KklVhkAU0kibhKwBsjlSwFM9jt0y
AWqdcC2KVM1R9n53wVIuqiLn+AZ9f7IZtEJDjG4tTzf9NlBKtagR9d49lJaztjWdw1vyw20g6bUn
X7wzDP7FQj+5IuoNyJmHLlDI0cXSp1/VLH41DWj3MoDtVcoJWlujRQR550FJbI5VpQnZGlSjnvp4
RVV0RNYtBOSycmKQoVPNI7yrlkdoDMdiI1w8qbjhXxikMugFJ0BAlcTrd0mnfkj69BUPCylOFTtK
9MCiHJ8e8Kj5cpPqgqHXiL64JPZ/pdVk1W63e0yFF9ALD0ra5RqITvUnAVCGpmGvEkrmIcwf74J1
SJraNxPHPtxZI8SCkPhVnpQPQxvUj3QYKpRYT6l6lqPzgovQrdG10qJCLFFejFKpbEtHujdtE/l1
qP92Mfi0AFxZKZ2JMZ5HWnkF4xyOXgRCweEra9kR9/KX70WRorZ2qjPlFFRc/NtgaxV5Bfjb1IBd
Zx6WiEQGnHCeK8zdaMvZ6bKdQbuK0WntaYvzrKWNvQgwA+KwRR3Yk5h4iAN1j0IxPcBIPFawjCK+
UBQuzXzPVUJQyUK3Ak31Q9HP0Z3CTZvphrFjqd7s6oufUTH6ruMNpOpM83s8/SdttWyArb46jWNq
NTfts1sjudmHFLOzUTyZGP24tiq6RgKZXNkDuUMBULrG4cfAglLsglEqeFpGLnU6QHLIO8kGf++i
wVR73yvpRq+3f+3RDPhZ2c/biKzBMxgq2Rh9/ozF3583fSY+EgQeEuQ++OeJB0juMjOTLwvkWW0v
DVu9hQOE/qN3DY8o75TFedUpc70rlkBe7L3zJmxxrUcoqIAjVOsvSnJJprjhHiR6JGL3h479Bdsq
Gc4S5RDQURP9dbNZTBFdqAN2zMzwlGj27L6tFKZbwuNpZB4n3dHfPcOOWw0ZH2l2HQQ8XpuFCk/C
WW4xXDNTNVdeqCpCS3vdhyOcPuiBDYPFHOyxLiAfcHgabT4GPYdNaCxL5mERWebfnE4477kjjmf6
Evc3eND2xeHSRslhSf+kafcHH/YXd9X5ZzzSMIx8q/DIeSj0Bu1/82rpIjf+0BcYFRdiepYkf3U7
mY2VzJto9DaewyPB8QrewLuZZXrd694qwm/vSVKR9CjaqXrouZZhGC+JyekHk2GXjYAJyayOVKX4
jHe1Yi2l3GrVf8JUygXeRsObzcjDC0leXdKaLVd7zszIPHPRNsDW65Jl0LacC4SkrACq3CXX1tl3
JthWAdzUNfH++vI82anoeHTkfeD60bUktmP6mqWcqpAASdusosxdvs6UD4Ra8ItTXK3D3CSH8rlB
CH74qfOrOuYOsSrWQ7jSl/3zXyJzXph+x3DHlWXMAbTj6AItfQSBE7ep1dqDyPFg4XaUA8t3ZsGH
NzYgCVOcx6/d7VFoxunszZqJ6CwtdwJrwPz4ZH1bXO5g+gDXikna37rVWqQQCTv+5wpHe1Ldkycj
7JWRra3QLS93VHNatw/dT7l1VDamOZv/74T/xlaHoSEeY7NYkOj6QTKqbHS4kihxakpmrEqwu1n+
MRWUNfucb9OUAJox+9Rd1qqhZb9nyOl1XqCxbvzNTYyufJiaUwBPFsFhS6eQTgs72RMEUVtXgxuS
P5BNvikHs/nsTvcS5usTieNGcX5735E5p/irH/neN+1yFwFsMDi6wEmC1atOgkUl9o04h28y+5LK
32wTYyKclRaa/a7xJQxsXEgZUStxWNIp0rZCLrdh0jGewLsa3+qJT5oZsaWKNkFwWkTzoqTAbD7+
BhG9CvayvZLOaGao7ZA6Gveh+7w61A4o1ZzJGP5HX/vVA00Jg5YmjagbSbhvjbLCvi67mVsdtXFy
Nj43/hRVlWbccSRpjb/J5zGvvzvS6nkxbPQ5BYLlxa14CEqVtQPgiT2JZ35mddX4Eq5T3QLR6K4e
my1RlySCgxrz7iq0ImPiLJwCP/2+UgeOhOH61JxwQfzpjhxvtM4XyJGsuqB+MMwfa0rFRSANN9zt
zAwgttcbFnSj8A+ue7eHrMxahIUwt9BHeyUb821M5El1n95r7Hh2Izj4ZNd74783i3wVJ6CHQGZv
oh4An0v6Wyl90293CskcpzRY/Ekp2Zoy6VwbnL+GUP5m28ALw0tiuQ+qagTUBFJj4TYlQ7z0/y5K
h1UUzVdw3VGouEehpIijvX8cjua+vPOFVJV5aHW5qTH+EdbmUM66/4XN+y4v/y3unyXnEL5adLTN
O7DVpT0YfZL3aqTM0lqWvs5z4QMF0oBvisT3/XU7X/WTOC8QFzY7i8sIsIwcYG+AKB3HiyadlaxE
JN7F04gF6oWnL2EYJt5mOV1yVhBuS8/TO0fCKDBud+CMJVLEocuMBW9pLX91OvAhh4uoVhI5E82d
iZLoX2MmFeXtGQqkAtrA2mC4hJvBbgPtHo3UOhdAfoXG8Va0rBKjqhS8its3Ic3eXT13yGBgfG6r
Wz6kHLsR6lTJkWCeThSm0nnGAQMu2bYqb0SV1svnZCdeYodT0nkkhNMPk74JmghzpPioBB9/H6vP
/+REOZtppYnl43yugoFON2AFseINkWCGoaef02KMMBqTW8i6+i5kxY+sR3Ldit6fjv97x06n6bO9
a06kX4ftNZ1t+MixcrGNN4LK0z//L9Es5kRDU6IKYYAPLkpQrXqTJYW05O/NJ7lSg8DOGHyDF59+
olrpqM492rH6CMqSXZOynhecDY3hbn6pTIJYXPIv/QGZXc9yk9/papWMsc6TMuCgBwWqPiAY/vvD
n/Vdo1rtc85SOmeVuUMZUvm3KiG7804fBIFcgPEtQntpbZCF0hqbwfKE14qeEe+gpXAsWEd9e4rw
ugZWUH0nMLRLecGxgwiCbnynrLeszNt16cRGzK2Al4SL6nds7GZ9Fg0MADMZZ0IhTEI/XKi7WWg8
26MKCLsiZlsQw2Kr2tA1YmbFpDskKzY9rik5+boallOt40Dv9bWDFqNAy8KVyXsSSbB4H63PlNeV
YJa4RyVUjh4GgAAqPzMRXn50dIpNmQfNOH4OUBtlyi0xjTdyf2Zo3Ew8a7580IUVM/FKUB88uxtf
gQTFuKtq+9Q+D0PnDhN2Ag1tM95QtkvZGLysCDGl8oNNcWkB4IvaSMoj8RjwpL6rfkN+EGkjO6sm
EossidQ0irnBC/Wv7XGKovfeQxxfaVAEitrU0ANZXZc3ueDs3aPSOCTGJMEsG7sP3IdJxRV+/n1w
b3+vCGABBp8A2HrxO/wsfthw9v+au3QPju7yw4A6vDh9uH+vlN7HRnkuemGmqgKHcKISm57uVd/L
OP14PpyncVatJ84UxH/u6cvZS/AX5HLXox3uNuiBJk0cQBMheXGIcp7Veto72YygOiTXW4/32kCY
/xBWVWusLGB+MkMb6/Z1RfLwaUrTRIyz4w8yHZvD6Qdi3amjwMzIPwzCfs1j3sucGkq6qzkauMJv
7v1JuEPJXEFfUxv37YbSUVWjVCtg//+k4PFxJBRULpAeOW0Xeo3v3pdeO+SbERLLMNutip911W4e
IrwYi9DkrtEVgsIcrpLQKdFRtxc9Nij/FDgro6DySTDlxNdFrxKwUwUfL0vyaUbJTllc+EKJM2cU
0jN2+kzeCBqXqjZCDmu+OlwspCxMyzMmC4pr4QXUhroCjkz3WnNLwKtB/YWeLfAAFf/3YTee/upB
rehSCUFoU9xhP/HqldE0NGjEa6xNnD/4kFc7tIIseyfHESO787EZTYLVedIJ8gZ2Dwm5CY2l8Xig
cf5pcJYbjwooXHS9dL7U0OKdik/KvaOg8d9zSpAT6Zsc67kyrBDT3Bip8fgGV03at7ALQTRcqwUt
kwWzkXVDpvWmCqkTt0p351NIh6KywUNJJiPaJiLmAVgX9N8c8TFIV/kGoGsGhz9nm/Xt2oBQIEDJ
ll9JPLcnU1h9/PJLwre3AZJIpHfY8OK1F2OxjUIofc3dBgYwYP8o2Kzs9G3+XnAjm8sJvyukmg+Y
w+5H6+KhtQLCk3y1fNCwVECpvSJptkW8BxMs5qKJ60tSOgTbKvJcd9dCf7zmlrs1bYxy/5Fmc/D+
yAB+x5248gJ1Gq6LACOl1fFij9SfcHJ+uBjtVAmStskiweU/b+/D/xq9Wa3RQHCQppVLHeIy9Z07
/EJ/NARaainJt1pDYXgCnJT9qRTdcN8/3DprMkYCz4SLbjgksmZIJQpWiMZzOel+egIX9KBusEnJ
U1W1y5+oIynnAYvv7G/rZKoTEc2kMXKUWT3fW2BoT8D3FC/O+e98QscqWE7uUs/7v6yJeWofmggc
GLuBjMFq5PJVRiSo5qoJeL8gSbOJGu7w7W1y8mKeISEtKwqslAkvzH2cxh5BiUVsk4tQZpcT7S/z
ZieMC3nFfG7P2PECYHzdaONun6n2ez+kaoYNrNeCBSjxHj30SDPDZPU3Yt0SNEON2NyO7LkiV3+T
LT58XCvzMzNJLY03pUY0EdfuaMcI33g1vtRsP2fGvhoPwqVMJiIy5DQQx4cIJupyoxxQcZx6UygZ
EupCdoyoL2Za9uNSUqpoH/E29KhX9FnEly2y9gV0bkEQRbzjGR6Q4hFJtLwaoedw2iWcmEuAcMMN
Ii7fJRxfVp+JbjghQxVeFSIsQYsIhXr3XovMbojghEWlRuppqehhBR17uA++1kCoKgbfPsaA314L
JwUrrfmwVuAaPfqYvx7nj9KzrfePRvcAZJZPebh8UOFxxepPR8ZjsWn9dk+SJP0asJUqJzCRUI88
+oOpfhisjQzZeeMjpUT4r1Ww5F3S8TUhIwLCEqPGhaFZQ+ZWEP3TBP8NR3EABeLafnUdnyfZQoYa
ByIOcr1Enmyoy7gaf7xBdbRKcm6QAsxu5aePI0Jl165bWN6Pc+rBq/ksbhePlrFSA0ItERXeGJkU
fqYrMLeTHiYs9bE7OMbqmkyyrPMd1G9mZwDwtnBr5fti/VX7E9gjM6fvP6wqeO+fk+GoZcpKpBeu
YqF8NEJUw1vnWdUUoVpsABPFFB0/kJflmlpeHDbnbJU6V8mi+zabFt6b1OtkgQfKZx9tTSE1rVo+
cjYP/uRhf8N1OwB8vKoRPgp3iJp8txf4TUq5MPIkxbPUNjejlsIP5EK6AR6Ktr0ZUdTwmdOKLnOL
z8SxzYuoMOq7OYYJ1MT+pQFL8qaLmEV1sv2CI45cYRhEkmzsD8dyyMwMG0YaxcY/uq6L6tw7pOHC
3ssNz2+FBu1v7MRDqkPMlYaTzq2JOZ4p5p6n6dlsmmmiUTpepEZaEBY/59/MGIA8kpNhfKgKzZ6E
omqOxX3/GMK6qWERRBR+4l1frWPnpwhaiNOIM1MCw4UQpllYaevm53qo2QgRTTqM6ieihHJ+n6qw
nu4B8/g5PnKR+tbq4DuUIqCCt4OhZmH0lbHo2SRQO7ANQVwapdOqDWN/B/2fTadwoZWZGj/m0Jzp
FlQL99auwIt1ETrm4Br1Od5tqEcOAyQ0o7CH9+TJakeuZUfXOc/apGmseFDEEVcxPqoCOJP/eLxS
z5L4eQ4Eelq/rwuVbUE1DbM9wo2dKHilFmnEEwA2Jf/w7irlmVC2edXCFiEeNZCMeh3lq81maYc8
QrWs2bA/gSDh0t6XggZYVbHwSd/eUyvSvmIo7Kj1M9EN3Wv+sGom/Up/EzQzznVlSP1Wbwfwemp5
EjvlJEPY+VAuaS1kwvOrh5tBhEWztLslAfxZybTIQMYzAgb2wVbBrvHi9/awICeZW4eO1a71INg7
DcLHPZ/jpX2tMA/9fxJ9V6f4v8B9Cr4fa0PbnVA/7JZAuRE/vqN/Ws029TdLqF5YruOxadxOPQqW
jp3nT+8pUuGhLsRpLmb9u2KbK3KsZB9yql4VXdNMhE+mmy9wZgzlWOURtzZm1HqHKTJIy3QI9Wxy
sNGrVeoKI5Xs5Blr0yN+UfD0okqj98YMK0QjvSnAOjaP7LqyvORcWszC5qDGOkjMGP4SBYizrkUD
9k/+Y2vI/QPCB5zKc1J2xSQH3nxUaMq/dbTqcFAhRGsNtjU7ymZ4Xe9N6CY0QdBwzDlCh/ZNN8XI
kKBLGAQFVZZZ+N/zWDU9kwS9EKd23k6AAnpO3tk2p4eGLeVC5NMtzRt8Kg9M4KQr4pPAcY1ubdFF
0ucTTevo/D5SiGBpvWCFNqjvvLFo6gAgvWKB6/UQO5D0PrQ7DZshZPjf1tcXt2dSOX6+V+3Vnhfp
CS6Y0q67tKXi+RNyEoZYWa2nI87yhAKM+pFTLQ/gA6v7sxrRCYxI1CkReRH/yR+D3RLn4bprUDS3
EnPsM3CTPg3ovMePbsIzvAWc80fXBJgRlMrs0+cOTaiyDEphDesYt5rRwjrgdVDxmYpzbRhZBclt
T/YrJtD8q86RDIy6w2t4JaRjIRXFJ3J5G039adgFvaXL6up1eAtMBESowCA9AX4cFFGswvgzK3op
/XJIS2vrpo2+O3+ooHectt5PFNQmV1dHMxr4RFeOXsSW8VcghL6VlW4rEX5Dpb3m+OUhFCLtmha4
gn8kWHseauhqJoy2Zefi/n1F5Vgb0qHA14jzpt/ALOkvwE8DiITB++qrEtcVQSwqetIUUlZTTLqN
DURmZx3nDlFWmTi78xPGtszXCw7mzKIoTUJSSsdSbSopOlShmDzmmLYVv32WHmzaNc4e7W/5tuFt
KptKYoiR95akZMxq41q2/hKINrx+/Xjq6Pf7b1+/ncwTK2iGd+hi8d/0Ghsjjfi752tqG59JtSQy
bCjo4wiuJ3MKSuGhQj7jZv21Bm65Qzklk9aQu3PhjeNlprKYD3Zu3wkLe30/7yPlORO49N8ojs5N
DrDvb8Rs/bvbeZwwCQtUwWsvYO3NM4lOBZfJ75Vomwk1LJ2PivvvQGBZtPSq7/UqnXDfak3uQIQ8
UGrBvMvIqsr8/RPTZVJ6wHGEgu6eVcijL6iXAdV1TirNSA1d15KD/f1TBRGAik7hnnKyziIsJtCX
phdTvaAEdqZLDSYUGXabX5KRZ4uwiTUxniqHeVC9t2mkGiFbgPwimrbo+gd2i9wp8tCw81ap+m/d
vT24XjdarJWIeBvxLge66drmAE/amha26d42NgilhnCeg4Jwo3xM69M3UJOv+OZvCVgCftebmCmk
2a/add7IfXja1sowwQ2I8P8eb65Xfc0usPkgyYy2ogPwO00A+1WKFXfA9r7KVxn5Dh4x+WBY/e1N
QfAV7D6/Xp+k0fF40T521P8/Ae2L+Xqu76lOBAouSsuhplmHBtXsx8bGXzbQ3q2Vr307t+Y0jzPL
WVrz+4fDz/1fgvhdveYKOcpXpyFvG9r4eENfn6AR65T7rzTNHq4UWvOXAy5Cv9OQvzO12NB7+Rcl
0v6e7AbakArZsshG2mLyiLTjm3dVqzi+277uhneLN2zqT+tg2Fahe6lN9CY6e9xZYZ4fdFb79B+G
+oJpEkKkni95HITP3BjY+IkQRJAuYFP2CXxMtpo4pLB0JbxT80TyqDSIhmPlQCnOmlPBC5X6NT/f
pv/6+mr4sABu5Xm5RUBtXX1lN6zDKL2wTnDZWBPh5+E3YxPU411YpPLr+OOZWGoIJdQ7tHXblkFF
TH2rW4Y280kZWstg3QGSGgX/v0wkSuWN4Q4TMgCilW3xOtRZ0fuOBOrhgPnVPQyCAZz/zyGHQKk7
ZoWD5RUzp06Kyvh2Wvezep99no547B4pTJBKeFM16yAeesOIqzUOL/DrmAN8agOmZoX7h6qdycwF
qL1pZeK6lJpzzytiu8P9qYuoDB8ERh7+uNHjW2Yyg/0CXEcYZ7VgT0WEW23qvqpqDlV1UeMRYpbx
PKmIA83VsIQvUWzBhnTLySzv9Hz4ncdFh+dX39mtSY0xZZaWZtK4R7Y+2Dne4jqPKp07w/kO1jnK
mI7rSMN+7OeGHBNqPJNa9pYy/GeuFxtMd+aWTfIZU23I1HfTsn0UECBv/Z5NnbD6FK4MBEprwoNe
UP3w9lbTtiiaFLmLUGp6ThqadLGIyNLmP5wFWdLfo3dGsc0DRY3D/QdxCyXZJldR8vKH3kCjPZdT
RJhjBhJyhW9iVvep1nJ9rR/+MXLUGrq2o8zUbdlBcULATcIyPw7yzxVr8rJe4urTGX8zn+uGHulL
RdsdV8iCwUwcAohW1/oxjolqiE3Y9zOD22cV7YyySo8T3kSP7w2wsyjENMMumKxkJKrlWyw/JaYH
zo778rWCMkxnw4YS7CjVAzafk0Y98g/EWXe6knk6IFO3b12sLkOJqPmmFSYnFfUq1tPtoJWT0uVq
z0njgmlu+S7VtEe6jueqfh1Z99OJih0hRvAkX0SJHCSrog8vT35AICjbcmJ1IlQlIZL1Zi2neWZR
ae7nVdEsrGFV49x/VFH1mRaOTJpB5Rldpl8J5wUPSHx5Dy2CCFHwbva7vyhtEAru282HTK0GM67Z
VJx4Egkacaau6Zj38sZiNc0Cb5RbVaqmQFsLrkUfzTIJSIunqmMVUDVrdNqqoaXD6j3yqQRRtyAl
3PJD1S7z+jb3k7ZQUpmXYvSMxOtztEmCcfy4cAUSSmI6N5Fv/MRUIqLcznbS7CBSRj6Z/czZoTpA
QywoUW4PkzYfjOs4xomYj4o56gc5OuxYtQntcc+PF7juPf2K5NrYXX6RiCb24wb4txQ5k40K/M5g
pwYWtAur4Hf8emGspR+gTK5mCYnRqjJ2FjGy0Uq7hkcRVqb7e48cvJRcM49nDFcGeJx2/8vtpu8g
o9OXmeJ8DZ3ePRJIhJh6TJZ/6Ke5qgPZXoGoQ0oQmjF16tmJzr44K/F+AldmOJJAXtTJ3bVEE14F
QMtzAEa4PI7Og7htASOGFADnT3u9zQzZrcasPLvltY7F8FYFsGxTCOTghAQ/TV2wEO9y/UuFQodT
0KcBNIj12RqksdIxXacwVAdpyA1O9MahZVPXg/kqM65oHah2pl9C5Kkx8rhyqrgKerkurDO6Gsr1
yfiq5sKWYx9PPUy+SmSfY8Z89t0PC6Kb4qM5lm8YoIDZKP+Io+3DGaWlBT6RhvE4000wJTVXZvF8
2fLAEFGQ8o+O8rcsQy+XMZSJD+T8GR4K6m7mKBARTxi0msKayjP2umPMrvt9EyG8SlsayaxzjVXf
f3erkHQIjl+TK0Geu3vxRXBMkhgvStjqRfFKUf2mJ2En2f8PyPccu+wfCYT9kT4TlY9i9kB8Mjw8
Grfem9lQdxCin3nmJ1QPHmr/jjtcKtu6lb/aB/F5Kwb4q78MTHBTnRlZ+vpPZCGY3KvpySXXVPKf
BCV8/WByfcEIIhS+B24uv2WugL761TWUjGgZYEZT5uK8sfD86DmAflMq1eikoQKwW3VDKQkyiNJv
fLZXcsHoFYFTy6vzAyutPdkmRZIwxjwdIU3XOS4+ELR3CVEho3pIUA+DS6+tSBFjV/xhWU04zw43
vou1AbHNCFfY+WsElQeeXGYOUnkaD78OveTmRoWRfo9xBxvoK+oqJ8takAyWPP5T8E3G+thVpGqo
ABvXMuecyjvpWxPu6NOL6ZvKaLKdQWk2LnxFbFVnlS2v19DErzStEDwRgsFcgVG7EKrH3oNpxlaP
MkzONfQBiEalJnsF7dRRTldV1pg4SFDi0GAQHMQEYzTZINlpfSAs489pf/mM4HF5yelDCStsm3cc
M57MgZMNTl4SLb0pCYmRXswpcEjosJquBg4vD6nsyxfloUw4toMLxtQesyEkj389sNXST0gh9TyL
Mk4naJ4PRxcYa/+HDb6bY9EGkCCdpOtpbKRqUhJMNpc/PJi7A3M3OuPqL+tip3bY/26tlCP4St6P
EDDDCxjZI/QmaP664rpHvmjhzYvTw/2yhNjKJLakN43hitOHDmTAqRom+4mQU54HT5sHAY+dAdIn
do3KYmw1/v++lsu7FRTJJIdxd8VsLOJYqN+OoABKoaun0nd8v3PyHlhb1IB3N8E6QmjZYvsqJKjn
XOrcaiX/OROMpdnZHdETtdl9cc0wh38sjKXMKCpjMdKPIR1p3AuwZv59geieET7XOTfLacCCR3hz
7o/OFzLsZRTybjc+yL6Q/1w+XY7lR20sTxj5F+hC3uwWLc+Aq1grUYKQhStn9UQD8oEfETy/uc89
dgKpdi1NqsMfODjH/spe3k7oxwIgCepUZdg+I+Z1OzIbElCTLuPAyw0lAlAf89PHDuA/Huo2UHiW
8O3KRes1Qv+tCS7Hm6usA9Grgop/Usra1vq4cphxWjY8ycXos40F2ABG08Np5sg7NweIZPMIrRgN
KUCqOWGKHmDqzmIzDT6I/PPLulIsZHgtQ9Fvh2Bwm2k1twVvmYdGIKPwuBFgKBjPmQYwlb2/OlC2
tuA/8wtbZ8FaWTBoNYTK+Hgk3+GWj76jpRM7MSX1kDeHDZz9fg9+Nmhfe3dD7JLdAzqs/hqu5EEh
TIhDCfBH3rOBEFlEetWtuwxLWR3eBj6virS5Q5MhQ404nN/heSpAch8BFsUmCqZTafosRC4PZucC
dq1hCgGZzaX60jwR4P4e2okSWqp946PecC5OL83ZKBsBW9VJJRw/Yb0ozBtriyJIlO5inBBQMyjT
iZaP0+Vil7sDZOpQ9hD0zithuBSd1PL4SFPCVJbfMYSqrBfydrSJdSde2bn0iNNv1FRljJikfKNL
GK4wAGsINgDV2dLJ543hd/ninIu3mIGCENvlh5dC9rxZj1TPPx1yCqYv7+zbPqtXYtWo2DX2BRWR
6OvIIEhQR8xsCnIy9nzDXFi3lVDo8r4otT1pXPOcYaaqZNO/mf2aBldKLL4Hfn24IhxnMkKOobwM
opbAaPrtU8+2h0MdpChOZgQqbHhWm6pmp0oVS7ALTivOTGwceo0bKASuheSG8NI0zqdjRSz4B/zr
qk69SzMhriZncvvCWxgmNxOo9T2Tr0Pbu9jC8tQtd8pGUHuxnEp9j+Wdx1M8UWFzt8jN3YtmOlFm
xWkK+PTfQ0h4ZH4eMQUzbxnaCne3ns1qb51NGPuWNKQMMIP6R3qHRib0/3ee0gAiQQbhf1kIE3+i
YNkkBJflzS0LPhzsUWSZkfSqDd1xVgGwNO/j+fH3DYldymaHpAdZmfubjswrUn+lZQEd+JXFxwIX
bLxLrDISiV5LYxkszzTTgwAdCBJmq1clT5S7dUvxb2IRW9HFppYfzVrT7vxns4yvN8SGpovBz923
nK/wwptql5qLRpJIh0cyhXyghDNmWchSHZO+h60HwAYqS9YH8PgPDc6+sAAE9RLQaXwosyNEHFLy
ND7+rX16O5n5X6zt6gxyyFwdRXjW/AEWy2Zi7OMkFmWiS6KmTt9G8I5mZ5YU4CakvUZa3l6s5p4v
CvC+rXr5m7hvbsKOo6ljIgzUZp8nxM+2RVrluuHAMI7vxXkAcLxV5pbb8ItS8FTrAS85lEDGbflp
sn1w13U+Yi/0RSBaEXX8r3kw5qMVsRvq6rN7y9IfkXNXZdZPkSJ3PG4rSomhDx2Ff4ZRVZe8v8rD
HiipDeAxqIGPEEcLWZabjFxPKLXuOrDH6qCtAtRzyyKDxDrxONqSxXbfS3C8JaKG1YOkQpT/kCCb
KFSPeqao+WU38l0cSJ09gTXwXRv5N/Ed8tA6O+PbBDbX6D9r2vBtctV6IddK/PWVKyHODiyxw8Wm
tStkocd6sczlpJa/vQ+USwqweUR5KuCSiVQ1vMkPgVgbyz+uYliQl6QeUAN49rE0MNTcK82fGLz7
HKad1MeOKHFXzh3ghnKJo7A85QXVr90YcYxceFgtZgNZg53gbbO7MHJIlHx9r3FByUs/I/jYzQvr
Xd7j0dNiw++Kjv7BH9H2vSff90uhG4q2UQEc0sjGcHUSM6gA5MUrZNNAGqsdp6gogCG1kFZ6L6C8
RVj2ah5dPt2HAC1m7V/0WJkDKGyQhS3fhLpXs6MQAKC5T+0rxRsyLyj5u9vwvujK3Ht+TlvuSwSG
uEzosdm5CvDsnswCUJYon20FEEZ/zapKSIhnSdQGR+XD1t8Fp6n/UDyPfMUCHmAv61e8e3USrYqE
OXnQTrZtyNcwIGgRPlPSQ93QncvfEZOIVPV/INeoFHnJwWGnoYCUdLW2+MzBKpvO2yS87uUDXZFg
yaojP3ez+0COywF2Tfq+V9yhglf5yK9ygQ4wS8LB1ssACYsdU3RCw3wc3/5iHrb17R1eccqRQ2iX
j7DGdODZwoyOFbC54/zAbjzN7Ctw2QLK2TezOtOUVJwFjqyFtu8NOXFhdYQM0J84v8DeLgl0qich
eCCanD8cVze0iSX1x9u9qODszDpuuZdM+mKBsQJRFs3scqykU4qg81/Dy+IshDzFlnJIK7qciKij
R8bGt6AIdCDTNMgBZ3MrJ5J7owp5pVQaPCjrZnP2zyfEj5WqBXH6gDiVLrYdsArp/093PBuAEcjt
BUeAEd4Tv8qtpQsXwZYWVPM4ZUWNFG+ccvxWK+YUmfe91EXsNk96b9E6kkm+NjGdPz+Yw5R8cjNv
HJneBvya5DdVxf8UCK3RODz7TJTkgrX1wnoAcBIFp5eYqhn1HtZKO43oFtCHyIkvtEG/ujnXe8Bx
MvD21oHmBKaz0qpxENhLHCIUBwP8xNzSXz0okQo4KhWMwuKNsUbMycNn2F6IkLRnu8tSkh0hmm1a
vNrXLLxHPmI5IYvRF/B4g58JHA+HscUMP8s7mtyB9X4f9sUKaJXAntRO0ceF7cY+8g00elfQBp21
Pg2JOuhxppUBL6B+wgTfGRNM3JoS6bUkLjxCJtIAZ9QYcxieLAkRVROfLFoOjWSH0uMEZEBNtJCS
zdYxF48hGNJp2tMeJlzKYqC4lJhACeRCyk6+doYjz+kPTUDb6LVvJ2RZNwXAHoVvuohvkVMUrJ8U
W+bqY9LQ4lUuykpa3JlyUciwGTa144rcPhaFHqorEFD07eTcVidupEtwfJXeDrxTNosj+qHGLcgm
HFqi4oscH7f6+BK+zTSHhXbjEDCaq/CTdmsu4XjGNXATWWf5I/xD0e26EgvfOeh4SDrgBpWHxFTS
qCLtGB9JE9mkXxn9rAEIKQ34LXrbM6aL6Qo8IdoabajcLNyys7uDTLIraYQmXNWnBDOwovjqhDKq
1E0DqmYwii52MF52BZQkFkAuSEqkcrpikMv6kREHD00W4lFNceFQmow1QKgvINxYKcrkBrRqNDvV
t5z7XMTYJnAKGvIsIoMgTVxahQpHo1SEPsNPik2S3ZnYHiBfE5kop2+rT/LZOa75Nno4VX9FZSHE
mwFgIjW2cEcXFkxl/P0UaUA2w0Rtc2Vj48ZlecI5JbkWRmEvtAowCQs3RYVLFZUctw4pCu/Sx0Qi
QpSpswgs26j93sexdpmufz2gvjDhXYZGn88grAPxun5dxUBcgj8+MaXZlXJktkSXc6BdRSq8/1/n
utDl7yvPkVECPy2nIptbAMmSqpyiKAh1REz7hk0xs3/PwA5UBCBuv7RJ0EQOHiXE95c/yPH1XDMm
5nIc6rgC7RXXCAvQOKAZOwBrjWSeX9pdVbL7Ee40njfgmV+LknRNLuEcxETvycGE0hnxMq6q+u5K
Y9Jvhhr76kXtyFTV7L0D7MjgmuTxoEbSnwee7oID9kgkRSge3lGCq/JS3iXM7akd1vmVSUZVF6NT
QaAm0UMDgw5RiObqP4N14UtmBRyO29ZpnloKClJbdhiOFAs2LhIwoQwiXdZPoWiKcg5YK9zhHZwU
qiKNUFXqCrIHbbyxbHPK4x9uEJVBI8706N6zm1dDGKaF5uKa2vCjv8vGPu7R48vaj3dfQ2KGwkqt
CVGyVAOO735um7DFdmcGMVg+k8AsuvWLqXkzE+8lPzidiceUs0srpcnJbpg9n9WacgbROt00l/l3
XQ1J1mJN/XAaml+3fEEeCKUBHK0T4+CMhQ2OsOf4j8nOg4sJy5QtKsabQ/mwW1NikvpQPiTMR06z
4YH3Dnw+cR6q0GRCld4sF8cFVX4zjWAre2/jmszhzRn3RS4eDKh8ioO5VXCcuYhUYX45lwcAXXwa
HBE8WB2dQePPRMFefLxKYVeiciFO5Vag3wf28ON/brW+AscTE8doxRCXqjtBCEnepSgKC2jWuaOk
kGfkfVb55bMRYn4cj/3AV/acDA0QEkQ3jLk7IzXRQBdMmBhudbMxnfPdryx7c014dhKUjTofWL1q
8/76GHfj4MYI6+v+32AGcLPY85nWOujsmB1AlF/3iLarwMomstrd6YtYD77DHxCMjCI7WE5gZi9i
0TLJDa+0KV6YmPiRlVgAFnM80iu2nm92ez/ILlq8J3XWDm5vpP0jj07V/R3ot8Y7hvSBCXlU32my
F4ZJSf2aEFXcoGKa329tosFZvB1lYBrvEOeutJmw4HuCzMEWp66KkEgJpQT7GixnPzGoyHVND7f4
DgwH8YKbt4V9skFePS9SSYhILipBe4Dx6AYNDaoi3S9jD5PV4n7b2HTwJCylJJcYhOr14Oun2hNY
6z4GP0tkZ665wfZJi8F9RM2EZFop5tTd+dXoSdoTp9uqpeNM6fGlrPSQmRbBWxGF1CFLohHoeRNm
ZLOxBiIrpkxXTCXqmHdVw2J3xJWIEfYI6+BqK7MZ/dkCBRHeOBU0H0T8oLgquiPi4hbLi+WHUhjB
HJ8l/9ogWs7au2sBaouK3+3IYWHsIozbKNeVpKW9PE9lsKKIzfZYDXN93Cq6rUYG61lG5kzNqD49
P0upgvuNcy6XOKbgp2Y+voflH9YdXZYoIEREm8Wd/8jkLo+wY56R4RgJKrDtTDKW0FvBpOeJpxP9
Yp610KiEYhCP0QHxNIPiuukDXuBsPQ8VDKsQaPAxZ2NDnJNtVdMlrvWnsTXhPldMk8OIRVf+i16N
9lemip+qOaqbzWB3JMvSHy8zqvxuy9Azce1sn02xoFzVZCLQsIu2VWMAFJ5G96dqMvGHY/74C5eA
Deb4jTgV15ax5GLwud5AN44VD30/mWPxLXJJvQ9pHPRDnj2/bSGO63VS9dC6aFLZT8Wd0iFPhscD
gl8j3gob+W3N4mYAio0FUY6SI5ND/OnfFMV2Jrt9mFQaoLHGQz6ikuOab+/LzJ5uu3FDMsTSgwam
yamzIT52wWa7/MlYYp5/yTXqFUUeR45vablqhulltKQJ1NR5rGZHhvN5IuIilEM696vIEzfZ95jf
S6LDYmlmCw3dvx8HzthwiMPS/oM7F/8kgbLtucTv6Vyuln1Q4vnOgOiyF0LAYAvOxJcQIp6Zkb3H
L6CCLvUjbdyaBT8TspgXRSWh/Wj6SSCSrHZXD7XdaibQL5VGF9xZZGbtwQapndq92R6tK4KHnmvs
pTpYPVKKkk2lWeJqb3ZQBQNLRd9PWk8w7x5ws930rvFHEs37h7T4i7xhONB4JyjP0Z8GSn6wg8r1
B1MCWoAmrEn3oqVOy8+1BTF2nsT0g7RgxluRFE1teSKKdd4CDbWyrrWVcvPU+TEcBkHTShdAboDr
9/8IUmhaElU10MqGlDjGFE/ZlXuxbgD2WKW8CNLmXM2CI2kGS13gwxIgFzgDhb0U/ZqrG8lwlQXE
OcDQ1NwXbQiNkBVY2bT23MiaqgP46MDbbQYtj2zJbDJeLmoHQCT51WCp53qavQs7fgktXqZD9I4F
kHbO2vRqH6S1uINMb2v1WBwpxW6lvOe/JmlZcHX99Q9Z3ngUl/zHXwpOkU/dOAuHr+QaZg9AwCZD
lxdLLEaZcfxNNlpu38nQIKAwMl6n1QAFvmjUG7aP0DTk5ctKScFQw60PQhaPSQ34ul6/QOTpk5mE
SCNFTr4NmXtZy/5HHDEJ36yCcAs7eoRY/PQ4HHV/SnSaJetjjCsd1ObjYSll8nePvzXZqF23nvKu
lFw3Xyx/+YGCkDyCVVu+uRhl4Nua6vnjGnZE1vQbwX5UcbbyVPPjSz4fQYipmb/cRfjHZntzXWI+
J3djUtTn9UZq78bWk3vT961zWLPisqD+RtqTJdv5P+oiefBttLXMPjY8In6K5aFagGO353JHEuEX
143ymRlLf01TxHsLc+4b+bI4yx54BBSiqfuOOP2O9eS9BtsArcxOGw9JYkDS76E60mMQZjYS8Z2r
Jqpsps8QT5xFwynxOQHnUKzAsreZ/ZWaNIgWb42z0BJ4PDZGehWBZGDxHl7VtViSQwTGXFrBkPvt
izGIkdfRatM29PINlEw7w6PDw4sttnkHRrNf+2+PVGzWStlJ3Y6OpoeY/QXcCyAxQ4rmVg6hB3wX
oBKBt7f8DjDmKeU05EfDHTg8l0JO0XaGzkK+wgSKHCkcBjG/opBMiZkYZzb7Q3Zrmb8q6Fw1CA+P
gXx7leoOFrBIh8FGaA3ToNODuxkEbfzpob1msRl2IeTGeaoMsQ/PxOPQvg7VVGSVLfVweZ+cyr+d
htUukYPjjfC90HQft+fsxI38bhWDsz/2d1QWHkJbEnC1AQ/42Lh2r9ilv8Qz6UxJT5bZmpvcHSSK
lbAdO8/5TF0o4nl65KKGL0pDUvVYi1HCmCTMWIB+Y/RL3gHslGJ3T95bNeAD9xtfQyTW5ue+X5zW
qvnEjvO5LYTIxBVpBAFSpJXU4aRouD1UV10TK3DQsPEE+Y1A0BHTz1Jl5xswkHSUYQWnYz1rbBjA
ZaGSMiEmSclFdbtUeirkdkDWTqSwWi6r6vUXYcXKqiC7YGVUDMo+lCHC+ODhCBKjXjBL2MizqIOi
uTC0fwdwv2CLM/KyEBbQNXLuPnyZLXV8q3knMM720vrWVxCJMIVCEQSGM2NPYa7ZRgzoWvY3NKyh
9zbC5bH35FIApuNtX/jJ5oUBtbd97CRmv1rVg+IM4d4uvBjnYSA53A3QfPcDVQfLXDjvHRmvi548
gRyCZxQjGDfQFFt1aqT/E8eGUgIXPS3PhPhSjuw9VgcPLFm4TD3A5fQ+Pq3HWGoVjY6tZuvrtQz6
80b5zGYZoveiz7UJSiAqI5KHh7/XyhpA0UvPu1JfQj7v5mEWPDqyXK8VkFubDIhuO9fhkZ8nACJu
9Gv11IcOItJvvUE8cJTQkIL36ChNxOxl1Nt2TJOc1yg/VmIIjnJXSDxxxqrBOHYz5J04wrZVWYai
hL/Hp+yt0fMvBv5mUubGER1TdBA5IDnXiWDpy+ruu1DD98dlyer93UbyFVBhFKaeVvCCdYG7MoEj
6zHDN0MxOvLIeCTckryJeQV8Q8S1QQ0xV8j2Q9VanCsWmZReUImKZ37/KzUng3AFaLgcaiJNTsMl
3e0SFEXcV8wuqXgjNu3g158nQIZ+k5vz6BWx+p5YT1FT5Gu1iTgMCe0Shl5KdXTjjsVS7lJUyTa1
EmjaeqOTJnjV9kjaHCeXkE53jy2u5nxzoZ1mRe2hvenkDqgV2yAanlMZOUrBsRb6gmlggrlTX7P/
90x2ygD+T6SqW4IjwUzfLWuDfi87f/86Pu9xaG6N+quMyL69Df9sh43kco1087+G2wIpL128Eefo
F3mIWOQPYXLKx+SjSNeOrdYx3xh7sss1ffQXeLA8tCVyfxCXvaW4Ydd35rOE5yru78EATNR1IuGZ
K7YRMPzxSF5r1baSsp2hMeHW3JzTDSmqDcLqusxJZxyAJb+aVZjpZ2KGbmFpI5nQGkFMaew3R4nM
+ZYZ4LNfVrTivISGPJkTxWuE7juesohSZSxeVrPoaDghj8Tv420dy9EENk38doKc58cCexZh3OWf
CNBfzIke8rmZXeDLluACHDy+fDVAF5yMFzemXrx2SGqoqwG8L+lANJBUpZDhPSHXyJAfbMySl/u6
stXPaiyDljpoRubyNuVR35W8CU/tyApiJE8fTQfV25CRPLvonamJA/k627lVhG+AfUdfBGisIn2D
oBhmGvmS3HvbmfYSPF7gQoCv49Q8pvYjHldl57fGu0/krJaP8UILTyss2mOx2HmidMgFgt7g2NGe
wv71CboxHlU4I3Kx7KAkiS0kr63DHqRY2vNs5CcCtmfqEHwOkqG06LZT+A/rlrwRMYRR/1d4/wcj
Af5HXA1lDn3VjZDppNnk4NGjfI9GdnlgrHMidiol28swd5T2/oiVe7jYiiQA0mr9bCeP3MXfmFVe
LetDktmMprWkNCh/6WERYqL7pVDm5J5BHLe1mQAdupBk1OYh7WkdvV/PuqKhLcFfF0TM6RxyQXZy
rP7Fb9zTdwFxiS3msCCK5AivT9PwmQyzUH4GwuO2/ul+TR/ChsE/L5eQ62dhvkvmjhxov1gzRg0M
7Lmc+tiivyH9JXR+WHf+2fSy+tkcL5eDEHpyFgcOpawo7Q7Z1NlTCTu+uQRfd/Cf3Qqnav3bZPrU
VpXDbuQ1rcnlWiLAwYTf+PEXmGn0JHAcQwv7aK29PdoTEPXxHCEcBkINxbBZmJ9Tf12mv2LQGR/D
zLWyJ78gnLFRx0U3uTH5BJVChx7As0QMzXIm0YVbBnj0iZbKpackjCBUTbSd+qBO02y0Yzb52I7+
sfhPM2Q64j/OJIF4eFt4dp5L89bpp5WANTacuB/l4b9W07ccKMnHUCs0T+6H7B8CT35h6Mr3FHGs
FR89pG68pX3gsXb1LYOgyY6cpUyke4TxsXWFMT92ZETRcyFqqzJswVpXBSj9gyznDc3oPE82eO+y
DfuonPAClIgVxS8Jzy8Iehg7HdfCKc92TmMcN4cca5Jt41nyD9DrWHlhch9y4YsnXw2pVfRIiPI1
PxUrM7G/0ZroO+s00WqeJSuhXSs2SbEMgo1P7wIYqiXlVGDcfcQhbf0eR61Cu5orkrENN6k7ElQ4
MsW+oDfW2IahCE5S3LNKb+y5rGS0XVLL4voeD/kGBvQtu1ko7hFXhKBZn60mZid0/zfkC0vB1CSg
EtypMuJ+jfZfOok5AZfs+1BrJK20Te5VgLBx/U0bRie1u7ZRmJC3Dbk1zK6Bw4BOD0rpyUnTD4/9
4ES+D6lF+ljRpGZRNMQSG2rUDpJEFNiI8ys/1EeBpxFxf8Aqd1enAB2RRTLlT2KEiup2BALhZGOa
D0V7AZfeL5SU3SJpCVtD2nf+UPoeRvq7vjecsGssMGzTkIo45z5/MglQaSK88blWLUVmdxP325Hy
o/svqm/Boz5TKxD3ML1mK9ujpYDpUggw1RLlLSm0aHNXA8Jxqo+vNngBKpwyOp3vjvR2V816JIbN
hsqUCjRxrbqmYkTKDkjtFjN5+Df96zSRYyU0F58jIlh0iWlMGKMEZ+SGx3kLeMJyzJN1jlfB++bV
VaPTg4IuE1bDgZJls7MPeDPdmvlkNUUJVYBb6aalV6IipNyk72t0Qrc8mq/RwHATbSnefEEH/K7e
mcWC8Vo3mm72saywNdcJwVj+4A8qC/ZOYbrxU0ftt1uJRWKnLO6WaKxzEgBmjKhAjcCA24rviVPu
n17t6JXLjrMu0i9c9T+JT8trqpjn9Xz2gy2jSci61gbIHbil+YRW+HRF+c8ht9SlMD5JK1Ud3c7i
Nqu+VQLbW0+1vvowApCw4sLESd9VQyre59eIV8wlsWhdrAA2NX8cFcCPQoYnswWFjnG/gb6gFNOJ
zHjQW0XRaOh/wbSC9tO8dbv9qtLWdClQcGd9MP0BTgylfE6MOsNYvmGYYEpNPFFoWjkOCteiBzgb
FdTRYeabKnC3eXTgirNusfgGGYt/V5zNWJe0SltpGfxOfVmF8UzjNvwPyFW/m37lSMkp2T7ZdEG+
D0Z0gFCmDSbKr8CoA+X534uDokfVQvjuqvZMm7h3ZSSr6mkTJpN+0QkEr8i9Qn+bRX5YZxgyH1kw
w7U9Q1usRjyblMVU87fNKQ1R+IfmNcvGcHX3eAwp/LcQeeI9p/Rt45ajmOveDCbOfMg1MUVAG/2K
r3Lt75qq1nXzyrM25GxR0v5rORPDSu4cSHQbbegN2gPPzFH3+iHpl06yAb89GAr98xhUOBrup1gi
n0pcB6Z9AZXZyLMVXmvHgyxGr1MboR2zStDJss83x2Q+Hqf2+fwJc1CzpSBgplSx31isMXLxG8n7
B6FH8q59xxkBm/kUnxTB4RTcf1vuzZqfoKm+sSoOtlUN9DHYmAlZKlHSVoXBJOG+xaClO8FhwBTD
J2VKqQAa/x9OUdGzarDg9p3D9GFtyFjw+QjIGF3GYUyMxyzlagk8ZGctZ0S92Pitl/O4Y0aoFzDM
n+8PvFL/EDXJmeNGgWdO2MrzJGYsWAecVG1d6Gj+Pcx5oHhi1FGV0zRNrbbII+OUmOjJ9J8/uzjH
KXvqDQe0N3ZrBuN20PKs9mAlbiV4rAbrB9RpauvxGJaRd8Cgh5lmzSJi8XEf4a7pz3Sc0RGuPYPO
DagCQiDQwiwLd9Maph/ma0sQfDwOxEgmXUHw5kCLFHQKswrA/xUUGPkBnkaD30SdCri5ELE42TA1
ptH2h17VTD9spUyysl7f1qbyrRvWDTItoxkeZTRthtL30KdbKkRThxHfRWgBHAKJYUBETRnIgj0m
DOVeqQlXCxQFWwJLuytmksGjBT/vyaTVr9RF0j14941ML1gWq/f9zMPuJnQByyyobY4a9mzcjIBH
QXAT5HjrMN1qfGKILR0h6gcAPx2zCunmkX59Iphzt4uMFSjV7sCre9g8n95FztBMOZmTC18Bwrrb
z1EbOYuTmOwxmnwpoWJy/8ZezjRxuQ3QuvCX19IEGHb60pwDZrz0O4WOfeTY6EXIE0e8dwoSFAnD
4e7o72HSKRD2/tBALC+MdPu1GvzlBXGjs6f8sIeAO8Wa/PkfULgBbLjvwTGc2Yi1tm8kaPYjNuIP
LnC0/tmC2KpjRUcdsumHgTV/6XgLZPuqBJ6FVNiki8JCM+QqxjkzU/OWKk31Si5OO84xzaWaqSOG
17RRlv09CFqrRbi/yzePCGeK7cbNWGz54OJ/jrJ3WpOIIX8sbySR84+oruLFwp2fw86+zhkydo8Q
/TO8Wf4NR8AHxQKbUoJD3k6WGrhBvUYTbd76/cQBP0zMzjoxQeHKkItZ1dnhKhhiF5vKLwXBT4lG
ZlFHoNlvpisp0LX+03tABjmr7XyNH4uKulpw7MftRBxyuC3yBKbYVn1lt0rXqvsp7FbxD609BJlG
OILKvlRMbPbGIlfNCyZlFx1uSeBGg72OlXf76ph+3rbRlU1aCSBOWPehWV+86OH2j4gTwFR+yEm4
MtATgoFklmBXUdPXctAYsC06lv1/o41LO79PHzb6VBCZDX+VrIbfVdhrel3bhOYoTlbCG0h53+uu
6W97Md/4ViURb6AXmjH7DDdUvthCaU0Zf3PqeAU1MnSpsxvXtfM//efYMY/QCLIjT6MfwedC6Dpl
mnNcOxfcXfXhZjRozvXB8NX5MJB5wNxvbP+C0zy8OPAW3e0ZROcO3BIom8yAKWRmgRRNs4DjZ7Lb
DeCvMyZBHmRgyA0YQO9i1DOk3fQm5PLNQBFqP8+NjQxB91c9EneVhhy80ovZj7yxywTl6kS+L03C
4iK4qBs9MJiqwxDlMnAGwBVbGeuhBxxt+B8M9cUwjfNsnQmxQW+dPSS0RPPP77Z/H45IaPUx4KmV
POShZt9ws8cUb6RhEi5nIqaEsiiIH47UFw5hmp6WvzaTYTTfjw/jwc3fLO9W3OK9pRtWCrugJs2U
+V2TWagirj18jQCS4XLJM+8pnGjFMskblM5QQEpPMdRpFFq5DSjua1Nhtq20VecKSqcypC7IoJOK
Z7UAwotOXtqHnbTgnvbJMS8BJEk7ACog8fInYP+4WbH4QdQuHDDgPLGcuJFWrHhbEg0LEwrVB6Ux
OPO4CFHCn858matQlH0wOOYYmG99Kn5OmvsM/8L/j+dYiOoSRlHIGfQiMsCKkykXx1dGkB91NEot
LN2OyWYfRHbKKSw0mwFuQSiTdllTxCbJCwy4Kq7d0hbNr8k/9hsSz5qa6anj7/21/c/FJObYMZ4p
K58Oln6ABYo4Im0kRK8CIK9bOvz5gjcQpSRRyM1vkPbV9KglJzhSR0PZelUQ7e80KzGn6mQiTbGo
YZOfWVJS/4rVdTDsWklRqGOsgsXwzgDREFW/RdiXcxCgdjXQVXIt2VleXmN0hJc75kkoN4k6oBeF
BijVBTSvmvUFuYMOUlOegYx1Sx3HK/83syUtT7GkvVnjJxK/lq/SJtqzTzobR6tRb+0p/5fEOG1n
OhWs5Wor3xtHYYAPPnvvA4w3WXhvqV+E3ypmkB4Z/8pDNKFLSPpZLddq1epkjOe0OyFam9Iz24nH
2YI49S58pXtITDAhe4XqPQzfTOnejcC5Fjo2r3HTML4vdjMrHAG6qDRx2PCky8M4cM9NL2jM97bH
tHmdD0ymBY2/tv+iFj3BFywRjnbSSJiUNg7VavUtnboAgxFQ0/J5pIePqYt1dqiqLo1+uF8v3MpF
21RqrGPGecqAjoM6fBiisfPzIxmT4QSev9f5hxXMatz0Nr0TZJ2Y3jvEfQ11ksTVHmxlIrShlT4F
vpoaeapMunBocJsAM6M7obg9Yw3u5BSNzdxDcxET0AcGZ2wNpx26/8D8PTdDE7K5X9SH3cwhgvJG
dVTA1QwTJq9bse9aI4TN+g5ub8pK8uRqJW8SUelQ4IV2y5y93pA36wYQ6PARbahC42Ce6HjBNNgg
eoufF9ZPx4NhvmwTTaQr9l9+d4iqpHVuWrrgBrC0+WxMpJZgEL5wY+2BYQAu2CJOMEaKawgPQlCg
b1XTSg1BK2HvtgfjGSGESwTI+dEpkPUhofMYumG3g6gdP6dYYmlFe//jP0iEzO3WaFvgjVk107Vx
1McEsv3PUyNNPIK8PS+8Bh2Cm/OUK2cOkQXQi7wE5+RuIKYKlMyiG+g7ADhd1cZkvn436wOSgg0E
vLOeMr/os9GwuFabu7eVkZ4HTpdQd0KBe7q5tSQp+dwVr3uaqQrM3Io7uBz430eXAZqTAhzNrYM2
ClZ8pSg2J1RUpjPKfuGd5lB2PrhQQk4MNRRtZSrIpc/+N63DpKbhms10RXHn6vzO/dWwnGG2wOJD
OuttgTc8ZbNYv6aO+0VSEWjRjjYPSSKMzP/p2DIDIIkmGJsWftRzKAYgvWbfDTtel6v6QAy1DbHJ
RWkZ8v48GL5Kc6nwWIUwpySlT6dfRxkTwKNmXYz2VukWTmK6ENkzMS+u4aMQ6BWeQrhWdqh0E4nn
MTiZ7hKqyVPWsNTpbCjFFWuXksvx4tuKrYksyd7T5tQ1QDI5OYFLd7l9Ri8uoDNWGlwHjkRpttBI
eFVcrNajGPEqAwJIAb5/CKAhSbFYSvhfH28L8q+BJke3jVlcG76f+o98DJmvD2ofyfkhia/YyxI3
bZth4hmBwMCY2AjszAKTNihgVP96WIqgZ/RnF8hGzb1eLXSEVER0dQuPQ6djCsQ4kWHU4XARY7VL
mnlteml+VyVOi6mgEy97HwuyHNWOKRdk0cmn3PrckWk5R0nAEodKWYOdPCd8Jocc6+qjJMKncdx0
TFW18m/Zmbah+0rx4c7WbO3GLXahK3T+gWwrFXfKyWtRzMaWBwE3GnQitD6XeGnDwbWEtr4kFkpG
SozlWz7n1pPmMaV+dMXE06BfKfi78Qr8rqunUgrTYKFGd4CR6s9cIDU3KV20z52QHWbnuAwisQvF
Fgl/NjU0bX4TjAGpCG9gzSDoaBxs+hLLdVYY73QVgM4Dopc2pZcOhxbrPh0/Us5bjp/dkH4FU0LK
E9oXUhXjU0iv/nwP/j7M5J50iZGeej7OywN4PGoF31+Cx1gNqhyQ4ZhqmL3CK766YCfoaQeTpd2D
aZoRDIxNFaKvdDikWvhQY/gkGhy5N/McdkVaGHJCc6MXtgCYJ2ky/L26pMHDARTif1WfyTefkM0B
f2tFtaDMqgTsjo4ql6lICzZAA4srpOfICSJEpWXL5HB4I+1ZhbYu8G2HXZxShBuFCeR4RXsHn5Mu
60yUPF/NgPomseWMkOVwKNVKqPZudGZ9Crf8RV7c1OikiE51FQzSaTHOcJVeVrLzOWwVWoR/nz8i
rLHjKNbUGQw9BQj3yh6w0YsKWrsi2URFhoX/dftldW63LoRpCcngg9dKwbE+K7WcleguMlRzClEJ
M2oG9eZh0Z529d9skc0OGMmW3oH8KHKqPYaRS/oCVQYZiGONTxSlCdG6jkCwwI68LRZimEfp5v/n
WcwoKfbDaVqSJKR5vFDId9R8VUpHe+djQnNhx0iH2nkg99DXP083FTCj3+bKI9fArcjBNwTbWbac
hivzFeUM7rD+tFzNDhGiwjEWUCGZ0vbiOXMoy5Gu6Ltfl8EvuYBPdlS+dz1HQ7myBx7hmh8V+6MP
NNs9avEM+H29rGGIsCpwkyByy5+CbtCiD2GhxjX93nZl26eT579CmC7lKlaAdD1plrVilG+l+dv4
7aizc4qcZRysB+SB6NgO79KI4rnOhA5CfTPW8NL9yC2GyofLFpx8/o+OE3O/wILssFN6R5Z0hb8S
HpMnBE2daNYTePCWcz4y49IV3iubtJV566WQN2nn3CQMvlFog5IzqxTSUpleA3AHeZa2Fnt2EIRS
bNmFu0IzMdqONprEAomrwUna7Af0MPLILeo1+gb/tuiPlS43CazOGgFBiDs4c3z3YEOYz6igqCWk
mYymPKjArdjkFbRIcjEXVWYLiyF3nwRefyAikya2yfxhoC/hbtRyhxLkPK6igittntkbtMPI+Jgn
wnf4NGc+ZxYujFTPGLNIHp3iC0TeND7caAL06bUXv2pVjIo5nsqvpBBrbvdwEdAEa+G9CUmfIJFQ
NW1S/nbunfCu8R2NGXwIXuz7rUt7LD6q8zcM+tgPRQAiZ9F7BPDZzVbJ3PbwFwwcCcKNvZcjP2Ni
eZzTaQ3D/tJQG+/IlHbnqInD8ycSOmdXTiVY21aWTuZb97LvQnX+lzv7/Px0wQOkHG0PjjR8NOFg
Yql0l9upw85Sa28XJ+tvmuT9PvLfG8ZAADg8PXrz9qcqeabteTui6xQeHmEwI6Gy/BQbWoW1Rp1L
t0pZtm4A0ESPQEfPjioyBLXchbBRWj5Py499SbMc10EOIcp/c9hnn2v/ofDeoo5cnXAPCqd/dFOr
jlHZb09OY/PIj2dwNjJZ6qNv64wLUhdAiAK6dG4ozbkNS+JzlN1W23w9nGcoaDLTYCO9iDUkstgJ
g8x+OHxkcmPrV+Ri3Tyx8v6ammmzEB8Y+9/Wudb20O/NQGeVWuZabRRYW/mrX2/TBm+XWceoqL/Z
0BBew0UhmHhAT5d5uvhH0m30ilfSX0KBG07oVu3N36kS/nS6JKWOL8XTp3Mr8Ky8FXGd8q3rzVr6
LCYXFDwTFVki9yoGb0O1M5lyCaLb6JMfax4DorwgQ6bXxKnF1Ak1dIXIUllYfq0Qn97bV5labUxz
B+AKXlNV2qGzcQmqaBqw/FnmB9t7vcoudRbGbfdilZoS1IjW/agrCusnnq/GM/GCiOlag/Cnbrde
HbtUTMxX7q2AFvn3f2CEZJjheXXCj/Bnv0Xa1MmtShCgfXC80dQThgaKCOIaVIuHMJGbcQXR8hPG
nKWb9R2S/hKmtX/WSBiYpSJ+wB+d7IpEGuQhAZDbCiVCZEPtSz60t7H4Dz1uGmZMlD0cOkMQNywZ
wqddzU8T8TAzjvxo+QBYl/A/rQyv1nZ4aYywcfCxFg/Vf88rfmSe7zWIlynBShTxU8GOq62+GYtk
bPhzQSYY0eg0O+6PLX+QUFKZCmBuablsz7/EsMKsVyAdhryeyKz8ns+HIr4OiszdimK3KT1VXjHI
nDJilBl9oVtJ9YgtZBXKkCxNmZnikMNv4PuxfHnMvSF3QSR6kZOtPnpgDs6dSFFqa/QONMQUTVmO
lmrWvgHECUQi+QZKmzAqO4jtnVidD08AY4GrTd/gPyHDnoNAP94V0BvkCo2VTD4hrDh+R+MihO+R
Oa+4oALrYo2osT/6oZD5FMHr90NplAc1MMOjHrpXWD4Ygn2UIr8D7OHaWLzNVs57RsGJHOe/LyZi
rmJB0cDtzkAMuy6uu+9l/HQFjHJx6dxJDphCyMGbgHikl10/PUNEZsZPjwuL+4COyo2+w0BkIWKr
IU/LtKgEYR54KqCyCsEquQW/g+43LEAVUB1c+X6ewR/E++UqBUfuSx60pwpuVqCZSyLCi+fGRF9t
ega/Y/MLVkTmJ7/bVSMDvB16rw2mkbyiEqO0k/PPczFXZ32+ZGIR60/swwp2OooNo3QyTdMv62Hc
9skFz2DTkVSFjqW6i2AResUjodQkX7KM1OpaF27kpkfJ5KYEW+dSy5+hK/Tvofzvj0iwgtGj73t+
Uu+djYZN0OfJpGwswz2wd3TsSPzD3Ln898ZmNXhNK1QXp7810+g58x4bYCekTINB/JFeeVbtSF3S
Wkk/SupSp1XmfAtKI9fQVZslKn5dVaI57+UrTNuEgIwJMZYkaSUcv6zoHapX5l1PVYnVQR23OSmb
JIplvkG1PBuTElgkoDR7qdhO1m8NuNaJJLJw9Ri0/349QIFhsvaK1Tl71553H2PD/NDcTCCSOhia
NADouyN9o5545KGTKXovGkcOCjUB3CvcENO5FPavkZqr2jXqvcP8cgAqRlhyk7wMB6r5RnT0wLI4
yFQthwdtY5N1jX5awvsFJg0hFwxwgdIvOqa9n9PvvWkilpy6CThOuPE8LpxcSEwYvsxImrfug7zc
iFzsvfQyeJp+or49Jd+BjPX8Uw/4JyV40RE6Z7KaKEs54pwHsMH9xR5NpdTiZZMKmYNE6knX9OA9
0jqUZHhrj2mhRjSm92qPN1kzgAxkllOXudqzs+jMpgaGUQe6GnrRRbPKrLD/iCRQ3yjythABQ3u5
bNkedmtd0mA2Ywv34IxyLba+7LU0ijx8xp8TMSlUNNTIdude4g7p2KkABe6RZkGUI3RAnhTXUqju
gocfmL/cNt4C17e9bxsL7xdc9Ehc6Oq8cPNNjW345/kQVMnJhblGFYXl6iI5u4EMiMXnSnwshMOf
UB1fDr6nFrEe9/I43YdTqxUQ5gt+5f9Gz5iSn/j1QXfV/iDRFy/JUaMWiqiLQwfgq6bE1yHnT3Qi
44veqMYLFFduLa/ERGMM9b2I7QGxxNs5xCYAXK1BpumMeqskZIr//hJ9/b+CozPbxeYAi1foItfQ
6kek9KmWUImDuICuOsIjdlaYr4MFzHAQoi2SBPcEjRP9XBySDAHCVLdryCNKPTzYCoAbofgryUJa
4xhJM6aifwMsxIOpuIMZ2+NFmqoOsTMUARWKSGaeaRzFBuUS6qSGbV8MK+E5N3m10lIAdmDhFGnU
xH6N6dq/ZL1rDnRXq/uqgBWbUPBqeGMNmiUifbGc3Mwxwg7Kygq4xJr88R4Vo3kma7MRiXJjrNbJ
27SS3nn72IR+Iun+DJ9Am4sB+MIA9li8vH6VPD9GWZNBH7iiKrhMr9scTHiGVDeYua7sDB7m+LBV
nutJXt0PuMpA/9VFj84WD48VQyj2HPeJvWGwJV0/OBaTiHg6WDJ/rGO90KgSu9vcZ0HgsITF2BF8
PQriaVQBSyrXRDfBBGw5WlRYKurp2a7e4Mkn/Kh8ONuFg3uHxqm1mFReIYUK8Nb0e/bKavnPzSE2
9zCcQp/MiAJNymnnMRCDL/KQRrTaFTDswsrN9yEG8ZS5K0GRrA0K89QdHiwzIcIX3tNRlUP7E412
8WqjowXOm8QH/KGbGeC6Rk0EkGvsTbsVc4WtX/OViJDr3rHfLdUG/u4VDKUbSj+2wsNa0TJDdEQC
bIFPLIaChQHzN5NfriYNeXwuorFppNaotZukZDkMuRkLXG7qamMoSmBKHwBhVplQQeSJTrV34jz4
4SF9X2h9E0d2pCKTsszVI5Dk5O9bWxi2rnOWk6UO5o+3WQIJRsaQmY8UMoYpvCEnQUdfVB20T7Ka
wXg6BtQGiaY2FC6o5xnMI3Z4ci+M63qg8ujQEn+o6eVa2YvooS4K/DN7CQR3NcynexGEs5CNsJP6
C4m5HqZ1qjf9CsnpglTwKUyav7pG/FyN1MjeI48P/zmtc4tCDIZKm0bvkiM/Y/DXSY9VlFhJBfu1
35QG2eOIJR8VDFJBddl6S34ToT4eRePCW287v4ENTf2PgviKc6NmqHicQk5D/syn/cPVFQmt+x08
MYfgOZ44kUnWzf2fbjILktxyO1b8wwEMo7uvvOW5PBvYydyiDriIcNMgtvYs+oULel6GLeY9iL0H
YK040K2vLXBO4dQITV7QDODak4ALcfYh+YbJIYputOZyr46IiCUaZh5S5qECGKHqO7chbyPZq1u/
2eNEDqrh7WQEI9rb+AKSnmG4oF2z2zaVHQNtz5CIMuZxTduVKzJ45yqQhAR4Xqg4OgsATj2i75EY
oMMv08LPdcCUvv+oIkFXbYFXmmDUlCaCqMMfcD00mfLtOLf2YVzeWtowht0uuPguga8zavx9Joru
Lqg2RqKSRvGgLT5em5m562nCKFqfipcKTRwllfnVsiUf8wVEwglxg+hfu/SZorAAorpOdp7Q+iqr
wWzIU41tYCylsVAPmkSiO3sLtP+80SKHAUqEIJ3c2dDowcIx3g8lbR7jKVVqdhLlXVB8Ax2ziw3+
uN9E8Fm/wgCrvz+0/pNwrWKhQQqKO8kib6UDmyVD9EQbaAvIFQtcl4Vgu40jW5F3yPpNAYWQgkhs
4fimw5HmE80rsvF3LbWcHqMqGch/kNvMvjxUk6UoMSJLTdDAuv3YeljCagpjY2FjEYqDQmfbJ0IC
kN+PAGjWaZsZz/JokfgPPEtaBThI2AUgfz224jHEna4dENqJy2/7/Bq/H0dSXPGGdtDHIXEGDrqY
+OMA850vff85L2AejuoG/aPIYcOf1YYNMFwjVsuuIyLoBoJNSsyMvt5X9WNmRr71nPekuJvrIywe
q7J6DFuZWPAG6Z5Z0U42+1LLe9M3D+zxRsOsuKxsgtbMT5sGpl+a4ZUP0HBtV4MIVWO1T93PpUNP
2dWhID7KkvzyMu0XgJZzMQtSD9cClXXafJyV2MjkdBLCpJWvlnWRoofVTdAr0Vn4FlBmV59wp53Y
GASg3JlvrLj9DmvfDWmwljHs1cfbR192NuvTiwBTbxYmprUGI9rGd8vy4xqRQpdskhp70vWnV89z
B8gK96846qpJS2EcCPYcibCwexdgTBgS6LGAtuwUUmgzz3/UclT5+iR4Qixe+386EsNiY+OrM/kq
fVaQJX1vt3XBUNy4jTepqNMRrPrlJ3Y0lungJ5ogANpyN18v4Uj4/w/YLTIo1laESatRc9vsAqLz
ZLyd9dTAce4PVRD+YGE5HwfP8ukshjY/oJEvvNK7ICwlgKsda9QXul0KRMwht3kpPeyAPVuM3TLn
2d9bQD4ISMHslQes5g3EO6G8XtylsypDnlmQGaK1dulRIFgh58gbw6zHFN0/n1u1yl5GO908YCKd
2RHcR7zKZD50PMCCOJSdjM6KiZyKbdpxcg8bVsrHf8a6tNDFgP9oZAKWransPFdNfrsb3dY+2NYn
BG5OCcF1tnD/ZK/hmvj7KrDcTJz6gXelCGjUjCeiFQT2KkxKIYViEKY3yGtCjnx0u06sb0+ivebL
sFMHB2C1jz0w1t2n+uy2VCvd+eKO7hkJG/BpMQKgZo+4kcmrei2XydpxNBruV5WJUC+D/COyIiMB
oyNkaTXieeX6AM6DPbew8HFdiM8R9OilhjmnotFq7cPweZHZjYDkbPiLHa7X+DmkexUkoX8jK+lf
ImgG/u/Bmey9aoQ+glKonVXzxThMw2dJi8dgQCJZH8/BrvX+2FLyaPG1ITJg+TRW3EHDuSLh7Edr
P04MLbK1HWQjDz80FrYYafCmi7GB0kTre8AwApG+wxWKv/X+DTDTVFLL/gP5SFest7TGdIw6kSZQ
0ADKinkpJ9pxaThyJeJkKnDOkeKNF8YB3SUkzXu8wRoLm5UcPFFKJ0DNMvmdxa7RX4yeYuZ9BrPt
khABvQIUm9RA3090J+/4LcncGGbcgMVnFxAjJfC2H6Mq49nPlnWOF8n6/Eq26So0yiw2CeZ1/MrF
4oeL9lpIuxlPaCnOHTn3+7h3pQyUeJrlTCdpdgZDp5q7aXHYkIbQJBEjSEqBj7SkES92+q8hRWWA
TgPV8ad1fqQUHWykTdZ/cau6xnDEND8ZU0+TD9H4OOz7VoLP3sO9JG/2WG2GvarsEA1xDyG4gnYU
Hq1ixzLbsw6QsCGlKet11N1P2ZuMj1KdpmA3hTJwSHAytrwCAfzpqN53Hvw0otp2W24JezxhhB65
gIxnrEhK74YsCduu9nIDE3/VG2LmXK2DlF1DJSSnm1Q0CkWtVwvQmIb9ay3tnNakRVvHM40mWUFE
3WikW8i83Oe443p5rvYKwoUs4SdfCHvdskIJyIgeNLy3yWhIaCuqAPGoEUBMwCbroyMnEtyWl132
J3l/CSCEe5N75Xr9ctQFqEi3ypb5EvBM2i8JmdB3LJviks25d9PxXEcESfjliBR47V3erEl6ZaUU
jo1iwdWGKi/BfNqCRNcmhhLWA3LeDw2y9LHc+HoGYHWyqlrTWqQA8012XtalX99/e7sinGcN4ViU
ynlaacg7p6bPb9P5dZELGAqvx9cRz4hw6oAXJFaVN7aNl9MZN5olR8tu1eoXP+4bLxhyXDZMyq2F
bdUUnbu9PPlZ/iHia74vDmZ6GK/ow0rCRxr7a3awkjRF2bqjczywjPva+x7N37JTOiR52vYn3ANP
n817jVP0IaXcJYGzPeRGPtrIZ4AcASMr2NgO2fXlbE4Tbs8QaqY/KUqycI5pF+Gi2rxWmfZtQOLR
ZofY+m1x2oPerZJyHzzsWRCtwJbNAfR46pFc5qo1e7X5bGfvsOdkanR9hOu0ReNfybF3oWyEuA40
iE/xHnmKS5qg8l4hTrLn15MRqll7mWr7AYLRKbLr35AChHLc+OgOmf7TgWS+TW9MaPMzibu64kOb
9Z4Lj0EzT+e6VdGW+oiGoOrgCRhSrmCkkvKDAvv307LKI5zTMDIFhwajtqvLiOHn9Fj+GCHTrh1e
vI27U4kpJYTf8YX7hjGpkIo1dIvCf0/Xw3pz0Q2+bVTrpglQ1sceoujazIY6iWvZimpTS3AA3isA
i6ThxmN4tRYEB62KNU/gF0KIo4fnzI+FmQ8xAxXd0n2pD9QcjK4LPdVWWMkLp3rF/h53TRayTAws
oCFRT/W8F4fFGltbSObnFW93C6xzl+RKnB+xqPXNnfnqo43bFtThDktR3peN5qeBgA+u3MET2EFK
/cFqJcQXnQMF9FGai0KysrzGy1U1YM8eJGzRmPP2mNdjVB6zSlmFUegiwvG45kGJggoJJk82rzpG
5SCz5oa8B9iGYunQ+VzPyiqJcIhVeQx/CFED8sel5NnIcfpas7TLfEo9A0Gd/7cENYntRP6CEcsF
CbOUVJ4naPyJYJ05bHv/lIon6OZs7gWEg/CIxZ2W9vdPFgY3xufoh1okgeKoGpJ+wWHuNSdLFvoK
e9HAUxMRhQY0wAZpjjKAbQf8Nj+fxk3TNyGrEaA7jvuGocLKDk5EG94i1vwP/C9ebmGbuizwOhls
OtBnheiWk9FB3pwESQ0vVDW7Rk3Y5WFV+8uIBPRP1agPadrpj6x/cWYvrYhuGIB09l7oerKBC/M8
Ww3fFkUP13w8+V/9LndkWV2KbyjqBx557D8rfjQLrvLq3KtRHtm/idiCL5NR/xBUIifC/3rx0Y2Q
0Or+g8UnXPAR4tnUAnUuD0ArSdlNtmvrpqbAnETHueIiEwctER3qC/U/+sFGhcRLOgtgbuf+ffYS
XtOLPaxdquqj1eAyu2vKoqvZ3jHzb/D/CsJVfytRMoNU8bxQbPPkgKBAfSVwfodnOCYsgGud9sD3
uvhj57v96/KrjpLE/9Vjzf+GZU263zC7znqtvZdTsyIeMliUoZ3frr3RKARXieRpYuD1q6ZUi/z4
nDJ0z7zyjsrT34y6yny3VH+KRjz7jAF0Y/VkSvlA5EXg2TKn5F6yndOrQ944o78tFvJNKgZARQXn
mcnk+rOWm/Q6C1gLmRddjMyzBNfRrYgXJhWLK5jvARJEPYqckbLwU9w0bZW4TdwscOKv3Orchjj6
JzunWmMlc+Yp1yqjaGiQCH4uYImpect1Yk3t/2fNlJJal3WJmCrpMsEg35L5BMuU8dgJYPFTo8nh
s4mlPd3obXn0omYZLcBPMLP4WxuNOfHCyzZHjjlLPKd2RE1OqyKiFJahhfRyEhKeh/vVjYR6NPCK
9RexemA02ba865dCqPZmmSL8Ne37EvmIXxBcxwvEXdVdUDbWcjpqOPACgxc/Z+XfHWsnvS/imKgp
DaduyMe3ZH3mrvvEPFNxyiP516a6VMNcD13mP6a1eXzK9aGvVvDGv6fGKTkORXzsQxuGiHzuqm5X
acKaOgyN7qB0RgOoC7wwg53idqRUmNGuub8vtfRj0GTFhbN4ouhtijeHeJlhBpMo/AaLxzXfBBrm
XpFXhiIfx2oht+oiBm2vKkSflEN0/JGeMeNa3TyUHSdOdQ3bRqT92GdEDh2gd/Lh2IkfoBqvZAFW
+Q+bZCiidafE1nmhe5cI1hNNFxYTBIrTyQbzi9tU3CLfMiORY2Zp0guKC6b3yOyBEH/ApACBlRt8
DFnNYmJoYjATUWFQidAgpJ+zQBbD4Qm+8BqqQgXdbcI94rVP4+1aLoiopfGitFZS1KD5A5vHSChJ
MhizBjg/6zKpTRYF+DHKWLWPH0ouao9jlb9WngF6jK3ySN+FrXcniy1iLXcVumX48MmF43C9Ju+a
myvZ0r2/q2CUJGfJ1rGEH6f7nbJRgI+AyklcD4YALW3ntv/L0sdUb348S8lN1sKr8jkWbsveiHTH
TiaugYZYU60gaVauvZi0m1khsJbAkrjQ8aS35uEzC3nJeNUzEpMK8ojLs51khed3LA2enzNl1XVT
CTwQyq+dC+Bgvcn1FwRu4yhNQfnkxWNPUCZiaJbbJPAG9GqlLQVal8WjQJOP2tjzexZlEFG6GWAQ
0hbCgSHUxOpCIrwttfQICRXSszlmhtizIvYuUeyxnbe1oYvafB6BB3SOX3K5QFRJbchdMLIyPZpx
yDFVOWkmi9+R7L4J1F7+iYYTW6f9TrxzP86yN7EjmLqNuy1mMwbKIqIhryUiwO+yfdlN5jn0/hP9
oyT4qYkhegVX3GmrVriANpk+FAWZb4+Q/tb/vRHWz+V0D6yChcLMvUVRg2YxCQ11mDHDF1mBD06q
5XoWN3jk4bVm8ZpqCjEFu880BE8Vg2PX0uQ99iLmwlW9wbwHiUKiVrA9LRwokZdhZDl7LZyXZjQz
QD5UqcAiTJP2ipXxRuuOqV19ISe4e72D7YyXgHSPEWvPeo77wPiyt+saZHzKAL705SqX5BvHUwr9
nma/upUcMcoTYWP/alzyhON/FCNKXG25hRRIrxxWlZG11bNTSbtnfjAwt3WuEGVPTLXaPpGVhBQ6
BEVz6UxZK9nSsI099z0/rhP7yjcUIsIxWoyzpnRaUfiddYZwLgoHVNutbfOJOezRKzKmyxEh2+3E
9YzaXlSTUsIvk16Honfs4u8/DkS0ND/t7f6SQ0Nar6gx0au2yvJiEMofZlX6I/XSTUmYUSuEaPwW
J0eVxE2iQcoxCPnmmqRFuODi7C3lDmx+XMPGI7mnOCxC4hm8mMcGazAUYBmmxj1Y0hrRKyCKe6Lu
zRCixCkAMJLsW7k8S8EIBAbT0X/iizIqRpx9/AzvIF1TpqPhfZ53yL5CU+ahfNu3uRtpDZ5Ac/t0
YgVUyOIjJBDbAOu80zEbVKDqAlMfXKxHArN2vZQhdMz/5i9lonBYMUFCw/rhrbskFvALdlF3N+Wf
M2g5JYVsRQfz2SS/VBbdEDG5NnFwrWjocsAxLm87khus9iPTFiBqEUQvTIiFwfvPq+VO/iRcKHjw
8/s2m/nRlptZM/ET1ajOQIX/k++0XyohpD22ot5iAtdmiE3PuB58pGPTv5zQ0HgDynjeCVfRqabT
IffeZOOmlfR+gYkI7sByImEQi2IQCyaEgsOHpT574mqhe1ph8Mi8TUThPKVYjU9Ujv9fi7OEPpGf
bo5KiQFriYEm4gT1KApVL/RDAyOLXHfS9oXIymk1dCVyyBsTr+WytgZ7EgzjW3gCPiiLKREJU+e9
eNwbXXvkzNN29xeYnhlY8LeViyP52s0+Ne1CS1VRyKuezY1YJMG74ynAzNJgFMSyl710DvYuatyJ
ocVVAWwkv7PGBwHaSFJDkFrbh7LxtzXGDfk30/3ipeGmy+8XgVxwZ8lT5HCeZ8iyFewvvdWpRnXe
cAoOYbpMIombWx/K4lo3glaF7inzD8IHybLsJLesDvoMo8OYX67pZvdy+7W8FfQUvVGeIrjaPGYP
DqNBZcuDffu9y+LL6CgTz4PzRxY3B/P6xJwudwBu/+tbBfgLKaMKgwXicra04vxoXeNQjUDPyUec
Avh/srb8wUOZaae9rfk+kW56t/byaALY6kINxET8HP87Luq5+/ggc/dMkLfooFivAWmQO9rtmJhO
LRMGvKiyfAlanwSe9dNOU4NmVAVlYJKWybJ+UcSKuyZvl75ys2V5kQaWzYahWqylVQxgEAlo/c+m
hbsOD31YH9rnrAfC0bgla1am9THrnvFusF0odPClUgMm7YCITh0271CDGawfc4pT59i7BhJKdNIw
ieXj2epTMcBPTGb9vvEOGuDen1S8Yf6IOH1zgztDDP2HX32BlM0tx6ZtZc1N7UTEpPx/91WYA7wr
xiMlXQsp3vs3nJj4KT0tw+YhbqyGHNWdQtrOGZPHRUcCvYK01vZ3AC1m5SNDre93TpYUEGsUicQC
SSCnFOr2wnizrBlQBUSEX4dlgK6EFA0zKGXDPOBlqXBnYqE9pR81jTDlC16b2KijIpgpMXLtUEHl
ZDLdi4uxQPmoKux/sEE+hr4YA1HaQ8XBhDcpaQ8oSxibVdCKXRYIzuECsaKX8rqRC359h5pm2qdU
cj1Bk/KQ9PD7LbOhs51iKMj5LpB8HMA4subkD+HIzCVXpSWK8qkOu+nAbKbFFmM/bR9Rb5BrccHu
CeTwq3/i0Nj3ZNoBY8yY8h8TMtFAiuFfh+m0AKWwLp7/82wNiXcB32KFoKobQf0TEOWj2Ld5zPN5
37gM2L5WIdOWjNfsUEI+4pgvQQJ60E++Vb3pLkVnotn9q4qsZnEPP4HDP3FEhMGc6zO0h8tGxVdR
zp/fkhz21hnspcKKmNweHZ+7P5sbGBTYJLnzGurQIoeWtKe5dUQYGqwlzRnF1qO2rq+xrybBPVNl
4g/45/ihzkgBPXuFWx/LL6XQNQa6hqYZyMUGlpQcKmF9AiQVxbnCsWARJ9OLAhDpLq2heKXZLm5V
TozD8IUizyH9e6OOIXU2F+H2D1ME3jJ6GZgx+G5NC08V8Q5TriK45ewY8hR21hH6pbPDXP3iy2Io
7qVkG4bSSIG9YUoyCzegErfvsziAzRQOtjGfhf1t3KNjFxbO9OVAcJbd8daNjf0016zxa0JhLMz4
2Xf2vmfJ722ck2n1dXcjzzD+fK2vwiH/lsz7j6XZ+jCY9mUGEK6ldSkQRbz8NezTjsQocHGwzgJX
OzHjKGUPgbZ+vvYwCPAVh20ByWLUPg7k2WtrtJgdVKLgURayFy1BuEUSXHoufazx9xysa9kqdVat
1BKQzcERMutXe75GcwFjgpF5nV6WiZ2G0xS6GC9rMQPjXxLdkfIfE5iPkRshSLtGKVdVKt4Kxn33
Uk8eEI1liktj09XnJidF0gHQO67mWOME0OnwruRNRoKfJB9/l6JuNyXsg+K4NbAzKQkf3WcRYiEa
BhPQPcjyf1F/qgC/SBxeLhkbawxWqnNxa/cavLR/ncoZtBGjSLbFku89zmzQN9q5K3f8CSZ5utCU
yauQBRZdSNnXdJIZt6utitxD1NjbfdEYExtAKwFsHCIVdV0zicm93SvgIeKjFEKgmFaq+Z9h2Sgq
tl0oi7049p+i4y9iFcUmF9YQ0MCy1ClG4xJ0DXtgg+JvbFT9w5uI3FoavXfCKbgfNFh3YABkkkMD
KRgyCxH8RfFRD4a9OOBu95PNRnwDaqBpkKVD6axYHIxNH4uSjLiPwbY6PVl42cx4a2t//PbbbeTR
uTyU69551ZM3woMTzHmghF2qQ/R8JxVM3zU2RZK7nKtJmDsMdM+9R8bZt+n8Tw+2cy6Yxs5VA2jm
3Z+pAvJ8+KabfDLRtBa3DwAe6ZPxbW0lehuxxjodaJ5U8cfN+UoQFILSmL+XbwWqErcMCK+MKsy+
StKUvGK8u77UxCbnt9mDgN/JOdGrmpPv7ucbnB2WVqEA1dNUW7Bxgq/QJLLcrNt73ujTYUZiv8RX
PQjjvOm77QwxjpEVEQ6EDMyxSI8pJpddYw9GVGiEiSGkPdFpuoL5n9QL1vKMJwi85ywumR52Q407
y9maBK9rl6cQv8J//kEffz/mFFBx2TtyR17Nku/Jf8/nE7jgj1BsOe2G7tWlR8IUSznuSfMQrGvd
YOF3FeAgyJ7YRLDjXHqJSn13Cg0vhdrboHnRSNzcD02tMykzqmHh7D7YelbU4JY9eHCR/95Bk2Bq
4GgcU4kjYyOEINTIb9MxMR4YwJzaZiEqYYGEFtCrPWrG9Qwj+cUbrFoMw2DqNe5xvnyzbQClcsVt
PcpVVoyb40UV5ZvT2ZAkwToIonAbf+5qd6adItXExW7MaZQ5bfl1LGE0k3BCGdkyU7U5tf6HKIJr
dvNlhOPRNGZ/ICSS3AG0q27m7UFEuV6MtMVi2a0GPtvdnMare1W0s6aOCaGSfumccUheJm/HVnMp
epR8c3549ZxfYn+rCO06Wb5lnzQtEI0CmPM4w8w6AlxnFams/tpmudqV2zqTwI2PNtzhdc2zKtwx
jx2fqLa96Rtyi7wKBGsSwPNxK3e4VYQ2JkM/Qym2CHrW/e+QeKwlgrlxxNbFXJgmb0zn08bBKv3c
eh9QKzIKOvF3kdL8W0rGwE6u7FH1tuG7xCp7TZ9/Rdihk8NZ5/6ASfj45mGtzS/loHnZ0X5At8ep
OnGBZrltmaDF1GJbuNgJhPxjS3O6ivGbrl4LMNcoXTfCi2FNhrJmew7stFisaqXjYm47eyNSs1JL
0q5ZR1kRMIbSR9f39Z0gRME9dYYiCXV8QZkNlwce+Lpc+zY90t78Lvj2BH43h7hOfVlq4DWjP0lu
eTdBAC3jdFcLZA5I/BIiIcVw3jimRnlENJIDa3j9nnprOIms/akclwyxOP5JzRRP4pWN06By1NsF
t32d2NUfQNAusbPDZdNIjUEeGihCGKC8vFEoYZB2FjPX5mF6jJyoI7QOtvIOpdFMGae+UMeyIAf7
yHbyesDzibM5SFIzXWx8d8Zu0aCPL9evqJlFyidWOJdqrnE4eMq1v0kioXsAKDEYUnAkseKIog2x
7/PVJ35yZeVWbB3hU7677OlxCzsVrgR8V+SglWCzDYnQGKAbXtjXRMjGLO2OoDdQcWrpUS+eqyFu
C5NAalPBYUu2GPoG91XzI4bNU6AAi2rtgBjEJ7Nap8YbudcB0GsSssDVMOjKsfAHlUKDyDKP2J8s
bF/VJrJlAttyipMsp02hcG5skaCahu0S4bfXTjSX0PPPuU+IVB2P3H+4cxWAhGiBebLd5lK9QInj
aS3qDOktdNQq/cwiFbyMWl0FnZgFG5DSPcDlaCae3ILEG/UD2HzzgRHIVv14JBYZcs6RYtTRdO7Y
kynv9SDMahKUvQKBjujrCdRl7CUyxYt4VUKmdzLO3jN1v935t4JxJtI9u8AlFLMh8Bh73N3LW8gB
lSBc+2WvDzr8nLlu+3AEFikWdo/5PGrjo025J0X8QU3QjZ4tsYwrGXcYGzDk+3XmM27IaYjdaZJj
76i/A5vV/AZ9ppEa4WLasETrmixEFY38xRRs0vlQMwZoOBx6GEYu7/JizvIgGu2JYlLN40uSiPcn
dj/s/eiwMABjjBTIs2BJrM3QiXdwFmWJZMYyy/9loYwT5clh1G2z0mhsLaWDCrXLcEWTqShxujNN
3BUrOz0XqXQOWmI8UbggkNFlq9F+3ZaD/tk6V7K2/00sLOjdjlGaUTRG9xQDVcKWV2FW80Yx6xln
TOFoo4GdB+XQC3XHpXTdsgKWAnGekUIAw57YW0+uwURFUxLThrtIqvC7StwJSNk7PLFvDF+YZec9
UOkv5v5Kv0uaMhV9YMTRb1LVPIfHd8xxIhFey083AB1XinYt4TmL0TtLV/k5SiEOOLl3JBSaBrbk
+mT7BdWNHFhTrhKlvdZBCPOoz4KTqwD/FddWRtW0ghTUWoBms9ucLrNOKdtSaDG4c18PYbme07zc
XpgCJGOqRC5PCqsJMJAQFMgh1CR0yiJZ/tisQ6LoyrUXJrtD/gwJlP+7KWZuuTtfhCslbYy8f2Lj
gdBopT1atpZyYR9/mCGSFhrc3x9UNxx8UIWrvg11KF7mXK8bHeueOT8pqtrrfyjq9MrekRacT3cH
tXaxXbe7nOfIOhuwmKX9nrHY+xDH/A+fpSSTWjOF5w3a+XOfCrdzNirmcO2uPvqfHREbobSN1Jbr
vkC7NdN2yZNX7zIm8Q38j3tfS5d1CLJRS/9HfY8qkc9xz56IhP3LJ//a8J3dJRTb2KCcVl1kXJgg
CY0MTL0NespMDsDpkLLvNGG9jnln21t8zjxxJCGl8+uCEs4uqM1nU59MUC9+iL5RN120F87poxjC
8FZBED1wJPpQtnuHLf+h9MY0LAizanHrPUR1/JoZe16amBSrAu+1sV96lR+y38K4TpgNc58JXw3I
E5xe0T0Gt/5MB+exUgdu2txNbRzCDQP5Bp7cFERmmCgUnJ86TmUTxCczyvukHSjlL1PIieD7+476
L5L3DEUXeAGNudnOvw9pD2m7P2yTsNuJgWYR1Xe8iZC2aFIKyEi6dYZkP0WDr4FOwn+qWuFdx8xu
q3iwHTer4w5mWAOhvwlrys0QQoQ+BKkL8QGuoqFiXTD/NDc3KxpiBg7WyFwzqub5jhWfmSgwapXh
ns4ewigGP3w3O9pvv8Q1ny6UxCD5hwTjkOY2jCqoO3l/2P6ItgLqAMcvpPJff1KD6qmmVeuwgMzU
IXbOqr0giDTzkV/tgASA0BrSqF61T0VIbqM+mms0RHBwP/3XqV1R6vynZx+APg2QV18f3jgVsSU0
xnxAsHC9q64KKJrr3pc3W+lNgMyATW+WOOJtXKbhIlM9Wr8ENce6BjB/bCGtLkJ3cvRseyv/9z5G
DAIkuCSWVZptfu/DbTa3lgc/WCqrEyk/9DeGaY6u7exJR3bVuKRq5DtxKhrYCNjj9E96bLjqFn7e
0Ek74vfSCb3Sfrhp2VUcAK3EBwvRB5tyPXePOcKlcZCpac13cMlLv9DVJe1CBwDHr/l4rx8I0mKl
3H4R5t82Lc90jkCJp/x0FlhgfieWleFV0+FBK2ZfxkY3bod7rH+/O3CaTdJG82v5LLimzPJAQDgt
jiNwaNJ7qQl6kmo6zSrNnEl7NCROxEBz2bfVBS6ZL44Q2NXl+6QHbSBZRF1skjPoH4nrYqtPUvqx
H/uLayHHy/KGBam0iGX0+61daY+lTazn5C4QxDmBwNgUXB/vztFWOb+CZlKu7fbzq7ccGD4+OJM8
zIlMRgvLuRlOGzHebz4Xl+4eAp9XgyyUK1VO6nejQZ+Y+naxjpZTS2kY9P7GAGnNQsTe35Lt8QWs
OK6oqWE6M93j8I5qP3n3Jtitq9nlgnA3u3co9wtGG1U6sApSjB7fawv71jzA22dSqFczcDjtnYJx
YmtQXLm73vNbEAYSm48QfzC4jdxqBy4hDFMmg3ecedcXjtHU8XERes0hFCVVZAOwZ9U9Iv0I0iFb
5MrGP1vl+sg6X4eXGbk+wQfUcKh50TLsdlmXh3/wPfEuBqvq/77J9Vto1FI1JGlc9bLHvDUD1Ta7
wrZBBTR+UbC0dUX2dGGFUQ/5LH12EAYauq0hTYLMdRIXLrID/9JD0nk86ZelivBylpVJMhqLqrVY
X6xt0EG5XLeHXicucay069vUnGT6jAXn14xbhA08X02+qSlzbhxqFgvu81nq0cQWD1IqMbfJnvI4
2FndPXeLHD3D6S4kBj6fbUYps7PfVywpm3Xme6JsBFgv2qF7AkW7LM8zVqLo/aHIcozlyG3Z4ckO
8enMmI+XYgpgpwQR0AyeboUqly8Y9U7mNU5PQJxZwYKtycmF0Z8b9CiqtcKAbYok4EN/XlF1kzIo
6Z3ieJiGwSHppFkOPYMLtDTwh9aAFZBHEH6DMcI7kQYjbow5OWG5M35utd0GfOFoKZwhOa0j21Td
Uyv03CCffXpAXCcPsG4LqVHdp4ThP/uAKJaPqK6pi8H12P2kCF5R0QHsOj63T6b2w24B8W2l2Osr
W0RHj8ypWowH+8YOZmwpUYYUQKbwChQouG1VsBTNVK2E51MHE+YvzGvvhUTtFcgW3aLLI77j5Jjt
5yj6rXDpW6BVBRqEMYtfZ+OTvUN6W2+XVOVWKDuB5uMn5DdnQ2qUiHz9tr7tMTSeNdFzHkrkvLl8
Y9lxKavQYWog9OelJZMEOxosmf6pJVZJj06k4tAvTR4Ly+kJiToCjiVDfa5dT6rFqbHcnBUH9Zcb
PlzgjMk0X7ER5fS/uBYLmIMf6QgCpRxSrF6NpY9GzJQYCQSm2cscUq4O5EZPq6ZELqOEGPum2WLM
wrs7JlQ90ULg2Cwc+6gqDK+x43QC4pkpMfHQmwp2jHJQH8nEGriLHYbF1gvK6EuXXPlAQAdi+cae
OISVFLqOTNdaoPI2NAFgNX5zSUOAFGiSZLReJrO/Dq9m7yMROEf51dziXrgL5Y6V961t2+XuI24P
zyrNTV4PYOS9WNax/xSaHtAGMOkN45tfKUCsE0WU+e8WsGCJucrVjg5CBFM35HMnk4gFT/sFeZiw
4mM8E9o9BQmRzZjk8gaieaeuwpVY+POKiszGmFjTNHiZrmD6zUX4qA+sI3a171dm5lbcMFN8qZ96
DXu8i6OhwuURhEgS9NcUoBFcUyt642aXXtoOBrXpvTs+IECPaEcknKJrkhL/B/QI6/gDkEkf6Dk3
Qh+9WJJVS+/sff/7G8raDkFni9hMinvHFfn29dGqZ2J9BwCCakOxjUNmveAalhLNrrJv8MD0peuO
1q4JXOL3ubSHN6SEqpySyiTNZcHZISy7UPg84oHTNYxtrnDUyXIR++gulozohfUW+aFxeTXpTNmx
hNTrDep1dQOAsmSBn6LXYkGHUZsuLHI3qB+QZ6YcWhsg/ByAgRFL4P3AJtnEtKhEV1GKSDHH4F+S
o25TnNPCsZKWG8vu5OshaMxe2HCF8fR2vvxju0O3GHZaL6CpQ43y15cHd9IqH0W/TKwHhSpuR8H4
mSP5vbDD5y59eo9f4M+VZSu2nTqSesfbqv1cuwff01laAA36KjeYmP4oq5czckq7+V0YtEkFnzvT
733E3EsgU7h/1/1x558ZaaCydnoUDZ9k81guQuj7rEYsIunKMG7jfq7DkW9rgrTrPdNb3ZPlGyRV
FCJuwEdsJy/lticVvKtpAV7TIPQDSmQCywErNuDzs3y0AUSEjTSL0ICJW3uo+gbXE0ZNfWFTFKZ/
55n4Up92kU5cOQvF/2pOPq3k6H3JhDH8f/TYbqV39pcdtDojkqd9bVTUM9i46y2A1HIsCRtcUSt8
m63l3iKcgm9sAgELKiOrveMGpGp6Mc/FTMPxIZkgejRqwcqUXwBw6deyjmz1TstVk0gE+uRqyLpG
FGn/YMhp8CzbvrnRE9PZ2rRhg4pmSxRWYfJMsZ2dEsOP/pYzoPGyMxRwszOeBIyfPcF2e+6r+i7f
PYOj+1IOW23sSSm7n/JJY6Qu780tsEKZ+yZhSeduJJXyW3hLnsCdXWIH22re3NNE/dw6TRRwQxQ9
wbk5nAPxZC6LGpotWx3I8rBN2Mg8Kc0j7JX5tj+K74k4OVdD73vUT85JmOCCVoCNHRRtMSCyBpf4
+Gl+h6rORFZeAplMNU0SiKixUysopziUsdW5ATapGxELe1D0V9H/MB8IRUxBvfQyFVlbDnUrb+T6
Gqz9wPURg1p4SeWojShwhUgFtbgw+KmNmittSzFwp/sTjYew7R8281K2eMHEP5SX+EK37SGLsgDp
dQkGt8somTJ4vHgF3IqKMdl7Blwff0TQzMFqd8bzesEldobpPR7n7k9WNk0g2v0Msw4Ig1tmgpV/
hqyWbAd9PBW8L+O/vcgYKxyy7VqgQrwGPia077B/LAs9z7zSdgdGXFv2ZRhA8BzcCN/WHFnXPlzm
goo6wQDEC3vO7gY14hvdWhQVNsGp40Fl5XlDLk5CEa0uKiQTsfnsPu6gCsT3uIwgzvRJQxMOmQ1Z
vh3D8dgEmKfjpEDghXubaByYH2PuwxCqbxK0uSjRklAYMR5ugbOEowtL4Kn+m7GQCdSl5sOurp+j
6Tp7gsiP96aISSam/f8mdCUgsQjbMWDNIfoV+s6yN102IknjhFBkE1f7cUjKZT9F/ogk7dGrOHqm
gQhKYT5YsrSHp/3I+xwKsaZDoYhnGhOCgOO2BWWfB6zc0EhGYfswXgwYXZ3POzsj2ssNA88ocHbQ
XhvVoaI/HQsLNPlkeC4iHoK3mOwHQCFtbbiaYBEk8Xcy4jMcU94BWwVuTh4Z+nFrQI29Z22RKi3U
17rHvMFY8HZ2AkqJvdlzKXjs5nk0CSQmPOwBNEMTkSIJMmY7jvto0Aa12bV2B+aCOztlmzKoLOwV
oz/RPCeRnSzeeSSt27RoTH34SatguEehd41L/MYTBxWGGa5V2qnlVmT7pdPiv95D7WZCm+8kz1eP
T4c3ymFy5uWbgzFDMJrfKWTSOQ3PmgY10SX2lts4uoBp/D6SQemGJBIuW58xXEBMzikQGWDEcclM
NpFQATDn9Ot+9zRyN8iOBg+zrntPr25/It8Be9CWOUDzIY0CBtzF2Knm2ghqlxMYrbWY5/igHwka
ueJlkD87JSeq7dvPJb/T9TY2/5641XurF16arFyXEKwqqwCDsjyfBdtZm2wnF3IF6CWQIycG9Sz+
NxaUBq+IENcOy5+FOzRjo5dtOfdY21HY7jMGHdd+lxQLqIjWRXp65CDcu6hoRTlEtWuiETwY7BkK
MCWCBR/oYuj4nBUuhKTRpIblglZmELzxvcHJ8bbtaLRUvHy159zCnmuMmQm86qK/a72c8hNiEpcB
HNHQrmsSu36NplZWGji95Sk2DVqBj7NuC+39FLDcgjRrzIQIVP4UnAxxdBFmHBA+A7XfjfXzOwwW
BmkNWNlIODK8FgIEkc2/Zjzq/04zKRiI7EW/lrAByIrnQEo5R2uWKQhm/0HNSMZcPCWNZ54DyA4s
xbB7mhrJh+JD27111CC71EtxrUrTp1m5683sDbSKdh8JS01Q67a7esYVDV5IPLVAHFpeDvT31Chm
OAv0MI750cnlkdhlvp/BqxAnwrqBLTnKchjdYfnx4ln2LBTruQK14R+FUYUh2k/+MQZuNgrx+Ji4
GSNVofKy37zd1FuYQDChES8VLS5M38UDYgj2o/tSz+7HgmLLItQ4KzsreVVmT4HweJMOPSAC70WM
rsAmiNITPDcfi7BNDGDoDe+b6ok8oz50PVG6rOArXSjmxE5jRyEa21zto/TOVXAYGAUkm3/rTHQA
iYEHJwjGmBZZX0h9VCdpjNcvY+QGo/lmlF+JvilgYXH+jtgOLHRcMyUgm7zP/gNsnL4ZsjHEu5Aj
JDHiqghPil0ftUKn6Mm5KFZ7QikAgbySLpieblciILKxS3ZFRC0EKLOAw4giSDOQAqoZjuyMWprf
ru+FisYQ5ys9B4CuUNUNGQxda6WMw9mDIHJP9sGp1L+Pc+q/Eqja8pm1DVhRaaD4NCE6kf5WwSGu
B+WsD3a5GW3xHx6x56N/bY5eERx+QO4j83CwsqQgY4s+XpyimsYIIiVIGLmTOAT5/5K/yL6CzWpx
3IAXt/KWxDdskLl8SfgnGkD6whvRtrZPD/6eZxHlRdtyAlPaSwMf2uGfuC75Ax3zX3h9zqiHwi/j
RROz0FtQYPCV1PRU0SbQmE1ri1XkvSS84FDbQ5hnydZa41NI8Z9Nem+dnugfa44qyPFaEieDQMEZ
oYqSHYHE+PPiYyLSJQI2Oplk+jaJEKKIffszZSlmf25oBPvVOpfZWjRnho+hu4U/Shq5pKdgxVUL
oDyhiJnioEb56monce2f5kkudtYKPqztEGTuj6U0Tgs1tT4I28LJxwx0t8c+T/DstMLjloj8QZku
qUZlvOWqTSfn5erkDsYb19GhwZiuy0RXkM6UVRkPuz10x4VRCZPLM1oKODD6pTHmMjMhadW4kUlC
ynpQD8HWOnRB9e20ZwaTsJyFfQ8hJzetfNXYUlhhI7/0HgGWpNxM2xwqQ4LAbD6p4wEiETlywUox
RE115+Jik7UwSNeD60SihLdvAW1EoPFc3CdZEJa+tr0Cc4KaN1C82SLDyI7slR7x44RNAI9ridbm
3rGZa93OpktOThbeKgTM43h+xYRQp5NZ0IU1FUeA+yr5zMG6sAkB+e73AvGsu87VCEYaIsAH7JCL
DtQjn5076BW/1mbal4aQ+wgelmfSeTohoLBE3KtVgmplHz8X6ZzpLFxaPylpCQaW8R4YCeofHoOZ
A2kG6nonyKJfWTWOlwBQV+qxxDPWXgHMBpycb0TrjxQt57+CJq1kWwORs+fo4dadlD2sj0S2oYk6
GBVzmNGGmgJbkYNwtyV5GaOgVgCdgUJOOaWIwAK0VFozt4NPtETgP64ji2qBM/77CbsrYUi+IM86
Jx0CpsO/+lxGeO2MJWrg1kBEJODyp3JJ7QvrE2N0tTB6s8krogjwJFUz1I4xf01M+ZP1WKX1LdeB
Cjak4tv718ExcqHzNRUbSaw8JiCJVcSLS158xkhuSlVFR/nzepIhxFw+z2CIgHHFkrkALDlmUWTU
Ec/qh5u/P9A/x7ZSF8pVhzfF09wM/eIcxJewzGhrbm8uKd8cKBkIFFGWSYqE5Bdsc6booLwA46VT
Q8rNxat3VRxLGXNUwEiNfOIewzn+pM/T1H24+2lCGJImXgpoPs1i94WVwfmVe2z28xPMcX0GmFO3
qp1zYuVW4l1arJO4cOiszzEeGTWK6VhsnZdVUiS0UjXRni/H/+96SY9bN35B+mAzOGvgJHYwwlNN
DhDB26puul5IjjbXzf6Ydn3PEiQFo4/s/8fTxjOEq6TRxI/KdDbUGttoLMxdKpQy47hbw9K6bJeO
t3M9Q9cfoKTRWrd1fscn/PNUdH510BToBHdIg6wqkS7N5XxcxHNnNnZZkGfnK/YgPQEp+MRea7z0
cSauHQB78G++DUKpog5HF1S9ZHOiynPTIIG2qsOXEt23Cxl+3+AbYIl4KzKAgjRViHdQmh9SMy47
VRCu/zl8PjhLfnWWzUm3KXPq6O/87nP99kP+NaVZXUlNt2B853ktFpnzvVWhpZm72Xs4cvJx6Z+z
DleKKj/HukoaFGiNnNGRDRbgpFzJXwkgF8MRXu+QIZZhvbxF8N8RV8qUzd+yXhJUmjMmI8lvkEd9
olIf6oITAPaDGJrxwOcCO+V354CW0w6yxUkvRSdJKRO3jdBtONRKXouxMM3NGzCaqD3Pr2+kS0B8
u/rd78g31Na5T6d5FPygcImEIkG++NWyKd32o7oWyLhzracZRBTHqldpQShpvMk3tIhTjrzxN1Wn
BP+Fsr3o7wRoyVXulI0EsvOjKcWJSBTPSRecHWXdJ9Qpm6RnLl5C7JQlfY1i8EjPFn4yfmdwikVx
iMTFnLmQ/Km/ng1k2qbsOiMpRUEqKtSQK+D74aSqZfzmlUC/WpybiJ+O0hlNtx0M8r/VU5ldhEyW
pRTPYnJ4XMttGIvBq3PP3mMxHIwi1gvDjx38jS86i51WbiuAbFg1a0IpEU3+J1+LA9GpcVVDGALU
/T31FqDqPYz0fIVcwpAyoibIlix2Ma6Thxuz154TB6G+xtrxe9zhDdKo01ZyxQkjvs4PH2bLVkyq
Mlxw9qYrTDd7kmVXHUIA2VZn7pKsSqJ0KwTQ3H5Dn34iywP9qR0ZZF0bfSUGpRX1/+uUemLg387q
D2rt6qUiwkHvUtn4CijrPqmueJyl5tKDfyoVsMRNE1ihbaI0tJX2T1J06oAuTmo8kiFqSs/R920E
gQX7pPs1AU7BDODELqecO8P/bSsVVSAuqTai106THAjptRl43ixBu+R2d19YEhZ8cpXDXVy0F8Hg
gbG+yfJ/qL3PTJWNjI/t2n9PczlHa+R/dN0FXOnC0eCqYdzLmGLHVIMRznFuei/pBA8AKs6TmGiT
9WsDJav1OWruCloUXIj1rfRQhoi+5uiwlTYcGPUggO9TIXzsDTnt7IvQyx9qYvEH4Y56VLPJQglY
c2Rpr9OXskvs+o3oJ3+MWHkh1S96okEOt+4i0QMcmjKjsIce2kYfIAACHwdlWJJlCtAmczNuud+5
XwdEHaTZg3Tq0nIeBf9E2Z4BTcr+/D57gXnsN4Tk2lHxb+a4WULTiIWB1+dYKZwX7JNZAYhEunKs
eYC7gVnHn6SAwzDQOQMbDonRTlE1zirgALMj+P3zaqKAbscj6B/LlmbG5klYkcL/9etpREYqAcF4
+hWQ/n+b534X0bWDrq9MT8dTk5oHjEKGVQTIEzlQ/2g/AQCWg5mrnBaKNQjXb46x3GAN/zOE9Slj
B9jHd5gC3uESuWD7Kw2HwC8Sa1+r8eOmc/zOZdSMwzaYuNtzhTErYPJjdDQuhw19MzmIAiQOxckT
vC24M3nCkqFUpZDtf74Rk6XF4bCKle/wez8q2swQ+T9r+sXbomDkDWBdoYbbp9NCGvHGuVK+iTIH
LiKAhCbCmCwCINWQ49NScYhgmZqllF1wanSmbYoSz1SdY+0IjdugGo1tXQygGksX/Ib1NLD7m4FR
vD5VeqfR7QtnLGQffTvAqGgtE6rxQyUybAfzyTVclOc4B5/gZLB6InTghpIPRuoKitq9hrL4xznl
/lBpgSXo1FGfjv54vBxCtSV++gy+zVlzje1GGWWVNa8qX3rbKLMr36RClV+a7lWNmVzO5B0SbXzl
+kmW2x5Rpwgw6WyYpEokqbc9LqTsNqum/QCyKSD5BgufdwHdRC+SmM9/apomSZzUZU3cLBDSUbdY
JnStQ3gp+7XQFvp8s639goYxQX2Cq7aJhTl2pxwhGsvwvMu4FXnVsScNhmYPHOdfhQvNUhxe1mb/
yhmH3l+eh5eVSkdCiKatT7qRo3HvbRKDESULMf9oPiWQivYMoR6pc66vY+3iHWGWAjKW6hBrOIX9
2bGC2Oczd3asdJ1SP+BxvSdO6C4krmAFNCtrJezJPmWjguyI8RD/VQ0X6PJxb3A38p2ChR18k9aM
/ApyyeHDySEvXMXwlD8f1q/2PRGp7fnMwTmAr36cPuBr2rKIF3iJP1FYliusyeJUhqZ5Gnob9XaJ
uPCHIKw15SL4sp0uH7jKrPS9UdJFDXpvoCUNmd3PgePAPP554i77/Re/fMGE7AM/N/e3ks3FrmyO
kgrA7C6EGvy/jgYTrrrjFChzSCR+lYWBVV8hrq2pvmjy+HdaN5lJWy15yZowPdu4n/EEDwf9mrv6
v1NDwoFg9S+7ryAlClZs1OPM8+oGfrZoP+5uUVvUT6pzitVoJlgYqrN7kRI2mBu0T/wswqSFWu8p
1ytxUTPDojxyBoExHxvum+xgQs5ZwzFvATWxYm2mpQ2QkFgcMGM4nQx7Ux2JT2TKp3yvKOiQSX5k
Zy/nb9bs6fYw79ivCHc+WDN9t3d6k3oWezS5wH4P421zFJONslfKiEX7BkuHcA8Mim9zrD/+YS+9
QSnL00hwOGfFlOuhkwSjm6O/tI4qdC7cVO693umT/8XspVZHujWhTPHmXJIltHyd6/MWnTJfSqXy
bFyK88O0k1vupGXyilveBjOChwZdm8NXL5yL1zumyRE61bk4fIXu0GJIzEaalgMN63ib3zihpsnZ
o1HoiY42BS8AkadX7VgTyPJnzjTR0rsKg4Qzl6/NjVsfq0IdV3APRhzdq+4k00wV9mqT6nHuDjun
8walrjOBwv/AczEB8aXOBiz1ZvJPD2ag/lo2R4JKEoPSz0RYbFkS54iYVw8u+pfsvbLDcX0R7Z0y
n+bR3sVQdsSfRqkYYSlBU1pzZM4oEYE4mi9NwwjvoRCbLVND4HbPAiDKMVFcaK03ddp0bFvw01eP
/8NBgl1OpnpKh3fhSy+2pevWKydUY73jnH68eerRmhDOB9WY+j76jVWxw9x/y37SfPXXERV0CBIn
Id02T7JI/P3ldkDM30vF52auMpBH2hUIrje8vLRNlGuIAOOWn8JMSnubJDDE2LWpbQ/hePBTh5Wk
bGbYE2MSm4JsOdGwppvIemPB92Ejxc/pupT9aj1BtMIYIsQZwE9/d42yt/9LJm9vLu2igl2yOoT1
jAfbCtW9Juss21FwjrrRmm+p7HwpQdVAiKPPLTUYbmYYwPl6U10bbgS5QBYYNZKCdex0g6GUfYBG
ifL0e421Bulhm49ONUwO7mk6uu/SFKPmF9B9q2fLux59GS0FW8E/StNCSQ1p9jQ8SKjfRg112Nva
T/60ZpDxs8/j1HQLvdFhtZw6d+GjQlRbixQPwmhtaSwvvOXuHsjhvXm37NqRQ5lt6MtYJ1Ax8rik
eB0TbozRazZzjYE7qxWKe1iLNRymS1g4UgT8PYLCsFRTqtZeWiXL2PJBeUazJeouFEpNGCK6gDUf
pT9Eunu9heQgmb6kxhHDmZFNx4z5R2vq4NXac/SXalURJrTOcfHB782qQn8qcn0P6fXJifqtktnI
mocSpNhE1rVfi+oRMPUkKvc8amxC6YclPAB0mGn7EfIoDA5wnAmJkdTbbaxJf+4633ZHRlemUGXd
LQ0l6xpgDGQpB6nDKFG0xLOmdz+14iohO9AeAV+wzfJIM+/48Wk5a+ieLqH0WJKxXwWPcjr2qSBs
Qe/kQwUH3B0k/lAF1lGGsHnoTJZ47U3Twno11aa7Lz77r5WsAkN106/FHPc+dPQaqRyZPyFsVHHq
mxRv9bihuz/nhwZXZy2t7qsmuf7LzgdWT3r81e30HmCFCSD7CHycZ080873xXW8txa1qZgf8YVBw
b47vW4yTACyCP6285PLRrneY4uPjIsCMrRLjbn6ykbAeY4UiGjQH4KWTGj2NtEWHcf2T02U/UVUs
WN9z6++Bmcl1EU45dt1leKztwAcv2bcbmBtVbsl1wQLizYoKdV1Q4VO7VVDMI2QH7ar+7Ye/cufE
T1MeL2KebsIn8pB1/XJRPIzCBSrY1eHr4LBwNADOdZRYHcCfwcEkhSqVLSalr/wGZCpWSsQzm2V7
pTjKhxGO+pwp9p4SsUsdbynrkkiMGpN/bP/60R9TLELYUHxUAi6iEADsEZYEyddapyHtPnFzRlnl
XVV/FsWvegdqECYMFfYOlVZ2eEeSJYkmp3t36Jpl2tZJFnqcfbNhvvlqRgBwKbnL+4hFMw5X+hK8
AjzZYeCcHOe34Roz6hTRP8Ea7N7cPzF4OLyptVmzkN7Euu1VeIEOVw8ID3+GnASFwNbZmOCa9xz5
/K89YhtRRfVoYAdRgKlsxMPo4rZq1tCL1qeUlVmpukSNN4yGsw6FDl0kdirtJdTaKCojnpQMVSQI
siUbJxtEEBARzVymwcb6RP0mnVcm2bJAkN9AaWU5gNiGDXyeobOoHEHvblOGTGhM5DFXmNh38xe0
+ay3BmhJr0s9UDLIC0lDZw0k4IgmSaUpqznP8aEhZk5COplX9TcmmPpmV7fwlHzOOIAjE0mXgbcw
GG5qQipDHX7UJ1zou7zgrNhiZVhgU1asV2AK+fXMJCmF6gx4UlSjC1aI9/dIGT2+kbYvL1JNzoVX
SmnODdI/JGuJwakiKjYB9v5Vzp9XFidLqp3lFN6X6ir69/+gLdMhgUOMQEbhtvgbu+3WhX2Ew/BR
95hL7xcEOJwHar/jQ6LlyP3TiOK15e+TQzf/XGFnvWCmGDdBobQoTJ/srl4eX+AYkBRarkXnTtgv
x1j+H6ddrUspEUG+NybRqmX8N+XgJMxxrYShi1GeTxSgvE+irX9TkM+No1XKx1FXQ4ZQ+Ky0GWd5
0ihHB26npFNoyIQFmm5pZpPRyR52ZWGjZN0jchQyPP5/J29hbKHlszXcfUK6deJBWY4xXK/4rbhQ
1jlGt0skw58Yx28mz84tyWduNaeL4EU8ID/N9Dpv9QhvsdVrwuuPEOQlN4nSpABoMT2/+Miwxiee
/nIZ4jjtKPGWxZj+p24xzomIcZnphzMNrE+5aygjTN+5hbNg3dOXmOLG6CON4hQWOPbW+f4t9Uys
K+hTf89fCy7F1twqgbFW4C6Chb2yhrfG6gWCKWIWC/Y04tQWojgVslGyqZ9q/EtQfdmWVbkbrkiD
iqAch/i4rqeVg/bmFPc0x92M3DiaktCMZeqwTZrcCLGeE1DguZv4qEkj4MpfPHnHvUZvmENRMNWe
BaLeoPn4RCYxvIAKLDOw51Wh/rshCbRPVvzILvOQwuj78IpC4ofW9DFyznr1bxbTY/t+izTHLvvS
1fpn1hStMZcheE7zKMVW93VbS9rQNuhro4jXjRQ6iyX7mJ+dT9lyy/WIXrn0CiREgj3FyucqWI+V
5ES/IzlTpkEbkM3MBTjbglw+/TLA42K1XCuWpFQCQeRwhgc4hfdgsInet9uqM5Qn/PWyeoxNdqro
VRDj5Q3PQC6b5RG9BYRLL1Oqzq+rD/zyx8GhlA115CVba8zYI9a8ysFNaaMbEbq0M+LYr1NPrRSr
b33b0xfykNOcfH8R+GurRMIjk+qjHh8vq5/H0ISDMtmzRLCUh7n8HdFCd2JKl9E4C/x2LWBUtU+a
dw99uvJzgMAKDUhcIoMa7eVeWdNLpzQSTOh3oEOKgKmLar1g1ndFrCeYJb6AP+018MhxpZEGaFYU
6EkgGOdKV4W25JrPfzpglw6hAgRb3joINnrOSHv15fw/HzUjlRJsfzO8ybN4W86pbDL8x9nnU2R8
9lrSZWZs045wM1QQmIVCXPBW08tncPQZFTosGYWiV77hWLWlOZeIN/SDa6CdDHabE+yjpqRDZ+0+
el6H8qrDHdShnIyeq80plwVpr76IZSoDBUyofd3VD3hR675hUx1pfhOqJipVGBQnuqcjlnjk8x6q
wrlceQ86olG8SBCZ++fXqqxcBko5iTWn5Pfr/BJkxli6b1XecAmCgVdCMDqt/e0YerF0RPznVwB7
4/fuewS4wt+SRZzE49UM2r9brRDgTLzzeyZluSWDrFKUUz+HACgXiHUE32lOvernbBkRvw4G7VCq
25i3kWzOGXiPHQFDylzCy0/xev9RlQJdYogxxHioOfNDqV5UhMZj6VEF3c2/NYSHXBNl9l/k7MHD
u+nhJVmLpvvb3hYeIBelAQcitJKgwzQXsRB8sMtVfaA14UvyfDNvIydYVdWKDjCvwCNr6LZ+SBv2
R6bOL67HafDUcsFVmlIJGwgiIz2YWIyKv8csH9xqvJoY7NAGh6Vmpuu6WNlH3p1beaG4YJhIXCZp
NQGzsy9BJkb2sBRVFkodu8xULMMrJtB9Dj9IaEFBNxTwYTTskRlJ5ocubP1QbuyIcD6UziCZWdHq
IevWnxTG7+vg+Lt+1r853C27a//2D6j6SylKF8cSA67+6bPYGfiMBa0LLF0WdrGXt8KAsuq+Whqj
ACDr1djAfPWUNE4+rcQFccDJU5oP1LWYUb8mcbGqOrAcko6RtpF8x5TD/IFFxKK2KfNbW1eiuBFu
J1utuLVsqwBtEooeoO86QRNMLdAmGPbKBszxEiN0fMYiwPU3sn6nMtiiYnDjGMK7QtNyZL9EIxnm
VA1F4/xn2duR+VrIxJbvW6hRFYeE5mD4HRkIXVSJRA8HBC7JBcuapnqBvc4Txm3wMOsJC3S2GvNE
OhnVPHiaVYCpBCS6WCG51pT1EIPyiq/+yhxuPLBBqwptBsz9vNHDTefmqK2p+t78kA7oWq8BV9fM
sYEfmUfMwrYdjrMmQJH9OKz9WqaL9qg2YWu2Fpp3epaF+K2x/FlocagK/guEEzpDJqOQp7J0s8dI
rOdgY0J4HEGgkyNak+O2BgHx6CfnWd7TQNnLdQdFIJfsiM4IO8GDfVUPpp3z2lPl0RsKTAbIOb9J
kGQYNwat76dVwdBlzbsbxQtXjDipmIjhXQsPfnrkYFoxgIN5q9jtPOBZy9ncJxUtJuwIyau2ebRD
rsiEqPtIsosK0cplpMSoZHL4IWyLiclSs3xtRR3oSIe2rRgZviSCFhHKNpFyjaXq5Pv3j1qmVSbj
vB5Crt+J4J7bF9T9PyxfezJIqpBrHGns0BPyjq0hho1B0L26iTBsoaqMfoQ/KwlutXogmt9fyZlG
AAAGMFPhCAdZWNMBrfMQrQQyEv/K0SHHp4NYIAWAhOgytkd3U9ohTRaM6ZgBn2kx8zB0ioVRKQwK
NfK3X+0Wt1o7d+e4FPckrUM5VSbuJSb16BXaVfBRl3WyyjRys8oOCpvt55izxv7WjuA2trBklCPf
7YoW4u4EH9TuPFrpJvPInQep61of7UjZ95YvhUYrcWjuORF26C9O4tydur1riXI9zfD63o0GTSXT
DlBUFYLzCaamT0JNX4s++hSFDdhDj79sBgHxsO0hVyfj12FePEyRMa+2Grf03xm8DVT6PKPbi3/C
Wf0KJM1gCiazVPJVA18e8reNWoW3ZQFIdh+kb0dO2iVqijJ6Ii4+aN4b76nVnLp9VXM7UvVV6eyx
ALpkfvjbxXnU9TlvQ6DANoNywmXRQ1U2qjFDeZ8HhVqSqoSQUnPXtaxdbgHGQtohzPbTDFV/F6AG
4nKUi7LksTuHmXSKx9FgCv69CwRemQfZR0A0xvGJQtvuDwkXtgWyL5ex31Vv2uE219UJKdYfgtIx
vZKbPnuYp2JHs3yCMK1h0XwyeRu51/buqw6CTPfHGtKjjP+yWcPJvIZonRfmpV3q3tC5B/CzuB2K
FLtZDsX6TPCFlpwL6grcz07E9onResxq0noCk+PpucS3FWAP0N6jdUqSg43CV7xoKICKu+v0HMeW
62Xpfn3MvCwdkuO9HBez/cwzEuq4bcVZrB2GJTrLS515maYd94q23VTl94hGiC++cnWzml1RpfGV
c/i9cFsRFx3x9JIuyTbCwcl9nWZGjGxD7maTIVyshM7+ZcQRhYBlKcrUxgOfOFs2Zo6x69OOsHMt
8+yhSpDLIbVm+qDVXb7eiIE9iK6kA7k9x1eUg00mjxhiTKfupbiQdn+Z5X14XMX9kRPOrmUW40zD
Hon0+VmOlCBtMT92b9ZnMaEERI5JWiZKIgJbRAXRmNxq1qX4awQAOh2ntYrdo7jYdR6GqYVfqFxi
YqO431MndkSLn5iebogeqhhTnt3KEJVdXe/3HQ/9fQh/i/wIkCHbLF+Omu/4faoF1vvVnDlUyDlr
IF3/e/6hNlChwqsfk5c7/bE7gX8q0c0w0gGTuoDsDstCZbXrpqvdPOnyrITO13HEZn19tD2/myNO
CihxvPYtR9xDZ0rUM1qN7lbI02M2bPwK5qYHSfY3x4GOsMnrn27W6h4xrxxyDLfyIVZmeTGQxZol
zaaSMIAte/pmjfeJMDEyUDrVw+do0iSHSyXD0W3LpPp54ATeA8PEaE10/zpawPMNXSldNBcU0bpb
PQni4UkQsCca163gI99xK/zxKCzPo3+Yf3s0Fuvk5mmGNjC0OLAU0uHjyS8pmBzZiJcJNdkd263c
s7yJvtTDCjpgkv0Y+x3Ns6sHG3TZbzRzyQsMfRzgZymLTFRyGlZYyJigtKXhXm14+5i8xCScQ0R9
ErRvlKeVaYbgy6ynNVlrHoOxBFwebvL+Yq81D1KIHCCBPs3+jLhPPX5quIq7JVrLN+lF7YKhFAh1
S/+HTBPNNLLai6njUJCZwULs3cGHD2QqlQlUFcmz8gb8tCc1SNNDz7Um8NyV9Ys9pWp2JBbGPjOl
WEsOFgsB4rev7CVHX2mq8ZkSf1hmoHuEtBautcKowKf9UuLFeZy9la4HpAzG92t7ks6sjYAR/TYf
QA9kzctK/mSvs6i1l+sChIACMMNyDPIQEG2gvrEYTMit7rxMvJ0d0y6WgSMqjp87mNDubOD0xPnn
AzvWj/YRR1cX6iOWuc+NkoWQRBliTE1VMI6KoLupQ/5WMxO+Cjh7sj8VhvZ9BgGfqdGx0hRDXlci
iZBJTpI0p9iGbtEpNYvrRcRWlQZQIcwQ+yOItXBYUck9acaMPHeLxMDFWoUj3Z7GIRQKuuvN/iHm
KlUIEYTSD6DAWcnHKwR2+0wPzBRZKsu2iATGDSvT2bwGOenmYaKt6DFQ+gl3so4BC6EO3EcoIGlo
jpmVzy3/xdpDwLnS0+w82h38keFEEjEOLH2f4ymu/RAnRILcOjJeVIKA40GXZJi7E6rFRySQpJGe
NRuRkNpoE6dPNRMgd7hVtCuhjcmDOv98IglqaIPSunkvYkKT7s793F0CWN+fTbYKME5kOurNWoNq
/ABpif6vvtsPRfaxjsRe3UREG23S9LJZG80WcO63QzOXF8Mo7e+9gTycciqvnPuvm31A8pYW6WXE
2VDCKJ1aRN/XHWYwaKHgMZcZLn90TbP0VQTI6aLX1V9YMToDQJNz1vEiO12u5m+Z2l4qjVuvuo12
+xDWtV3B8dlohn8QnbDILcCotAq+VeEQbsjE8DhywXS2na1NwbCvQ/XAUiA9Vtdj7B6xsUHR0MBt
6mBe5NWnggUxxXhflFmYX9gOo2AgjLtf8mXewFFWeSz61EIF9UTr8WJcDlNtbD4vZuw0LG4YHbmh
JF/2pmScJeAiO6cwGQ5yXW96gmeBb5FVOZEwPiKIoygfckggZimVjoDcafC6fAZaQ+YLVRYiHP7q
COSSQPRGkEBM8tGH7Ty2JrSYVa1nKZpyMdkHw68f3CxCVwzRb3ybrCQOrn8j4ZPyi1yMHetVL2Et
U7Ev7NR5vCJmlB4Lp/zGuTKQcxvFbeJOkt6vUF/Jae7T1L5TGMaVTlyYe4MCZkLtP8DRT/K2mouP
N4fIxIVrHKfvrn1qzYoKjUgu2k58LnM6BAn+cJY50LyBJbyOHf3k5VIhVrrCdmiGzSIkeInY2b1Y
/8Bx1P1+W/bRBKW+PDSxiv3lVj+N/3Q3cMYh/Lg5LTfMvohJM+Ko3CbKTLcMYwDhY34w+n4w4s0/
p7gjhh5dAt3O3TDTgVy+WBMuMwffr1RyEAI/FWV0dVeoABeGQGqbTkF0YjV9jFOEt+JIGeuAVZCl
IwynYgnM6PsRbuf6a9RXitMHl8dLoZt1Y0RLzDE/Yf6Gxxpn12T4YAtbmfItr3oON0Hqpsv40md/
ILjW2HaS2RZZ6DJA2/XsAMy6qbN5j2K55d34XKUGb0aFK9bFdKmTqzGJiSHfI8mGfAy+ldVvVLYU
S+Vhi0XmcoEuwUdjpfL6osmwe91wTNZoi9Q9zghuoitl8aTPd4msLBl7bvNvkmuHtGOdU/69IbdD
6/Y3d6slziCaN+ADwEEeeL33+BMiic55gpmjN80t3lTplcgMSwaA9sj5gN+Ni/WLiSOpTKTISoxK
R3/cMqSCNORX/ffdyOXfFh+EbxF00rQUpzLuXJCZQ4qx9qSB/mb8A+KEuVEQMXetT+nwJxwraVq4
Q9TWekLuiY2R7nAXspD6iMENfM5j7eTZv/K5UEPcdJ1yJyevSPmJ5GLaEF0V/30t6FravDfMXXPs
SXdMvb7icAf0CuD10ueTzMpzkWAAF5n9VyMrPh7L96XBg9tEZe/0j2PMewyK553RLra8sGVBJqdn
iUC5sKEVowaXNcYISMMPB2dulfJJDoWXFTZOxcCMpycNwGA1s1JVxcvASDJO87g1jyIdFvp3VnU8
wRiN40HeGv4ZkFZ9yPuNV489mJfP1rVaHh0czcRvEV6x1CJpWSQ5mz0dhFP7TMFqe9yPkGd/qLI+
OFPuQMod3z+Bc/RtG81cJEQhrdRaiJTXmW/eK3qMxTRFOk1Jkh6pNPMZGXjiFtVfVNFlLTOYGs6k
1wYam0y5fKlEZhgak2RGdEsMARrbRvhcaFAVlVhVEllFx+Nj5b29aMXawYo/ZiuJdtvOe75Q2wNY
bnpI+2g//WibdzWrTtQduWZXzTCXpt2NdolDazKRFb/wcID8xjvK1tt+J8ZeaQsonJ19s01AE4ok
42VZe+bnH0Fqkt0QbyU2SkWAcc9Zk9f2Rv+9ki1h7b5l5m8sRAFD+NegLsRQ41vPPxKp5cBxSGE+
leOSO7csC8tksV41HVt5r6LO02Q9D6xU7WZfuSl/WZRvpCeMdAIw4jqoyTP+scW7lVSz3YvMTZOv
RstnXZuj69BcB4CMhPczDbebwyqmJZiVFlCMRuLyOq7iVrVJ+z8LbR/dWjB1Sm53FQI6f3kT9VJP
+PKbFGyR/LEh1lUVOJUTq6PWNMcFc3EOcEjoH9scY/P4T58y6arPEAcyFSB/q31OHQq9Kf8Sb3md
dM39xq8YvfeJRyXBlHDyY1u3lNwAKzi6cIwc5uyP0ELyDxxAj1d+CiZsFvXNm2aJwORyO2Q3K9o2
cnLNDtz5x3tcx0XDdaWmu0wgqTU7NxVpUvpm8IvE126QsHjGvwZ8awkDjHSxjJOhyfc305ODG1XO
H/D1xxZLa1ycRxImijHq8h9hbTq18JJflnRc7UDYvgASG05gENKa+RUi0+S+bY4jznEIaz7PQHlA
JQYJiYBbtv2oiSs7O4cffgeH2wh9CrQBAAEW+C8WxU1CVjRzQ7Fgg/yBkP9s4UydrDWktJ3DyrxN
2WyEkRfIeXWAiuZKf0Q+7v55kHIcv83FCEPot66V5ZQHiku5VIYHX6cxyh8GAhqHiGQte7+zUrR+
+VX59zNx3cEQh4+Fxplvt/qdRYnG0bl51HyKmPhRzTXxwApNPAwb9Hpioh25TX8llhEib/Pjt8P2
arrrcE/vULZ/6hmbFOMg3Ujd4keEU799OaR+oXbSEqm4f76UHoDAATjLgqT5o9+2AVkIUWX+qaEk
k46MVppqy0IOBle2zWuJ/2TBhAyxWu3/XFWKQDu3LodZTYfQgtoaMrRuAoEtO2s2KUavAHKSGpfL
WslCTPHqcw3knWOHCt6liMJCPnW60EZVCF5XTWJ+3ftvbi/8iUwoDLAMoJFGBIbw6iCtVBiiXL7c
uXkAm2VPNvNz2jqK+2agfr/J364gQUbW43Phfm4YWm++xXq7xhwcqmbr4m3uTN7gaeUBZ17OFVoJ
nReBPcfJ/YIH24kzgCak0CBXVlJWBtt8UZHsBU6gGRIoz3/MBWlAMO4B+3EUv4JcIP8glPZ+0Sp/
0Gzjb/ALdrmG/erze+GPKbH4rC/OJg5gn8K8k2jzgi1OBu2k2QJgrXc7su90Yk1hHbYKkBzyaFbx
uW0qZMm03XEtxuXPckqUUjHy7F2ql4rxw4KoXVMQbfcaeeEiKGjv9eax807yZUgFCcVVfJJ+l6Ji
7euras18itk0nDU9HKlb0BeQF226mp20eS9OIOi4aQulgQnW2XrclDHIhzN/wuEA+8rpb18BZ0tP
y+V51vxuCXqUu04IRXoH+s65Q5iadlys19+cBWS8OmKrmTJkHTmDpOfGhh9oWnbTBESUKDTE8OIX
brvI8+RUlo3jmG6C0nJKrpRQ2OvFhPAI7uqjYHazlDan5vdVl3u4bFJ8rkVIdUD1Off6xZGL1uz+
nffxWUn03t1J6ROTTMGoGZYXp5uMOklv2sdVMWeazQjgUKhRewgibI3scBdf2EDu+SWZMa9kEudJ
ZGWNdP0AYSyrsv89E2B6cKq7GSXPpeXpV6mkMlXrOKgEw6tzFEm7IuhlVe/xfPO1L2flPVdOWn8R
p1T2MAANSqwiAnNO4TXFmVEyJUzHgJFeBxbG4is2hnCUrHkmdxcp8cHPa8drwZTjg0v9DCe0LZKH
Ro/KW7BRHyc/x52+E3P1qKhx5nuTNtseAJVyEBGvwLxcg7306CzWBQHe3FIYN545po+/FFZu3ZBP
HX6mcwbGMMMpxU+Z7oQFANyHIkFzACWOrHjajc2uKhSycCk3Ccx1vMylYOHtvX0mrZL+C5GcvQtH
i7VxWfrBp/IdPsSZCEdxWZx66yYtuZ48hJdPRdhYGIsNyiGzfNsOXuSSMHdN4LVBHtbNI3wAbuFN
gpp1xTqtQ9lq9fFMtpJu0CC0pT/R71d/l788BgyZExMOv/qTBYryWRIw3bjfsy2iXAR0I+zpMYld
+qmsr/b8cTrOD+Mq3zULoAYw025yx4KCy4maHOltBBpuEms9/dZzTnzDjjaYQaXaxf9NjQ0kk/Yl
fIPVmrNdTRZuDEA2oZ5MCaPeiMdxPuJGr6PmVN89/UGZNd26x97mvsdD3KetNHfRSvNxD14PU2Wb
o7xWTSGr41NXFbY2hrxeIzfAJWMrW/OHDQU4oRMoQmufOyJKhA6VlddOmy7HDX5t5k0vLYBB04f0
15oAgnJg0pvXLOpw0wMXt5b0ntpWeS4WPA0wFEhLI4mt83HuGBgkGoTKL1pDRl/IsNU6hqp8B632
yG1D5SIA/A1MFfZsV2nvoly+sGZtZCe8ISKMJ0VftJ5mcTgP2wLfEJ420SQuSmJVl6Bj9C7vMr+G
+wIk57jD8OZp8ljxsIsFv6It0uuAWMKkAd+ruLsDaUXNUjEaJksonpNgU6IfPj2jwmNwZpOnxd9T
NCgaiz15H9uHip4H9w2Wxi1oLNYfG1ZGj5zzSapXw8Ck7OsuXMoRmZcNjlclTq5ZF13yMH+Iati5
dbEo6Bim07v8wFEWbOW4OZq5eqXj7NlcFjcNGFrrJq4l6+5niAqLbBb1g3tWBl5GbBKdRxnU0bzi
V7OAwvoc454OydmN6SchuvTNTMn9t61In0rshBGd5xjykQs+EFEaSL+B+mH98NreIY9E8E5VxI8g
WvlgeR43POqBv6o5nxtrWs/H12bfKnDJ7L8BhPWHRLZ/RZgRpTdE1b+fPD1MnV+AHdw3BrSaieY6
0GzJh35T2J3Cb0KUDKM/ZySlrXYk8Oy3MxqikTfRKbHBKFC66q7B3M7eUHwG5wOVA7/S2iW41hLA
AmX4UJJqWUlJlfp8pRx+qxhBmuo1pjOf7/K5k93EESziJY8BGrGzMohfqofBUC8hag7SCrsBQbA2
mjRvaeslpLhGT3368btAv8e+o0XhcsILbtBN1bnHKIylEokVsGfX+I8WP672sqViXcVZfrh5dins
XAVnmUDpvmKAD2OyZ6OLrA4ULg+9iVlhMqY8mfot0ajYCDWjZmEJkqbv1v1jnKrqjhyjs8h8NyZC
pv29FdfKJ4h3avke1N5DlAqECw7WMqeVYGTPm4ELoyQceyNGE0QZSqjPSAWoeOrH4hhQv5x3uS3/
Sg15mtDo5QZug2jevqD+ErnmJII7yR36PlZEUvs7Uhf+MBH6Gcv1fmVw5lhIMRbidYboQ8QQnrll
b9imRL5wOLI/ex+y6/kA/BtcWBlnrFS680iHrsTDToFQbxSytWqVRQvpjHJzkxjjjRGDmcRYZXL7
8NQ2IdJgsDgS45V5fCltD7K8A9x8Jo7l48temS1YptfjTWVPBLxslaK2NiEr5d0zn0AlbxDTghcv
NKE27PxlsmLJyQWZ9Zb4ZPK0utQcQ84DQuTb1OaZ4U9BI0dtQ8FwR4oGV1jxhlCJaLBt/yvRYWMM
fLm+YcPJ6xGyxWUl9NqQ2PdICoABm8rZO7SyVnMDbJR1HvSO3mUvwZC1qulAJ0PZsoA5mG4VxZGP
pBdDcZuqkBOUgqe3EQlPa9KYpD7cnZU9ZoxU00HlqqqQdBAOt45zqePuzGYaSZaGRkbFkeRT1rFn
5891Z2XS0ToQ2lMHqfCb0tE/ssIWkxve5Z8SNCnW3E0TutZR0JSAN6dVtBnTQ2M7VY8Os0CyZNxk
EiVLYAu1XUOUK1WuIxfJUqj74rc1Y45482fqCMwwzl+cXhxQfpz5FyYV5ZrFl1jBLJhXKTAa4uN9
p/Fr/VXXSGRFc88zkqTE9f/DX9HH5w5WtbYLcH8sZekQS3JJ8/CDxH7A+MHJe5+fgis1n7uSH8sS
33eQ3E6cVLjDeM//PVV82Qokm2Ymgw92p9gUPSj8xvhTz6xO+QciR9C8tvxFhWq8Gbd3YpA9p+N3
ABILmKnD8Rl9a7eprPOGjDOtQbXDDulLRYFSgtWOnDqU9paOiZBxJxTfRmXLv/BLcK8HcOn2fEge
SEg81F0QOfhOh0x3m00Ro9Z1iH55VqjilIItxeP6Z6BY9WRNI4r6RBXGoTAJ1cqS7b4LEvr+rYMO
HCzEv5O7RkB1a9+RcqRw/TO1wnhu41bwwYJyYcuI2IX1tX7UmUYc020WQluF9vJ+/0S3pwVHY88S
REVQ7dixvKsPGk4ljwPkDDa/+XfTwVF7J0t6cWUA0Vm+y9RtZL7bhCWuZtXg+vp0wwZYevMR5JR2
91tP+O/lNIriRYfrwjDl49Kx6cwigBlPTQqyXmYZqJvQGYvnq/T2W+13JfXLeSwZKlVQf2dBTFxl
2XaO33q7Ds9jLWzTCK7YXtac1vopQYLhF3lSlaQjX+Lwa3tdMl6prJyUR0XSIdnqWyB5OSZi7NBe
WFNrPTPNqFPhTbeLvCgIDeEE6bWCTFVTQEMu/qH86u7vqhdQjIbtEuFYScuoV0911l/qv69QkY59
ENQeXJqsLT5HdDGHBMTlRkhn6Jykbq2+W2mKknapSP8Otr4y2bqEaaGcuoXV0ej6K24lVtDv+jRe
EfzoEdgh6Jaw7oUCK4YZCs0qyCANI2jvlWDEyZ39SVI1tlo1qyYtza065d2kbsOm+ei45urh5ZII
APkVC2/0H+eIUXAgbiath0RzUOOMolj/WXAke+OQMccoBC2liV9ezBGQc9LTodaE2la+YT513MrG
lcYsKSnSTxbIXLo4fSx7bMgw6iUHZZaCm28hQrTklz5OoisjlcH35j3N+niSfLflturizd7Qveh2
KaQAnN1T1m+g2Vw+jQfarHvUm5K5PucvoIi1L4RBP2VkEo8yPBN0s9dHApKLZAqbhI0sPZYIlvWl
1MIIAxCJjs+qzIGyjJrZmLDDsirGsNuh2eQ85ZKPQ7ssHYLzph3v36GVPZ9gpMEOJ3XFc/kC4IEH
8lMmL+I4pVZ0YGXOcNYvRqPeSjELTJct8hn+XT7fkpRj9xqbP3xJHwnPh0xFgM7ChVCRmR1ZLxOY
Ov5Bab4+CT0pG2Cv8txy9mfyEKzp0WfEImVLLs/eOTQ4IKNTBQenPfc6+gLEFMJQrEV6kB+c1nO7
q6P8/KmY3zz8FO58qMss3GUo4V4WEAMNQEt1OhkkXsOAJ+G8uCTpCrkKnbcFjOye4ptw9h5HCFZU
qEuL6hww8u6c619qXnMqSpNbdAotzdV0xWrEOwollGsy+yvVERwVRnMk2eviyf9G3vP0A2iOJ7z+
rjDhPA314Fc2Lv+4IXXfLujn1qMF8yiLpdyal2oJx+PlNPDxzf9DH3BGQNi+6ODedsz9ZzmArS4w
h2876h4DKeo/Y3YayCxCtbpU9daeXL9z0oLtWnniqB/6RCLwbKFjO36NzyTOnGyFKTHNvThP1HGR
Xpf8oVuJeB8y3DPTw7FQABmeQd9TVp6qP1peZeyzVtZsTmbfSFLcPvlnrrSuSIZrhDPxukwhJNrr
eOOsCS7PGfQIgaYyn5snsQldg7XJ9NvLCQtXLm7mpJi/yapPB19eBHxuCYhJgLWghST9F8sPUFoH
sc/9Zfjmk8S5nL1alIifKytF/nF2/7aSFW+alpUHfawswPmP/45MZXsjMEDVMYapbvRmHTqXFyaY
xMi+y0J4dZ9EMcu2tYXfMjT7VtuXjIvXJCzSapWpx7XsI8urI1xkC8QGpVpqd5wlCA3N/FAOXzC3
5jU/vL5AGeviHhJOrysrNGZPzi+tdk6Qs2PqcRtNv+T1esq+fRoe2boLDzSsBjBiWFQB+BN6kE3x
IdIAlRji7co/oLIy/bPrgmtS04idSzezJjN7pSxta+abFS1ungY9do9maDuYwXEC2LoMsVFBIYpJ
r8AhXcnn86TjCy3ect5Ys0a8DlBkCezqYTAgLX8Af1SX/9Twc3Z2AIRSFB+ytBGM9jUpN7XpGZz6
8uWsNCbznwzqFxpxmuZ3nEL0iLOnnE0bX2lkX7RhLi5yzIBcyRi7xPqcrIE+FE3uietY7ocfz4kZ
0dBzfsfeqBlULV7TdylwIKKR/YCTNiWEVpwYZPGlpCKFmAg6cnUmNLAKkYUyO6A3bRiHa/fONYtI
DhftLJ1G3CqhamcroyyVifoBPxZXQEV8/gY5JPkMKino62hWDKVUc/X+KXAHGi8a86vs3jn3eR9o
fR4Jc95x7eExaoslbO82Z3gTU9gIeI1hrg3jVBm13FhsOXAhG8RuknIQ8/GT/69Iep8b3wvVvS+z
EJl41OE6yHRALNmQQVb3S7O33XGTvzjmQ1uyCWfm0FXTI1I+CtLKMpizRc0lkOXlwjaYpg94NL6U
xbIIGV6cUponqT2zDrSmhQOSObH2acK2kdGTnxncRjhz1M1TT8VQlZNK6PQDxQ7RVzjnKfbhUarZ
F8PGgYEm3jsdtrToJzvHS3wI4P8y11Y31lrOSdyANoCWk0HR6gV3qT89tDPANfKM4U+Evfqn6gPa
hHaVI244rEwK08Ho6phDC3tmbzPGRnSx41WHLCqTLwoX2yRRXc0YUAVBKA6y8ZUBwuDms1lkBVho
8I3zi3viMQ2h40hlwwsov+EGag3V4Ak7rpKtB2g6EDWzOt/OkLsF4GjGbsyha7HLYhErWWmyOEOI
iy5L03VMbMjydu5K61AN2gXGNxRu3MJk6qOZiSiyb5eXu/f8n6U1/ruY5rVJGYae1GX6Pjtc66iZ
PFekRrp07AVTyjHJ3xRV0hzTsD6yRUBNUEjVkTgb6je3eiP5umMUyug1iJtvz5egxVxNMylPdfPC
wsr5yQRT4G6SZ8DJ8hMITvB3XDDsUqYawfflxF0XCI2iL9x7b3J3xzo4MyuiGv2hdSGI767uGrh6
f5/qJVMv0n7O/8XMzv79ubJryvQbYr4tWxwp2OG2wYLmXuF2J28F5D05FNjUN23PlYwr0ADFMnZs
1fIBBMSntejrB0buCqFSFTdllz6psaXj1rJp1rbdpZxKncWprglQEYFc3F0xEXmgxENDPxyRXCRG
drcG2uaq4XbpgK/7HYRzML02gKA0eY80bXbT4VQmwx2kEGTVwmwAa+cyHqqGPb3PFqyfarNgfO46
XHbvc2nqCbx6nvoW6TkafnlE9oI+NorvgOBHiJEQKbZQalLtgNrbngr5jY5zchqU0F3pudpXGN7a
KLXh3DXfCw05TeU8ihr7cTgMkCTk1C7XhPPEctjxcEBTTzxn3AebEtrTBaPGj5FPRd6PjDSVywHT
QoDgBX8cLNcTjx5h9FlXaTgRlWYCLD9vc73NHDQv9jKr0uZnmfhvKxLcH4bR4ITyq/JtefyBKgrq
kplCpOx6LQMv+J7pHe83cV3fsD/SjVg3mGWiyZf/UeYXHpbZwluL8KhzBSzhgLfQebheNYr0b5Rb
CK0oK0naZyYUdEdku0tx4eUn8foI4B5q+g1KsxkIrYY2ZbiZZOilOfx+YLsqSm4ZRtS7TBegj7/V
OaxzDHinyiIKT1o+YnQfd9im5p0j84QWnVXhORGurFsG3wHMBVXprU3RTwcHG33lwsPdZk+ra8Dn
h1U9fCmQEIeywuUm07Mrc4hQxMTNFeNGju9KpZcUwSRY2Z1W4ZLA/3hf8Rn5eM/tP9Ey2Ri8RdlQ
vWhSpXUSLBXZIWF83juCv7toa01rogPtEFF6xEbVdEk4+mM0WHxvz66ottPU4N5Gh8jLy+pxH9XY
6u2/Z26kHl8Zj/DVPQ5pTQm7lRONW1N80OsR4XeATiB1q0ELBBoJeOP5aWc/tWzftkXiHaVHgPQB
fmZfBrXvE4kQBHd0biUaIPduz+34s7mEADE4EA+r36Wdq4PtZT6YSqGN9D5RhLF5fOhqF1WK96Mh
vzww7lM6Bpnrw7XAA2G+yGB3VmoY+J1MSJhKsxAqsQFcOryazBmGkcmfIdh4m1WAEalQ9hJ77hsa
iRHqDtffcQHq3c3Y+lsdIaHORQTWW7sMrfFXBEFEpKVkUFYVUBlx+S0Ix6cJkcQpiefp9Wm086Md
EEXijE8AWWN8RXbTZRQWmn7sqGduwBOb9FJKYkU4GwL/oo/LAT4VlZQ9yfTk+FJG5znPR3n4UFFm
WdTuhxgGK/zmDlJfmx1Ud/Vc8t6+98nQEVluUxhoirrMhVyX4jVBos2gYKbmcjt9hh2lN88CRRB1
TjpPD2CPYfu5fjIsbDo1VlugfZ13ZCC20QTFgwtKnY4WsNN6vcGTXPOxETb/FEUOrL5X9N9BmXk8
fnYRROSS/gQqeY0IkU2Q8ImIVQFhUq6k4UOPqwW/bYn1Y+pDK51Lf6XVQQykbo5VYL+VtsfHqOj3
GCocJIAukUIRsr/arXr4v8pifoYwspqoeTtiJ99sKEJaajknkw9z6VDJenXXur4ySf4CIb19pLlG
bsvqnkhv/fszd5Fh5pbdH0Frh9cqntM+WLLuORfZIHoggDo/1U8bC1/R00tLbTUKNetiYznpmkHm
MItEv1a71KHXyWhg4W2OZVLvmbrW3QmSoeoue5cNXCSkH+VbGMfm/VGG1pprLuxQdTRmCAys1FKc
tO81qog89/e7Y6g5IIDYkqes/DBC/U5uSY69LOAjOv5H7r7Sm7qVA2jP0plvNzRPiI5w693QnM1l
qyBTQSjYXJLGWjVbJzfJndgRec/I0DYrCL2QJact3M/C8/PaUeEsFzH2xfYOb1TZHoK11FFdoMWX
yzal+nrFr+cQ35HPQhKjqAQGFvCc9UoyRoS+/cGe/LTwaaMtMXVQzKg9AHbOVDCmMl3KxhoGYtBw
afcXd26Dr7q/z48Opu/Ai6ftC/nd0FsEjkVqnOi0EJYcaRac/oq712K8iyEb+sxXbJcgF45E82tO
5vmUvkzIgvUUrAb7v/kZttRN5Va1W5/lOFpCSKvKh4QtFFbzheWM+8zANKFM5bKHzE7OlDQ9flRt
ez8KRQyfrKIASsQC8E5l9F4k/8jzCrsNt23rXRsYznCchkoBp5QND33jrUX1JAxdsp+TzrqGxxYy
J589f4NsgC8B8VtVNpxEgI4wnxDgYhhcvlqNCMiVASHo3pTYZP1AAYFWxV63SU7uy9d06eeIQ/Rs
ToHUlgh+4RWYEZBPCvBvAsmkluy9MsMMiCxLLchY5TqBRObm7aEA1JACkmbrVFcfd4RimS3e0az9
QyM8yxMDd+lUpiw1ORyF5QNEhc4FXeBScRKsSMZC48ovqtlPvuUjktTQKiHCuZy2KX+Z0m/8JePA
szEYL7Qbpz9pSGWgsqh1awqEuXu5d64PXKjamo7wf72ARWUcsKNIYWH2LfmTJFveqcnQiVg1WhBw
Qd0Zsq+laEWsXnyVQahVhTJ4JblGWfyDqECaiwhe0I35B1NpfnO9mHxNILQQlM5CzqmOOQbmdCck
Ye4PsjkDp7gazDB8/mJTj34iUjvowif2eFPTCuMIguVZJGwxwmeUOEf9EWOI1wDmbXtyZcEXms16
w35XPbaIYAOP425dE+5K6sWZ1fjg9+9NItnSk4s0o4IF/gl7Vh+WmR0o86/TZMrnnY5ZlxwDDQFO
b95zZut7jW8dENuDoclOdCH2+Yh1wdPZmm+WZOJY0vj7S4c6tAYN1jbLUflm60IWpXPiR7SPrZEH
flZsudSLoKIy7KwNacjjjTOWcKiQZS7fZklzxYOfOAG/g2Rl+qquVuD5qaTKfOnkGqhnR0jovo2F
97F1ZmtDD5oXqHMFIjFWMk37QueSJnV6eExJHYkzopS0AgROS371Ie3Z9cBEg/eWa/G9dBru7N0d
D9aMRz9TjhN+ihfGodCDs0qTk3zHvVmEnbx1lgbfTOXKV+eKszahP7M9vmsSjhsPFiLRNcPJ0Gsb
QCwxioA84B7MHXyqq6sb3MGkP5W2+bGpL6rH/yL3w6Anm8kyjpFH60mLT0UWKUPGZ6Uc3ayVG2Ry
FjsYaIOoGILCYEyuw4Spmt1pxORPm30zCzhM1bRHMzNycXNlrJUdl6aW+kIn6irdJSuwsUrqUfif
ih/hh70siMNEHyKo7fbZfuyxCvSuVLB/eTdvBTEiRPs5dpl9/iWG2+NSHIep7i2S/uIuj4iyKOlj
DwHmaDGOx6cTCBH3BzgimMaNM2/ipSDPfOzQWGILQnXFV4R/RLsuONTSKYzJHl0ZXClBErCkN4A5
tEpn+8KVKBAOOUv18tFLAd3i8WH22erPwH5qPZVABhp3oOuv37+qv74cnjUQ/pDoDRPgV9yhcygK
FDrIBj4BoL/IaV1ksRtKD4GQDIyvevIJylCcAJWC/XVs6Wo7lsa4eGXlgrvxb1gi+XRd+BZqvHcR
e7VeWSN753uUuDV08meEnC2sgoDBZc+nEycegeKJjE0daDCdkNww8Dx4ZsBcWMfED/4Qj3A9LZ2C
JmO4sWcojb+tsTVXkJ9TjWT3qEZA6FGHjKvgUnHOTvZ78doOJ/QTCXTC8TLFycS16by3dpYKCy9q
9ncC290aUWLwEjQ7KTmG6ALUesnLN+eQc9NCo4x4LMH/5okuYE3G0BRBDZpfZsF1SZfXrEszyp9d
zA8IsGDHVIyYPyaGfWPllEa4pG2Aev/32WIskCXbo+0g8aEtN5fKWnB0l4xRq3qfzMYhdb0hcZXW
LyQJCrQSz7oPHBgHpJPDAY58Zc3gcItYaTxJZ21fqOx/mf5HVo4rrd7w2of3gTlJXvvy8LKJRU+b
fK4kR15TgqrHwlDtQwgqI1/HV02z+3mjIEQnr0CtpHkNXU+pnRLw959soTk1MFbVDz8FeXVkNF6b
XYoprJtBUC8rPdhDKMyWHfPeKFKw4g9TDA2CdqLIYofMqv4VMOS8MwWJqFzaWK8X6agyzWOuw2us
aWWBlru/GbKbsYPj4379/c1w0dvjo4zJjQFB0j5marGk72k3d4nFUIzql92N4vglAUpowOEzxeRA
pOjmkvFN1zw4nbXkMBwrQGgnxrUWrlveQrr+VyUAF7nPbKCPD+LJ5Z1XqocwDV6sxyA2Jk+Kdj/R
kFiZsajRsxVlYYOdryKeP9NxWceKy2xoeTF1McnxGxDVgOnY6XmUTcLyYdjUoGRfL9d+PPoG0lXV
srhNnQpBWuUhqS7Z0KBeSN2d4AuMUcFIIKTtrTANIhEHpwg2QUhuoo9WWpu65QmPddjnFXsQn7RR
BW/PsdBjIz+hrU22f52Gf2HmGAmb5AF5QtefnptvYA5HlrLfWbi4QAOaBWVZ0uYUwxLz5yQtXUPx
vwxD7UJxLZmEU3WzTHqCGaOwcS41SlNzC+05/iekRsNrRJxwTB3j9LYT+OUDxsscJjo2leXsKu2M
ZpfW38JlCfC+d2hdna3ExTxpJroLAyv5MZ83xoQ0iFGMG8o7Q+5UhmSvn1P6oj1sJAnoaa9K1RmB
srgMqrlYupIipcD/JJFXr7kTBBxI2VV5lPHnXwBSVFJaC9AD/AA+ofLVQQykmafxfkCOIj0X7tt9
cap3J47O5XFpY3Th1Oajh9R3XqRU6TfkEjCYDQa/eiV3DCWCSyE/BPqUz+Nefs3Epd0ZIb2oPZqw
UM/vrKVStRVaacz+guuJoaunZfBgkr70vr3flXAMPYHDp96p0OWuWaxmGVbcnYmYF5qb6EEozST/
AkChE6uKoKwunsWWpYh78lwAt0WoHyafP8i0ZNy4G4gMH2ajxBPwPubhi5s6E905o6S7ks2U2Ngc
beH/z42x8NL1/xG7yJeRELIX+CS6uAPo37qvwEF8UEIZPGz/Vc0s4fvsye3+rQDtfLwLczB4zG2P
FV5MFiaKctQ4OpPlyfXW+/C1AKdtPOPR3wctE/w07iMIbzl5Pt6boJ1Ovb+ZPDAIf8lxyqzwgb5w
YIVyGgXgIyloG0xgsNt0rn3vvFT/+Z62RQnqyNBgva4GWImRlamSCESOviakRVjC//aLh+mnHwl2
ovjFEUOazQId08YUyG/+huxRcFKgtTj5cwGVpLlQlXGVN9VyYNDSH453MbcZ9ymCh3D4OeGSw7Xw
437yUzPlCbuG1QezTinZVd4RtE66Bf0QFHkeZ1ut4d6pZl51YDOVA5U5KQ53HB5UEI+WgtgWQ9nN
JzwBeG0aR6qfWq1mZlYCM9PKtvkhEmk/FqcGUrvoVfh76L8ylk+M4lVrtLyCirPksO/7N6pCM+MZ
Ef14PZhpBewdLlWiIeHP7NGjvH9mCDIyc16jzkU8jhb1Z/uFiK+gbwZ7VhtRhikvJmyJgc8lHFUF
eO22ciwXxnHVAHzCHWkLwZNp+EC+f0arJ3nyNFwGIinU/m2SP8XgpgKq6bXUtBfg2/PfiVHcdZKF
6pBKbPuXAYWq6TXD/fDC53c19oi9o4bpzQ63gtxwVJEkV+eF1W9hN9gmDPDCdw4jpzTNpzQSvj3h
5qiCjQcpQRUXYvHekt7SLjQHm7R1Vbz40zbjSrMjG1tSVVNHfhKCzRG9BAnCMZseGlDO8WaHIdPT
ULMmUKwDVt765idr/iEs2prkV21R6O5pZQL+qe9VJUmIlPxhTLNOLbNxrwjFncKTpoyUlJeGxIwN
r7xPHTqW4ULltzhgl98eomllkHrBLGpIHbUjvMkOrsTdTXmkMLCI53uqupX0zYoed3x1MOwowLUS
1cIc24uuvYxTCBjONDwDzpi9uz9Tkg2iUv2h0KKP7KpiWGLcH7szoPrCLdEro4F5I+xI1S8lIDrf
H0TLA+s6t+UyX9ec37hWoTtc7adjA4raGUV8BM7MhglGNcJN+uh5WHGGv9130kcxswc9lv13wwKA
JpJ0mDDttgal77UW2e60bKzKsKYdSsy0P1NbPHYQpsU0uswR5bXB7jKMuLgtyuE+0xAhp6suio0z
mtzeieUDBOi8UNaVX84KJZb3ZIVLQthwPhNy/0cMEhcRCCL4GEVQ1BLvS4fen+anS12r7b6nOH6x
qDQg3V6q9a8SE5e2Nwj+0IOm+n21UxtlQJ5Nn1xjL/1G1BHmmyMuHS90OEZHksCGo4J6/volZsQp
7Z3o/3OVvJv+fSG5c2IiGYLNFxd/k991KAjuA9E7XOV1xNsmFdNiN8IvDB9BNZf1ZSGBw40oMoxg
JjdS1MtgPjY8AnBw2Y6dZt/zKJwlmkLl+2A0wC9VOezMgVESy1G8xLlpSohDIIghH99fv4KTxVmk
QWU5hy8L4tsVh1Txv9pYExqSiWaCxhbZa21n84m7fbAxQJpm+nJbVWZfXg8BdXINKZgi1GEG7VAq
5cw+ptUyF0LCbLb1ZTIuKfu3omWO8mXddheK4KbSrXrLoDLfCNP4n5L1VcR9QHwfQJmbsXyokBdQ
g4P3uy0Q6vaWz9F2vPy/wLW30wwB1GUyIxsv+RjoyVISmIIC0H+TAX8YNc96IGfloYE7HDkDGybM
CpZu6VVJwRW/6H3T/GG5GlwumlwmdTzPxJADnQTIo5VXSlassiPfgj2SXn5CzE1J3WU7uep8+HDk
V1Ph1AfxzZKkNnEuhSzYdTtL18ZOLf/ebFtnWb/dp+QvFnkSAnXqITiYiXRuqAFA0cS7AYGFDZie
TN+1MMgVZ8Me1jVyxZqmpxAaPtkZN/jsHNzSYvEj9D4Bz9BxvgOJA9cvo+foJF3Q9fxvH8iRNo8I
gXax+ftNfx1XuAAsm4mF2sqbzHL0Lrncix/oHNtnZ+6i5xXW1Dt9LO5B9oZLLkShh4pixicaG265
25+hG9nek7TGp7d1TgunxgvjtbAVoVNfG2Gl3QPeOmaeXp4tvft6iuyq4F50G9Lt0Tt/AOsMpg0B
NMvTpxkUs1J0Ls/nrWslpfWFOIvmo5xJChR0QAM/jipsQjJy0BwIRMUGrhv916Kd0Nrnn9qn9h9Y
csTP156R60+xg/58P6e+WRpWNkASjHk5JZ2sxdTOC1ORoatCSaW0J31X9SJ5Br7DVNBHx0ksUB3J
N9AM0NhciOWRl/9MNAPeJy/WxuzxxpEJ2Gcmrjz2BkDxSEx1dMFZWkT5iL1RwisbRXwCPkAAnHBp
gGbJsApdqtCMGiC2u/b22aB14D/8ajn9ouJAXMlqbsoj7nHQ7oI3a5LDqEd4Pw+8g7FZcud3F1NU
2C4VG+a5rCQ6QDbYeEQPvyzkgfOZ+yz04V5IqONO/4UWFqH3OyqdGlfQaFxYI3Qx6Sf5t8hceNzO
HQ3piWNAebIDumudH7A69B6hBjNknPRlJydh8fodobdm0U86JTDuAsLSHTjBLT2i6oiU+URWbg/Z
6Up45Edzf0b7n+fbA8eJiTlaZlx8IhCBPO+JlogcAE/2svFDKr8AAGH7knU0L4Go1fGELQ/I/i8j
pZ7VavL69VG2NxiW7m/Mmw7LZMjdNJfp/5iLwi0APpfwoo0qhhh0fQjF/ZQ0kGmt306it/GVMv1e
JXCMnuyu7l842bQsaImVuPEX0VLL1WHN3Gp+/tm1C636iQrs73NOfzbkam5zzv9XD4IiFktsgykU
Xe9fc2Ddmnr6kqeHlxtbIl3lLxouxBHXMh8MKe3MoQySoESSySY8N0sQQ52Xo6kVPuZhQtJTimp0
PjhrgkXL70eOLxITc+yxhFcR1q1QW89j3HaOPDBme2P1aaVMi5zLh4qMsO31KzONteledQEZjgvP
7dL7bSbN9BV3Id+HTsKBzAk4VlsNkfQOMTL3tyFTjz1+gOj7MvSocIuUAndVOuL9MywMc3x4jD/7
K4aM1v0/dNXDxa44WdcKFK33n2Xl2gGX28P++KBrinAOebmlTTYmDCevygw85vcZ6C8/ZbeiNPyS
8JalPTh4n66UNSYnrA/0E6qA/TI857EYhDixWoOH4gZVQSfb7qvyGOQmDOKftD8sZ8PZqI5Kvdva
IDlJjlNIthttm0Yg6QYNoecUKDoxbDJCMLhUDaw069EYmf+1qF/LdfJsz3GPfSCJNusdZBwVYbJf
L1PeXiPagqeawmRFrmAxnY39qpSxCwxVzeQ/dqmiqRHPfZdYkCrvK+fxSC4Ojdvhi1cs2LdhdOXt
+MsWDN/oN8G1ktbtrsLuyTLFYfFI4ZzYeUzI9+QE5vvnRvTfs/VuvFicXjWRhaqOA1Lm1Dm4Y+mp
CKIUWGq/iOsmrMcdhcMOUJoGxQDPjTa3cPqSVDeLWPcjJSxKPanZGBC3W3Ni87PMBadHyzwJjctO
gWZs2d52nzdVazDVgg2PwgPk+tYxGLFxMWowq6AN2Q+lAGfNv6udtKjaJ1Z0tii+k++ItPBrdPtC
CONo9XoBdC7d42t4XQ+F09bVjLGNrV/5L5u4sHRKI19AL6bH4UGBwMBZSupQi4rypNVDZIr7Hmn7
rmtI22CniIA0gYGLcxwGCyJj+1gtLp9qv5zZ1ejDhYQBz9LINaJcmWLotEIQ44Vt9oYE/mlQz2a2
8YLNl4CML/QloKHrW9BGU833St2qJ7ePI4EGpMetxIN3uE+hUn3g6OAcy6PmqDWvxOdH384g/Y2R
JSrLrs4VtreXnv0yyFhQYmF9bGzJOESAYoGs8OIQ5hhci1/XWU9XrapDLqaKNusNuko51k1RgIk8
eWY+VV1CPC/w9ssjV700qHNq418HAO4aYwcKz+R3ZVzFzaHbUSpd0t9/cvNlrt0PB5HF56JeqOUm
pBiitY/0HXhgp2yRcwR85Yx1/l9Sij3jl1LXlJz3jVySz7dzZim4FrDmBml3zskMn5Gk1fx//Avt
JDDjCO5tAoOp6JUiUKS9docalt56f7G1D/xy7cHUgsmTDhCiWpfKyy+dPyWnx0EPXnHbzXWot6r9
21f7U8G7j3eYOmyInpbgJ4gpXxzAnmuKJkgkNMPstJt1XJb8twYiMJ3fIW+7hmGestjm9CxPLQsa
Z6uYAULnboSZAZyDPqNkMg5Gvj96tVxuYG08fDjosAIj9Q7KVIdMTalQXfCT/qag0WpKxyV6GatH
RUY2yFPjDmAZ4ZiZMwruqCsqbxrnM+xpjvX+9ONkG3SnLvfY10Ui2RBS8BabnhYvsUkJaZxETkPd
xs4hX8JBmc1r3CX3zSHUXwiaFxywWc8E6f2RJrE7UosJ4tgKXLEDYwNNw25DU1zbLYEUzn81jHUz
Fy8IYPLK5asoTe5YNashJHaG288LKLpoDmWH3EqkoCnqcGpo5OR3vMPiwuHnyyhK8kJPQXCeWiJu
3IdjGM8ZEMWg8qR73Ley7vOVGZO/hEeEvyYB8QjcGrGVd//qbJojqnzedGvXyCv/w5zAahx2DRou
aEjWdR5qJxr6eMdSRdQN0/XnJgtSEbgS164IBAQVd4SQB0xrn1k7x4ej7lre+VHLzTNoaPNZ+wfE
vkiz0t8Vgqxw/U2SONE7Wyhe72eg+IQlM5x7iWt8LCmlRrecBdAWbibQQBA7xiLATXeJ3dhhO5RF
8fOkqRCbdaT70LJfBQE+n2KHehf0bVJyekjSGxCf3rUS4X6MN7WjHZnCFL1UrPbKWWRqUuCbJjAo
3mWVDxxS3G0qr+VTMLBPsIc6Ev1ONJn70fHh35qYuz+wpms0IGiSDY28IjrVnFMc7V+GwoVD3aic
suThAK94DaYwwOrvz5FEbdPMek174IBmQhgbzVM63gmR3FUz6L50sS6KvASSkzAL05Py435XG8p+
vDHDPv+McaFgFCG+TQwsybwhumCpdTfVNpOOY7TdmIFngvH8E7z0vV6qgJxmr7X4f95Rx5bGU7LC
HXXYDMIzxK47aqxxzk5L76EvIZpYwRU/b1jCK54h+1iRq7c0+u9f6GohP7D1pby5FGBqbRnmd3wH
II7NBj7kpoQEX/lnGmYHaPEzHnKOb6VDpb07KTXsz+inkoMBjSOxqyggNEn7gZGsOAu8f+AuwUJB
xjl2LARXwERRbRopdhN/M4bo2W+VTRulbcLe8dJZ3QzbFL6ARLR2yyKNxMqhYDQd2HT7TbhPY0Ri
hcdzzxfSyoEQUHoVLae0KJryO4efv0Br57h/blVOcRaVuTKZrKBRa6xn/zpg11Ae5AXq25ZikTlX
gMkh6v9z08PtA+IIVFMV5rAu/WPEsg80XRBhbqNR5fK7muphURGceYSNX1tp6HgXKLjrxmjappO4
Sa9UwaWw8YxTNKc2GF7i2hLbWdWld98OtS72qLHA04DfKOcv2Tiaj06UhVEhIx//3k+vtLUYQbfh
3MmC3I8cP5DLah9LHiOtFeqvd/YZRNgRnm7Bc0WsQnj0ekc3EwmbBxKnKdnckVVC/sNCFDgJuLjG
Jf+qWg0kIdlg3nc02zEDRkfN+3gz9BS95u3CjXtJ4cMgRwd8rGroIOpy5Wl6rqQNx8nQ7mUSKlVB
iirbPT37Cwo4/zipjDMga1gAoe9qifEu5n2ha+oMXLxI+U37zSPwCjmYQZycJYBPogcap8C+eEAN
vX480fgzYwAGAjQNe0CutxQkjT4vWRsaoWIQE1egtW8fwUQj4GFNe0cngY3pQAoxNGiGzV+Xrt8F
A0WMTHhJNH/6xQqBUTWo/zhg/REAuqJYg+1G3e5NIT41mK5JrBypiPJNAPjNVTtndWJe7t1tYOB1
AcVN2eTtKESka1VUd2TCUUck3mionep04DOlK+nAjcdMXqkp2c38vAsB33lFK/fVpE6j5g5Iictj
oZqRadhtPS+bMp47FOA1flIRWMkAKiHwhq8M6wd4ExoQJlWILh9W4ZR7NEM+dwPCoH/JdKAoDe0z
vY7YfD7wG+cFmWo6fpoRmnSeovyQ5sziy043xcYf7/kX1grMH81jVwHvkuqa9i72tqEvq3KNd6pz
c9hADaQLi86+ZY6ob45xRCRGHK2lGnzgGfM/pp9F/ydb+HpocSfam0F97+jfZ/uYwsHl/5zdOx3X
4DRCcDNvHXu3JftERpfRXbsUqg0T8ypbNEg08gbQhIu6sS+UChwE8ebb5qv1Kx/SFheynCwAsGI+
zpVKeVcpzEUVpN62tCqVjK9xF2Ga4IjiRs8CS8aQd9oKoH+soT/3BVeVsFwLKApmDFBTvrz5gyAV
rVBng0LHtO7e8YS34BEjoh0apxD1JQuibPDn9+suIg2hb0/zV11rnSV5dgStqJE5BBAl45/LD9PK
rV8h25RNlw79+QP+hlUPuR1McHARW5wVw3Fj84FkK5NuC9XIFyBlaDxWlY4hrjMtlbTCzJzRQask
ODu47NgEzSUh2+Fo4S6RwB2CBv9QDczKOj+Im5Cz1riTWOLMa6/DAHP9k49WV38t3wYLtbAhYV4U
ZK+VVaMV/N6INW92Jz/g5adYHVX4MqBsV81HWGo47i24biNaGnIS5LGtfhIXF1Yfe/qcWAnWDGUG
GyHTQYXAHYDoMMhh7HMhxRcLl2gHaIBbOjgn/bEQcWxuU9isKq0tE9UcaD5NccBYaeS+jf+nQCyV
7gBnFz+dAvyWbmqlPD+NRr/Ysqo/oty4wl6GaF04FVbmxjfiBfSBfeMa6nTS3Ic69wACF8REStii
MZ49BkCjqbuo4YLyPj55M1n6RBoMM9sShnYU+VT+t52zGOWnvv1hkqMDyZjilxtX3dNjWVJtTtkz
pIpF4AKjwcKDlanb5aiYBmdJSudGN5eRbY7bbSyYivLBFWmapim351siOWZWtqlFBmbABrmoVHQS
LJFWzaOvx/XsSOX0wvk/0Fg5HL1uBs19byuydO4CpsAGGipWaHpxL48jLdvigaTeoc4afiUNOW/l
HSMKd0rmPSqExFZFI7vZz1drDjpY1gx5+vefe5iBKtihpdefqSRqs9vKihWXrEkj/V2TjSM+PZ3n
GJEWpa04QVT6/DKr4ZKVTasucpWcxlRbY72uImAhvLIi23aF3rfR33hHoTOj9JXPYm1HF8t404X2
h1rsAURCil/+U3F7YTWZCoR6k3jNLdFuQlPWlOCId1JFpZqrfNZsW/8RcczSzXx0DARCnrxq6+jK
s7ZYjJokliazB91Xqft/w56ntp1P80zk2Q9Z7vS8ESImqq7xQBShbokTIx6vRjBUw/sZGtPIG3RK
fmZyZGUuB8tRst83ce6YnN2goUlmiWsnIc8WQvC9exqv6owoPX/VDZhsU6YsMJmVEUYM8MBAGBS6
Befj9oJ6EjyNlRsmy4YQu7C6aWinOpPH58V/DaRWynZfN04Am/UfZpXPYBs4hue2NDIHBNCuIZLu
owhFR1OlFv8L8FPwUdEeVHSJEXWxxlQ1rCBZG3yXrGaYCFxCutpCtnzDmNsuM2+9A0763zxw9jCl
184AkfqfWL4Aq+n9K+bN1P+tXrM0/WOoGjg08J5qv5HuZlM+iTpFKhs0kjY6hkIaZbxfqdEJ46lP
Uc9z1uVISoa7OKYuoAvEJzK0ibOwobpcgNtUZjO4ocofVBiufk+bKS7nm7wQUNbiG30hYkEQ4G5g
GLcYgyewXaxlREiS7FmJA4yyHR8mKlX3V8QzTuYvUvEAns+BhtjnraOSy0nr6wKBfMAh71yVJm0z
NJg58SJrbSGri/80hRr6IvMgRBICgjkV9s7jtemIb3rFCytCi+BkfyGeUv1ukkSvh9Z3rwkVq171
SRdAIHs1DIsyqXLfS2TMt1wuJu0iPNLHezsK4BRFLQ3gDLGgblsQKnDm9JqFUS/RfPxU4fmAMyYQ
dzQSDhpnK9pAlKBJ9+G4lDGuD1ufPmUeaYqoR3x7VohqO/P2LO6S5VjO30LzhpxS6jZXx7Lnv1xI
o+DfFqFOdkzdne3VlJn/uyuzhzIdwOt6nkCmmAhG1lkT43E+zdsy1P1FS3uxlo4JnALdRNTHKr1k
d0Wc5hfIQfklkF8XDaS8TM7R2YcqEf91iXNRyjlGKRc5yHJTd8UW9wXigBQL5oaW7GNH+Tom3ri5
O7gzSqdJFBHfy9hC/t1yi0gbPnDLobEqlhSm0belsV/mwYcXK8w8Ic4QU+kINMdQiBpgzv8pVswv
0cD2/06jFHuxAqYlxfZ55qz/KCvenmpfK1J3IQlKZWkwYGGaWSaxG22xoK5fL8k3/1dsOW78Eobm
x9VLJyJzI0VE6hMNrs6Hu4Z2X0O6HPLX7YjrRDMQoETn70NwvIhGRwgg+4JmcLtEA82FP87b2iIr
NsmerIzlxqSgC/yZihJ89leR9x8MuPLLUxQN0A/rEy/lApqNBlBm2jMv+IhFsRIZ+M6KBEid6UWU
1F+59D5/wh3Ak6MY/rYWj2WEYxzgYvKu5k9pIrzVCHSm3CSN/OKRzvzvERoA/WOMr3YHWntOobXQ
inHLrDDHao49PA0FsNOVniExnrNfbMhZGyqn8LUW0hXFTv64BUIHU5YCwBdLtsUzC37pKcpVNT51
JHo66HqDcTLH/o1AKTVDEbSTVusEu0wN5z/k6/eLM5phuQRi1D68jFOCUxgpOKexxMDmoV7YW3Ze
a5Px7JXWGLtgtSXF0VGOiry/yl9dBzq1VEZeajgtyOtpKSSpR/FXKUc1CdmEFmhAWxDfb8u0PV/P
u9Rd1VQZn9JhrGmH4R79N0rmUkqjOMKb3hI1rZ9bK+3ACQ2HOpk5OSOEV3cJf6cz6aMy7MHURHKK
tzlA55MhXV7YxE9LDCb2NPhqTMN2Be7X1QDPbQr8ik9pEg27bYPL0EM5Hi1i5TkKTptAPTI1Wqtu
nLpcdqiOwDqPRa+QS1i/noQejmPPOq/sVjaQTL7oQZqEODhCEJ5N0QJ7YHCrQVLBA2/BslAba5y6
MDyp6qeiEOHBhTimIBVv8z165ck1Aw6hJu4ZQnfK8i1RxwwHDBNinDfOXKJroo4woMutHjJN1UcW
7t9cw5rzx5txlyS62Ihpy7+Lt1ysc90/VtjG7xShSAF0B/Wl1w7kHbfjqIF86tybl+fuiVptezEQ
sbQFZnGzPxylarE7qy9PjzRMJqM7WF/M9LLVq2bfuUPhEJATBo08IS3GJayhaGrX5mAFnLzYHZgJ
ZvCRI3OWmj2fRZatmlra0VKwKg07rFe7GUmTmXkDxVImIs0BmGagw4x+JebX8LEXi0W67Y3BV36x
t7SrwZgI4iiwmpYtzO2eC764p3rtoGHFBlj+AMO7Kt8vb5bhjNrYYoyFfsy8FvLNtzH54AFD30zC
S9i2mzHd/ae8QTWRULTsznTIQvsX1g4s1xKF/EiJ3/00fIbrij8bZLAfz+T+K32TnIkla/RmGziU
sShGKO567gzTLZ317L9orilr/XSzJ1QlxydH5lhLmlZQbbBodsst1NMuwC6XvPswabsn4n5My8AB
zWKFEyvT925Az4ocSzGmPma+pK6M6dAPrAag8aP9noRPcZV6tjO27Awlw9CU0BZ7Sdjtvc4lXi7e
n0XNQBxTMJu9E/JpifJEjtd3Z1SofMRoWapKiGoCVjGaDDfz8t4lpwFzIQEof0Lvdre1HHCqdTuY
pLoWKe7vpdtAKRolV+tt5zWgQRUy4qRT3RGPpBWB40V7mbuAdZqS0+FihhyXJ3O9HXNipCSqN+7A
wqJd0Nh+2ufGrhZeWWfyCnL4mQKBRYWdLrCa4h+hSDe6VtXdiCZ3Kf/cASDTTxB68RDi+7HxcAUy
knxIAOnbEPLFajI5TkaAPY0DPjaOkG/XpDoCdcUFTEzbo8xQqpljlMflfgje9fWGrVimA2/n2XdK
U7zzZSygGUAtIJ5yuyZQN+pgyowdJvtRJH5NeyZndoi3XWc6Q7w4ay2Q/jeT1SCpQvZtxQQMXYlS
9JG8x853yPuhdo11NKg3jr/VrhGH/gC+hgMjXkzTnWBYTtsbYeqJ354IgNHH21Wz95kwe0oYdV9n
cRek45oKS54NzWBEp8/D1ti8UUuU6hndKUP0tHqOU5B5EKKx8nfyif/OYA4mbvRhSlPIV3eZ5O6s
WAnd4Gk5Wsx81NtV/ij1DXS670TXjE8z5YFTFTZjLjOoz+YHs1s1g1Bu4bRF/Cj0kphlQJsqzQgv
tMkKbS1jSvUbmiMAS0gOe563qISK3Si3opjmcaDg2hf00b7hYM6uOedm/yvxBngOfbtq4x1TdmuD
tHZajwXb/q/45dq6Z+qfFvzWXSNH7M3N/B7Fzat48hjs0u8Pqo78Pr117TwUPAFhugblC/53rfIe
Z1nWy1K590kwyLXOdm2BzINtgyHmmKxzgl7wxW8x/c5d45O634me+xFOHYdJYmBrIlBQNWWYePhm
889ymzsrccV3Gx099nGcx1a8um/YEy2wTmEtPTb+7FzItlTnoZieiS4XvEwyHTvhD/FHcS7YCIhn
Y1pEoFBpU5/mEP2AjMTma7fxi4hoKXtrFjFUjGGni+n6pKzwMnCxVPFeprzy0rxrnmrrGB+BkO6Z
tMhGMsQXhZM6tMD2TYAsamRT0gVaSrnxiPpD1udtdEYKS8k7gPzsh+4juHGt1ID3loJjUEqcK4ua
jlvWsHQubvj/mfHXh1FM+5S7FRBgu6dz5B6u1SWe/xZXN5sz/rki4ptYJuuufnOFUZylsFkla3ZI
M4dWlC1giBdL8p+DDP7BB885+esqhN2mkD2Wqds3eRH84Du1JTTfpUXxiWntU2jBYTXWsKo5wJRR
nFT+g/sohtzGzXouT1g4/KTh3PRp+8w4kTusbt3xakISl3c6Ffa4BHdyeCq9GiPg0qRC0DIaId0L
Kre15Wqqlz2i3Pi+x/UUHm9HTKWwBHpEWWG5SFkYRH0JQjKiNCrb1wsu4PGomOVePgupWkoKP38M
RecL6X7MFTy+9+uV+lNrX/eKqvQqZD0IXDU7huiUP0hJG7SNx1vFbIDIhDPUeaQi2kmme70y0JVK
pNvgzndLGWA005CpdYTmXdaYYwceW1gI4uRYHUV+se1XEpa71xZh7W/zT0JwKcB1hvBajI2u9Q6l
HXZD+IcOAbNvdgDnW66jA46eo+4pHUgs8QbBkZrrXXyN5iZlyUamOwjK3X9gUflXE/vhNcdujGOd
1/WIvhb5WKAx+SOu8AIlODew2vsNDB0KSpknru20amK0bWseyhLOTW/lFOXH5HsOXfNNpAZOsKeW
2LYgB6X+wWFiJoBn+B9ltXjUTo4V71xABOVjm6rx+CKgl2EnYcA/twMLV8z/rsxpAjv9xjPWqPsN
v0TtBU4SchkZWGInEvkA24UT6eSHhnQaBAiEEBzxteOhHOKdsaJm6nBORGdqRYKzcsDTRpJ1KBR9
I57tO74m215CN+KsjNIYephYZOSHDFNdH+zq5Ik3hfKTBxxs2YaN60vGIOrvg2zsY/Rp3rzbAs+N
mBZN+RiysO7DveaxNeDLPSTBbaPLPebVTIahDABRQ+qfCPK25SCk1StrERdWmNrVUwmrGqCvqC7L
Ie4t7OclwY9V7/cRyZ+vaMayHQwqHt0emZXgrPSxQHGDSQo7raelzWnMHsdy1btJBKXwN3FDM7fe
LDTpcKUgVkUMkBZaGv8Sk0uR5TrqvAe1Jw1urggGrJ7XGEDSqakDTB6KY5G5A1TjMH0SEaeMHAKx
6SnZ1zJe7l4DYq9ew8XpKq5QoAzvL8ye4Pg+2gU9oJFXuikZb2SHC3RgtCQLOwWXs8Lbk4tSBamK
iCALSmWFpDYEvzpnNPR3fU+R6y/wD81DhNdVBLWtToiaxBHxq9WBXWqZFYIEQgxN+DTzUifh+kwD
ZfSamE8za/7GkR3uKM6A3FeXzUy2SlVPW6F7r/u7MnbVMLH46kVG/+OWYXvp/PhvRG9w3OJyIpAu
np02dqTH2/7l9MKoQxYgsuUUMWCNkJtzBIuc01UDW3VGw40YqMPREtVRn2JGPgpXy0Hzrozph5RH
UGw0QKwN7au3tlxFDCXwhlD4jpQ7lMk98RlAGymxXTb4DKvWtHRnyL9FU8YyEsFdblk/9/T5ZFCq
m5DEuBccqHZF62/+bJBW+jrZrkYa/+u3IOKJd1HRyGE77mR90TeINJJKmHigvYzH0LKryFHHOSx4
h2tyvdS3/I9ECCeuq03QQSNY8T52SKtKXQVPIIbHdPLKhcHvnL3PImY37hDvuOM+z5Jx+YoB+Bcx
TKhntPMdzDQItRQvgVDXz8n9KfK8urXCWUSxAKCSXuN6rVXMkoyVakZlIRNYApPgx9BHGAJhS8pg
EqV3GS0jkLInDu88yDaughnRfDiQ2FSzktb0X2O/TjFBpifOvmWsNL7cxBHDb1Zm1pwHh3Su6uin
XM2KgUtFO5ANxOK+XraMnJzipbybc3+S1QLuibPEXd/fpZ9WrCPqX6MuX33VRTL7qmDx/JqUjz92
bnMA9OvMKfYh5eonwv7MYfuRoCkXUW0yF3AMIs9K9sZ/ZbODPJTara+TvBtj2iNMI2g5qzkPlUVr
BB1xnQ6D6kzMea4gtj6gQ+syL2BydCZRH2fl92oPpRDzGG4cNs84ib5x7UIy5XsYd5MwbZXXJQQw
y1tj3IQzRMB448htYf+VcLRL0hWN4MfnSimNM1RJfRKeOXAL/qoggkf0J1rSC+LZLcacQ4RFRt3s
er4i2PsGQ8tkcot9Kpbdxwei4sFijTuYSw9sec0vec75yEzxCnR9kRVWRh8070gz31SKuMNFqJo/
RdEhtpVX+mz3e7feBg7fEGj86X9E8Z480FdLXdTKpvNW/XGOQSs7Z4HNp52/xApYArUO7kuhkxqj
xZz0rP3zer57VXnT9Le6HoVcrS/1RU2xahyABF6zZtgTVaSBhs3JambG1vv3+w2o9eo8b+d2ACgI
rRYXXddWFwalCmR53UFOR9zAgwCdJNXzQHx+wL1psgpX6Ryfza98U7WRxxCG9rAiI2ZhviqLVQ9+
eyVAZ5je3h6TIsLWCvbpl1cMpErT7xClWF67pfDv8xGMELW6ZzRW0BJ7B8o5F1AK3MIRvUh28qwT
Zp4f2TrUrlGybOsjcPPNdmsiInoXzfP7gbxOd3Ic4PCdFWpIxm577pOeui8aLeuhk/7ehkx/GPkb
WclVOCiIZVBvd134F6lVuvBJoz5+trkM1kOaZcasoF3F8wz6gk7Man4TQL3cHz8jeOLDJ3hAjRms
RsDucxXPTPqQ70+L0s4DGclJcW44yxyMgZmQil7jjWlhHt9DsBdMHvPQ5KylCsKuMD/7cwIPXqnY
wbJF+XBglwreID6T4Z+YzkV5e8D+H17f9Q+qfXbO0iwZfjCO9mS3mG/ypwf9QVBGfCVBB06a8M+8
zm2Pa4oSHBi2p2A2IkO+bVhVkAL8lr+Ax6EP4RAeSoDrXhQHHXje2L5vAZNv+1Q4TGsIEFkV0hT3
LgNKxII/S3XL8m9qmuBYsC3hfFAiIJw8uKX6wz+xWb5hUFXMnH20nANAJE3sP5bN8EBXTgLuK996
z4JeLAzevY6nTzUVpZNNktkxhZzldlUE0LtOfinVUT1QouU8nSz33LaHGI9YWkpp3dsCzZPh4BqA
ySpXhp7ys8g3+5SA31tExHcRbBSpG0IDe8Z3FAz32uCuqw1rV1HuH/v8JAkdVQ1zrs4HHXflvOcl
hoDn7dywx1SDmX1aAhi9MWKgWqftz2SZ2aFl4VykKBnqFdUlTf8IVzxywzqzsizXEG3/AFCCjq+U
vk1ZR6MRB+2A/x6g10BgP5A+UDEO24rptZ9eANWXJtaJvHBYQQj0OMsUGqx85W+rI6beQnpXVZOw
ofZNc9HpYjSJBMAjuxCHCpzKRkkalBdA0iLWOmXyf6RYa+PlSJM7Cp8y/PnpmBsFJIpQRCi3EgrD
kgiahU6GivzP+48LfRhTbZARS4Omu9IknfOx+/Da9a7nxSIgKjvaRCKZy5rdgr182Wf5MlfdMaT7
XsS9Sn3LtNj38VjFOGVWB0oUHocCphNVA1C8M5D6+X1A7L5Fn9PfWagtM5T/wwMq+NG3s1A1PqJ3
8++k3iK4XzIAWPVihsRffPNyUqqwk20X5IGvGXOGthRQKLShdXb26CG3qzjS33Wop/aDVV4H+BR1
mTT3dnZg8/3bXXDdngHQSljvn/eiQZfeBLrfjJOIEoqL50Zfy1lj8V0K29iaaReDm+HD0fAL2Yxx
taiAdWmXe/TV7uDn6tOR4QvlK11lqyr7VmAabqD7JiQsGyrd2CrCXR74Fk62x5l47/ciO/EDorD1
S44ofcdVrYYl5mpEfOde3k+1snJhCTvI28AOuATjAR3z6u9/Sfja1YDHQCOR15qGmmwj33hKryaF
BjUN26g04Af1BePcSKoNh+izUrlvE0xhcehlnHr+ecroQiZ1zq7c48lagyan0Uc2Pn4WLzyqTkQv
opSJX99dPPlEowTbbLYEtZ4NOWQVm5cL+YA9qt9bclrFfK7jSRumR/gy2K/QNdVI5198qd8SUKr9
zg0rUzpQsyzI+s2msol2R2MjmT4wbn5FMnn+tFt/gABOS09FJ9d6EKgLspeCRLRb3izSFGUTi9t/
Ag+DJRjtDOjJ2BauN+ZhM2CmB881fJK0q/lMEhuYrPPO/ANkvfXj+Ue+WuBtEGdEJTMXU9pmdLOE
v0bEBhFem/71t/HREUzEWw84/QGNpVroN7HLhhNxfq3OXjnxmOcFtR6H026nf0jj2OCwFCWQQTui
Bah959y1CX611cDeaashZEkocdxLAYKZ41a8ZCSK/O6D8ZOPQmb7gOa2mpTYYW5jZg/rQ/cr7C2u
BqOpLDqaTjI5hXhx5ZKKqvrgChYLsae6yN9pcPoDCzOsV7trMveksA5AOQIqis3c8mOJ8g49aawg
QF7YsWACXg00t8af7MNxwzqRVYuR7htT0J8pOe0IYqXRawLOWi56gM4z9eUmcWjNqiRu8DdKeRAr
zM+EKV7eeJPQjtOUmavap8GYCyqZW2UvjxmB6ilmbsOmjH72sa9H8CkGCy+fMufWxdgjty6w+ymg
xcfeRIPUGnpIp6dbhMqgjlL3h3KeOcDstqxkIsR8PwThg7O2/j+LhjuJ3MBt1S7RWeO8GiUapi+K
ksnhVAuCkzDr8TADUMJAq5z+qgBlS3EKn+NbHA7OMzM4Co0fqoi09GG3nsc5tY1msPcUk/txoFbc
ZlrXvvb7mcLMbB8tYxUbrqcTxijkfLExUfrsndQ6pG/krc6RqkF0LPQDsNBeenXyS/cQxm9nuqZa
ZsShUrfxSEHtMMx9cxWLhu5gxBbyJCzPEvvPnhwkkywdjoeQWf9Oo8JRsw6IXHtmygngfV3ahaeZ
kkSMRA3Y3aKv0v4leUczd2Scl4qoA9bS353OQ0WY7RGh3NH7PYODq1NhtM6jDJfru5R82pra82hY
wj+5bs4C3oMxKO2jB8MhX8NCZculyCYhFBaswpCPYOj5C9SWHNriRcQvL/xxdwHHfQb/4vZMqBCK
vQahoN0QroKQjPHQngPAV3ogFvS8UUqE3PQoLjo2AtIHNQQ6Ic0/BmKt4rOeontrYelOBWeuxmZM
JgBPYOkommPhwe7EoxmjG+YzFuP8l2mncbTuDyozv5yKyleI0TizJdaHrAAgAX4idNumbsaEWiUV
rXivU7RSWQWHylt/4SUNYzrEC9xtQBrqsam5MdHC51mIEL6quLtQD9WQDEklGn9I2OA2ZDEAiMss
0H7svyDuWGwTWBopL4DHca4RrhQ3uYFXUQth4N7lGxGc0RTazN7mgPyvokC/quJ9ub6320NYukJ2
2xTsd3HB6MDvXZ3VfVKv9mAILzV7qKpgsc5iYT2uTTo0UpUPK99caYCPgz4kQ9OcUmMtlpPvg5+5
IrU0DTu2DKYeGXQwfj0cABVZIF/xaUwQ8GghsSDplVw69DYpYHibAYfG9VM2QNpe7elt8eZ3phum
GFcZq9mdOXYP3GdZ8av0YEq7wwAK2TW5aqVx0eEfHo1lJVjShr/MoBHXzyGoR8l7OXq0dARZ4J7h
Aa9ggfss+gxMHVyLI8aoo+14y/ayMg9EGb61zCmX9dkun2PYhWJU0TnULlyI4qRIVzRHzizba7En
mz/YAMEPQ9ZS8pU9D+Qg77xx3LxPxArK6VRBbxdbWoFlmIzHhKQBYEUlWa9PhSWG13VwCwqr5dZ1
iHRaTaUAlft19Lz1tx/CLyEzb4Gn/z7qdXMNjelNzstTEhCUrV6Z1QD2oyHf3xoKOVkyDS34Tkc1
M3w5mZqv6j8rKAdooXorm8FIns7TWLaAPzyJdzg8kBpYtqMax8Roih4MuG/1+6OTugkoJn8T89Kd
kWm22vFq0tiGoMqr1XYEwDJUiB8MpZlTfXtGDVISkFuK+0z5GFP8ykVL0izahqhsA8XYeiEA4igh
bQqi6igJ3y+OGO5ym9c9CJBeaOLMYjoYDdTdAQfvadz5f2DlbuEI5MjEi93cD6AMmp7R0tEElu01
p9tJ00WgOrUb4rWuHTVzOZvHRBAR6SR0S5Df+FMv+HPF8gDbTm44C56jr1SATMEjSo3vAaUDxHX1
r2VpImTXj7boMAGQ1DQW0sbdEOq4kFJL5okMFm790+lbFgcU9otP+NzRJ0L4N2f8hdmiwkWDkg1u
DLAjOrak+CU3yijhWBWNqA5HLr7tQKgZlObW1UgaFFnAOnZ+OiXAsjD/UUw5AxGoOQ9zq/JoSg0V
H3H/dH7i/ysm7v9lrcl1jrcYcxyk4JkEVYAMIzJkb9BfzlQj7srYxmc/J+d71xJZ4NzeE79lHNIM
MfahHpijGQfnsU9JP35K1jGheU6m1n7CrjmhdRRubQOzspwtXZtAwkcnoYLnZZqt0AwLrXfXc55y
k5+9Of3s+i6tx/YKOt4ZTcyRQ2umghXcmzbp+oFfDnxyGLBBmLFUOjQotZjbfqFFgwrm28iU9yyZ
wALsrvZdHlj5/+m+qgBS0bQdIfvrcDIM8oj494FglbzH2bEMnkX6Bi/rdHJJAbXHMpum7VNsiS5D
2MgXMOIF0re8ayWJmkMvyUqJdsAXbkzJdmHxfwRUpet8tx5Jn/4DzdlAMDjh8/qYVu3TTl+mAKNk
vFTNqHnY83tQkNUhLgiSkp+GO8BdST1cPOI0IHkem/wLLvg8du3Y/FmNUZUAMSOq53/Ajz8uQjIv
joG9xunCa51akAoM6AmN0SNplSQx7Hz2L/dAqjM+CQFjhJv1yuVmiAxSDpLILcFVoNO30VFf2i4a
1nMnBjYW+DK1MCllYWJ7J0HLtOs1oaA3qhJk1jYFpC/kw+qZ/CXGHc4rQPc5PJ7Fh3kq5Sqs5HSv
B4lvesP7kfcD2kxYSaZj0JmGR9Qrjej+ilMZJxCAWvTV7dMGZZHZkWWIbEhY8QmtzzpWuVIUjNSc
eioHbeYPAE41B9EdgpgYbV+ybCI4EJp8dYRqV3gJt6qAmc5vlZCBc9ptMvh6Iz49y/IcKbUDIO+T
p7cPm+2pJgBXf2VHqFJ4KkVk9gljlxWJQmYMOwJtExAIkGmJD9nPmFPmzsTPXTDKwBrxtDjBuQWS
GFLkADTb9MYWo4dwj9M1/Hr3W0C6fWNpPmxFnS/d/rfhkUtLzLU/r/S5g22A9zH+UVX7BaxLSyDE
WkQvd+aR7hRkc5G4h68/gGoj6bhGNn4/7enXYahR11GQsiL80iYSfQnOehArCEdm2KdAqCLv3aVW
wfNOoUmkJYjjDBXlAuGl943FO+dVroqb+sUJ/zCtEyktnRqXJjU1EHihxClCtW0Y6G9L8W7WQE/l
D4GlVScGl6TxZ6bspWutNWxFx4dUohMsWz4xpuPzaR/ryV2b0CTcel6az9RxCUGb2spUwcxO+Cwa
0dIejvgmemu/KUZSWISacoh2ms7ef8N/NRy0aSKdU23lgOhtKBYqbDK2jCgpeo1lTz+f2dbCh6kt
2eUqNxEQK4/wgArSmv9CpL+zbBAnLIxZIIwoR2WFjL3d5A1OarfYdNb0sqehtlRtzYWPQnBD24eG
1zZzsQss+Cy+1FMyzcoja+B9/RdgT2Sbq56h3xuTXEf1NNWACdgCy7+aaVgZ6edSQGXqU4fADOZN
ASSRI0NxV+K3TUDb+6kTvSwDpdk3we68PfZyPLjZq7M3NIgg5Tp4gUt/j4aq/BKqqk8M3QjBY86m
SDe/0EHT7b5JYFs9uXDXy7rzZZXvRYkwY1npU9/Tn2di8CcJiwKaVnzfEVM2RrWRjku6s4y9EHV0
5dC5/ZJLzoLSvEkqtxmJQvo/l+vARr+uOULS4oDsuNU1fEN56OoOoxRp0+fhrvJ5Wke0iiyTN7bm
Y+GBC9TmDA4Q733sLGX4kRa8skkUrnix+edLvriV+N8eh7SsYPYUFJIIYAbde6GNFUTpJN0PmMOA
8tVapPIKBW23hXqLOST0RfBfAb0U06PlaMyCtFIhJOHqadFWGA6Z1cUIcGzHNt/tGGfU5DTAS/gP
qHEH0JpU3u2pNBuHSXG14X6XLUti+SL79zCZHpK9qkfAcOdWblbhrEgMjr9PAYrCwlhw068NaokN
xvaNg+oiXoD9UHbgAV+uzD/rcxwRCotZL9wfT6fYknW7kqtvZPy27tgXpK3C1Z7mjzbV2ncdPGRB
pL6DtJ4HTWWSvoAJ0X5217i2TiBFHs9xTpb7yP3ZvH10vzay2T/y6+C2KKetd9b7kaP5OpOLVuaS
WltBuZ9hXlnANw+XZzT0JO0IAbwIUz0BkZ0JQ4e4211g7fuLXddXic9LZ1jTorKfBUHym8cJCMG2
NipYFMWJb/vPFMPE52TY/lwBn8WJYD8+CuyVsFRCxRAWO2/kkR546n6GT6Z67N4pSqgvCBjCS5q8
iiNMSgf2thczuoW6m8B6ZYNqKeYwj4KGEMhSbrSkRrPelI4mlboIaTyoCBZ8CcrSqbLJe8Shm5Cs
aCOkVnLxTrEiKrzpMZR+yDANRK3tSKUave+ad9HAimjjKb5ucuU71YBZgXpqy4dF8xWHgDPqr6xV
XZw3vo76ziImQ5sSXVMAxaEYc/LNAVRE6lbSZcr26lVv1mXXbDbEzj0BFxiq/vaSdkWQ+lrQRUKH
PZdGzSZ3u67T1q5MczxnZVDIJKrXeoD1wr3s+S0wQBw7S3H7ghNWjJT7qufIE4Z5t7NpIkuGEznR
y+4BgYm4aiZnCukFNZHG9Br/TkZ14F13k7OAbv+zZKccSPCK9zz1T1kn88oEQ9yshrqJWqu7X6Sc
qx25VouuMqa1VUGOSJTa0r8FJzNOgdyzL4i5MJ1uI38Y00fy6tx3XmVqqpYp8wXF44vFPnAYkH/t
hiNYQNS6twALsJlp4WKK48NKtKB3old4Yz8q27xSwNzin2UUjVe9oSQ35uQK3jM52oNWS4pfWblb
/aoEJNQD22ZE2w5v4fADe2L4z6XWBaAKtbWYspeuKs9acXGNDx2z24G41Zr4Vfh2+FJtzWhFlMgz
yL+quWwekK+c3iV6s5f+nyZpdZgRCmTCEGZghzgCHhjZmPeCLWfkGb29ywRORalqq1oOG80mEif5
kid2pBY74AAarNfGRNYaGClc890/CDwbOIAOUnfgXs7Z3lO+GBgXfTr+jkwt/uVv+rzYdiBUpzC2
qFRGNksGjr54HhanXnPC7Ttx9kqT1NbQn6fPBPgVxyjk+PI9+FueHzC9aWZBFOTTR3BemDfEvhPt
osSREY9aYwDkzvCa6HiHpqVKVpEiIDZO89iu0JfrAlXKx9SXblWNpt+8P20UJm/GpML7d5+tqAs6
dzqtGDxlFgshtgpfg/nNa/HtG5h210mUO1/FueDREGM6B3xffdIPZ+XIdqH9K2yqs6jX6FCKDTmh
00bR1NwwI3dGCqwqrLVmEuVaDQepAOcu4dXuPRglPM1r8YsP5kgiDjlIL24zA15jLSCzkIcJODMk
ng8y8bN/bFhUlRl9fY1p7Uimlr96WYCYyxgfY/DlDASIB7KujiP1MQ8eyOc16DWK0ITmVwHbpNsL
MwfQVByLtB9wrvasHxOyjGuYQOAt43V/VaXRp9kHLiuYDr4f33qXv1qluQRgN87qASI1R3HXTCYT
NAOoCPNqYLSsUv3VOAoWQQX1hCEaw5gjRXuVPZA2v6oQw0FNFON/gVjXGXkbjGG9y/BuGKUvdMtn
Kh9RrOlVCscincQXhsXR6dW585VdTStyX0l3YakePw75T3BwCemK3CthOgv5Y8SfBO4mNFLBgbyD
2bmmZGx6VAsAnLuuWV9S9TWmejrXdbsKEW8047cmrb9Ajal1BRstgG8RdeKpGEiTYjwd/HmQTM/R
ag7Fvsw6YGcpMxlobl5lkryx3BI7Zg3LEpuE9ZpsNsI+T9skXnkKQj91n5GxEdy5JX6UVORD2/lP
RbHbh3Zc7GrLen/P+aXVoHF6u7Ia3osoxOAwQg0YBv3mropoezGy3m/+M55DXDy/+jHhS9NfRojF
iMg4RVNBzwZfZb70Chxjz78XSuQoWvcCeqnOalUNFuAltbnAMdWXrmSXwvBySQHBq2MQ12Poe9xe
hk4L+nk3OK2qvYeVOWvCSmn1VoSWSEW6efOyTBElD1HlQmqm7F70PGB1LcjVeahHJM1C92b2FY50
6p4kqjxLkj+0e3QAvibbc+cRus4gciC99myoe3FS54t8s8a+p1NwneJPlTa2QrWAZRShrePxU1Hk
YViyqshd6iv2BrBG8Huddfm/cjdkv1tOEYYEqNGKs/9yCtl9UYp6H8eu5OH9MtDeGfu/Snrrms00
SREW9p3A5uxrXcMqwqNUaMADYeBn8YYafMcC14GnsCsh8Uyz+4ppFJWnnc/91HjZHuTJhKuvvA2Z
hIyRuQGnQ5EW18HSjeDr47qPSvHb8Vw6gH1bFDVyMvJVyZkbQg0+wg3dBaa8YAZdfZqGKADsk3DP
Q9+UXqjyGrcL8+B69PCY+4t5Fx1OvpF2l+rnNgy9LS0eNM/H27+O3CSV3dHBh868QU92VihGFYJd
tgy0yHn9GAfhqfEa51VIGyp9gD+kZt3gNcB0aIWqIS/KuVo2PmDlCHe0XEUbEs+DD5T/6kYceP0k
7gGVUxNq6e4dhybS9jV14sgmGTpYHSQlHbS27O8UWdxMJuGbFUNpt694Y7xeDUFRlI6OrT0WcgyO
0aoEAAN5Ebq4rzXVXyiXtVvKyQ3PwbXbhXoRmd8dDSXovxZoywhcP9oN6IA8dd7Y/xUrWzzbEw8x
9iES3PBpvsc/WZApd6ZTT4YBZfqeKX6gK7H1Q2cU9+81AQgNuPIsGnBwsPQbX67qugSwX56f6Dvd
TziCnWx632AR/w8g53pbgc9i8ugG1YRTPaxAoszJ/uvd6S0ZbIJ/4bTQ57PYEG1Mlw8sgFEWVnuJ
QSHD7w9+2TC4JmpqmOsW0avZ7rbyH2LmMYcDJCrdPUH+cLrFxG11s+KU85EuRZzumLrpw0WCbFuk
g0dpmCWLd63EIqCUVZB8bCvgVmJ2j5qv3rqDGd7qCAOTiLblOPENPFbDU+KqDj6djSVJNbZ0Bkh0
uuPo9yMphkcY2QBH9vHGAYrY3M8q1OtiJHStQr+C/qmnKLB0lK9ciG5cMsiT66OIJKXTCju4vjpo
iefJ5lq4FoWqsixLSeqbPSDGZFoGeRntUZNWmRoayWkLrX33AItK5ax9e+6r5O5ReF9i9njz1lhv
NodM7rnpYMSg4YZu+CWTjcRmKtZ2BqEh4HpXDrvsUwnS85m7mj4W5SsCUY+nbR+0xWA7Md6aKqkx
EJg3GTbndo63miTjfBMRIkeZ6V/Z3eiJ1HXvMcoFhk8GuGa7rBTQCCPm5/IvB4BVzJz7pZN5+RYP
zBUR491W+XZzpXD+4GWBM0yaEO29HBJSQIPPlVPHjXCc3XN9N0Auh3Q54lweIswFRHXYrMaN6B1/
bQimevaA4mOpsCpqn93AVQrOEW5yW+hvhD6ZJLieRyq3cQZEosuAqmYyDJ2T9Jd3W1hYu/716TKp
4EE4suz32fscCvk6sDjZ+DwfehEMHZopsIgvWfsoQwJMEcAcsZrBX0JyAi66cT3j9IjqY58jpJ6z
NM/8uRo8I+AGkI0a2dA/wboYKFLH5Cdvyo0HqF5cHEYXoKOtAn3QOaUNW0fwB6/bf0jZ9+PCf1zd
EGaCjQUAvAyOfP2OuUUkk9+7OoT0G/V1913yc8POf3VGDUFdzk+YVzPE73iYC4GzIiwNhwoZbs6E
nEZGbG+c0vEJ94NKdK0zHraBVcFUo3Ypmuf8moIrydvk2gdH6OXOViphRyx1NLA7xEQ/gQbgqvuk
wqKddA3gfwwFlJU8VPTNp5sGtUTELsQAtxQj7TVhqCa7LKxstLse6HPwYAtTPDv6jtyMgCaLOd9L
+OES3+oPh2JE/i9lSpt1R54IvUVKzmueww7WbSecPuOwY8qeSH3EbhNd4OCPsHEuwE/DPJI3oJ/t
CIstDxB1RtcdS20PtuNjAvFdRfP1KkmILHkVN8/eLkbfrhEo6/zkWMtjWAtzMlHukQ0W69t0MVpr
blxtlm7UL2mPKNZ/Lc2CyR2x7kuN289qKZQ5YdQNe0qaIffPz0cSg+qg+ALYa1A9WtikZk3Za6vC
ffyVUCL2NLfkXZT09Exp1fZC1sqm44x/hfZK3kSYcb2cu+VKhzcnDbAgbvdE24CO6iDPoYXNfeX+
Py8fw9E4Rg3RqN0J0hx4BpB4jVX4o02L3+H3syPIh8N5FgFLigMj/UzgVPXE7TZdr9jKZ9Bfj6v0
NasoVzdTtLddmJmXEK6FXGZ1RIpWYHCXllHrHWqK5iOMUgR5aJmSyBu6UHgegaYd9JP6ov9rzafn
Ee2hNAIb4ni0OhJMNJMc0ZNbg3+gMo9dbZzaLKweWDoSwm/E6op4f1xpkEp454dj9iYN4argzVar
cDdfoah8ymcMCWz6dFX5+6du7Hqsv9AQ4tqGD98MF76nLUSHYPqlxFAAN5Bme+gcKk5BsDV9Saet
GJcWZ/C8PM0nHtcl1Yluksq9uhPnXw2EjKnqlm5PwibW1kSPPc4nytpucZLw6kXIuOq4AlopkY/S
nxbkyJrdCT3UN9GXySemMZAkAfMqnWZSPOVLNBOx3duzQF/Nj0oPGi30LLO78ygvKuVGbSkfLOKs
YfVdzposKmqs6/VDinhdGzpVKByLStYX5f+n+Cup8qpU5EKwMFJ0sB0G7yKj0rxmSTz9QvwqWeO7
77QfBlYKNT5kRIc3YPWMIbssAO0NJI3GrGu1ezjOhLHWMxz8mQCPOUfBuJEA5cF7FiN03+G1zLgg
93gBsj/9vK38DzBARr4bInyO0oQvxgzBl+7jZ9ipgvStpekCFZVU9fhm31zsbCpzRSL6xrP3NOnS
2wd2gHoY9l+VDKItkcbmKBIOKOUhl7gQqGbtykueXe0B9EK/p9z6szFHCUdbSn9LYdxjvBVprLkx
KA5UeYxxcDhjzIPsiiqXgH7H3LaICU2LtdaGwCTgwufeY2LpHw5Dl2lIWnMfjMiOdalUzN3ReCtJ
cmk8wbOXmODKe0tuIpwk19d/gjJqOT0buKoGTp1/fo9Thy9ggi9SK85aEnB2QLdJb6LefdG1QIkr
v9QGtB0fd2eTsMM4TNGU3Fd8HdRXItn2nARrEYBOn9gx6LiGVGQ+47IEmq7/aq2AxPMqNECZ2/Fe
ftmvXyW/jwrY17P3fuuSYYfkM4VO0WOcq7INxhVDVq1WYa7pgQiY53Z3aI8EWRAr/E/HSgDmZvEn
pQZBo72azfCFpY5rwxVQpOP3z41pCstJ1gFhgVHOct4jN5zejL207yGuurutfo4qjjieSLDO8RX8
Nzcz2dx2cu8f6OMoByHivvAHHac03A3T4+/KBxk5DU3U6oV2nM9QyOZedCdajrIyCai/JQ0G1N3J
BCU866IoyEYSX1+DezMPe4VBNXqdK0hFUfbqWYZczfsqGUajhlBuCcG9mQaPt5UuYMsE13/j+vaj
UB0gtwocRdNv95ZB8NUBvuG8LJh92c2UZquPZmx+RIXF17axzCLJvZr+GOv+vwchdVZgF0P3WcZ9
4kc7JXCtkVuZFtkGUK5P1YX9SD2fFiko7IikMX5YzmJmLDZ3bkYWWtlxEsupU7YPtUFjZUHFAzVh
cUI7CX8KZEBQeYOsv966/wlPbrF7cjszQG4qIDBtC3jYzV58Pf8DoPfw7pE0JouPFgDDfB/IZFK4
363IF42aCQZP6wm/aflxddDzn1yJpQwah6luQFBk2RpGHKWWt/Zj7J4UE1pdeuK5hBJFt8es6GeD
0uxyhktk5z7dl7Ek1M1HPz7hkJHGj5QiIJ7G572rG3SCIQj3lIzDNJb5o+o9NZH5fm88eV1jo2sM
wPRENjuaFjS/OvHR5/OhaH+4QTjL2S5W54NHdvmQRmHNMfj88RebKZruqXOqimyn3/gJs8MIhjje
JidRoSSbjeUpbcEt0LgxYM9Xr5ldn9P+JwxEJsrfGu32C6h4JjsIC3lcngAfJzCdCRnVCA7ICySA
r8RBpF7dStKP3j/6JN/CJUXfQuCnyoTmQlnPA+r1sgUUF+LwfshDAhJB0QjfN3w60I0CofkwreAr
xXPqRhl/OTRIBjfZga4sBkBtoM59NpB2335MrqUS0Nx2DwrwM+iT9rL0NxhxpsVg2HuLOihF+/0F
gqbPcTbBE6l5dkQGz1v8ShZHW8ALGu/dG8E92BxZLUVL0q+oFhNCiZHFvvW3xRGLBw9WRGbvM+X8
YXGwvpp+f/tWUg1wcfJsz2mcFmuCDq+eAyTSLsPgz+Fn9QtjGpYYnU76195DSr5f9kObmNa0SCCX
+xVZl1hVCcX5ik9W98avkxxLM6bOYGtnnkYjSIP2IQPYsRkTtCQN85FSLlvXf7EBtiUvjG0zI4OA
65msnW18UuWmw8baUNLibAWarJFKGHdqZsXJj3PVFU7xwSHGoGFOj27jt7YNDVlQh+aao5PdCshD
Ar/YYTSS68Yn0sNlkm9UWXhBv0ljZrE2a10vWzB7zDhX84xKr1RLn14+7VbS5PVZC0HoDXzOCgKU
+MOfs7GB3GMh06htka7hOb0O5AOVfqRYXDEVZ9zEpG1V69/A+UQ+MDiVn9Fn7q9lBA7GFwRnqLRu
aHUg88hAOJR9LEvMh3bB1nJCBlDqAJFAZum6jDlZDxRwaqRo7DnPU9Du7qXHojRuf+qMkoS6Zzz+
WiImjAt14DWJXa/MUK8iBTA3KQjpByVhGQwdkkiVubONo1okxqA8b5TxpMoLfs1XUvaXg1R9RzJF
HJvwvRD0o8s5na8zvIjr7rSODyIyl4M+OdPsnlLL8I7Y0Wik4WId11zFnlNiB4EqH6RiV6d/jo1t
0ieIDWpbmem/wj5NLJ2RQYktTY+fUWngG113J357ErdYLlgE+r8XmCJwFhnZsJuaPCfzUDw+bH+O
eSycWtE8EN7YG0H3rEJEL2uaYU45Tgjg1qgOFBaMU8xxQHW773Lhh5J0Jc6uL4MaNuRSKtkKIlQm
Fa/yx6fKwiUxx856q7D/hpMRVc+wmmDwWFfhPu2Ggdnnle0vusLMedN8nz6Ch35pezpFlqMsVI6t
FnDK+4SerFjaZT9nxJSWINuEZZ5QHQX8yCm96uj50YRDFoeVfv2hn44GM1Yr+Jpn14kH9k3ClRLV
zgOsUSbp/DEpZUgoYfvBqQCI7+Su5GbygER+Wd98yJqzxEdob7cSsCcJDCc7L9TnOPkCdu7p5YW+
Ejrx+/gqzv8x6RO1TC/KMOy9qRaIKEonlLKl2D0pUB66O7DIKuyXZ51cdcd4f10OqLJAmkX3mef/
yerBW0mwBjgxswkVlZt8fJO2aRqYSdK73FyM2V91zBCRI9xUSD58mmA+amM2lTQ1StYOwOzbB/JE
jwA6BGYS6ZsJ5LUnhpLoRg92yT7bnnwsYxC3QsW9S5mxkrxFEVpgELTdYIbOBTc2C08uQGGEPD6Q
rPhP3O23xXyG85RpuhF6DLUb7eSjFJRXM/xwN45dzjN78/IB5KPmfTVwA/WrY+YR0s2ZzhPMWpgZ
ABwrCb37wFZDESuE7DuZobBGOn7o57cTYzx5iXobryMSJfTnyMMjTvC6sS0eJaGH3CeAmlxrD90F
OYNz2pEjV1OeL0j2gz257a4QC3XWQT38tpgJ0dx63kIiJG2hrx1DJAw9YV/00xB5Iseuzmy9MhDF
JpyY87edGlW0/rxIruJWI+fAdfAf4HsXy9cIGszEFxh4QaGQXkzCSl72TTeJQ0uKMTdCLh/qlWGE
sAHGl893BTq7bx55+TrzixBOv9Di4jsTU5emebb00xwTvr0m6p3x2n+WU3ZYEu8Qm8yAbBSrdmhj
L7PyDZeTJ9rTYlGBM51iz2MrY7LGJX0W96bihzF2tAF3WfgaFB5VnajtXk3DrGNGZIKDQPi4qNwu
sBqYzBcyHtWsXczxrmrgrpjI1yYJIN0AAXTGluNC8KItnMqyLnpLVHs1BGXNrg3GD34ewTSUN8Lc
mkN/JUAwmGleYNVGYJLUhr9ouNYIxq+nh1M8qqQgYW8ZBUItFbFHQ8vSs08Ru2N4rsd4NB35knjq
/v7eOG0jKNNkufARW24VlTJNZw/oLxDHOxfZnIx6eJsb+ogBdBpT5rH0NpBzhHhT3TgtqrBUqd2M
Za8PqZ3aHX2Itr9eKBZGvx8zMIwIHIXN6h6z6kdK5JHLyRPZ/BO4WIR7ui4TBf02THwpr56OnyTx
4GB790atCGn/sFZV7xiDEwGHvA3PTfdCY4eEmQdXQH+wkBApIr/Ic2h9vYalyljEYAYeNVKyT+mm
HRZgRVtXJ/72xC/qe8+QPEkuqrAOKPJyQ3Ih7mBBkaGWOUwG4b2AH+FFRiZuDr0ggrndf39DLK30
Uy3iJ4v+OenNa6jEgNxj6VTNcVMHd72lgNWUiCAi9sJxdLzhxf8klUH5BSZUUy0lMpWDgWVB3yk3
S1M8Of/+AtNZX/bzn1yyJy5bjHoQA+LcGkxo6bwl7aX8deklEvBTaV9LksjYUJudn654CMid6M5T
7naTxVkzHpIf7LQaOeaDcLLeIt/8DLzsxr0H2hlmZraYiGTgJaIg2mzE+UGz+SU0SqEX6VFvnm8J
KxToVyWhdqEsh+X/AkdFDyVsUP0PmP2aRCaHKEectB+1dtQeeqhBR/mgzHQ0N0LL3bpCgidGFfYz
9HXoZeh//OKIC7YrwmGPbJbc+4ozrn3KjH2fW+RQCD/AGeQe4UCUE8S6DUGGj+2tGIpTRICc0ZqM
/5/L2rm0eIVk3o2l/xTMdA1mJHD5gdLrkqFtbyYKGT+RL8qU4xVKwI2pyypleydO7LMjyFNFWZUo
N+toNqcHwsJ+ihFNHPlNLWSv1zn1kjVViYrZMdsNekUagUy2sEQoL0izJVZBQLfcR3w1wNhCJcEf
WvdtrNgXr3A/VXzvXyneqV3PKkiZfQwfiZvhX3eQDB0DG11gI1XQYJ7s4MIzMKWrjEv270mZl5bX
KXx0uP93N15UyjRxUClkPQvmy5RV7B+1rZEdP3pi24sgQvcKM1rzFH60uNXoLMj17l2K4swetH5f
GaELqOeAXL3n/PMb0WMgIJjPA5gGrfJYkeXFDLzlFsMh8/GUV4wAF/Nbl8jzHg/AQu0QuKALK1dk
Wou4NoLPYHS3me6OTu5NvfgMzgDkwpiCCaxcGpyr7hcKeqkRd1x+ro7fPfgEy3g/bOINkFmggfpi
UOA5rdHZcrg0QI8MbeX0uhKSRlcM7FnQY6jdvWrqiRjUvPiIMSsiimdw3Le+aoMU7Zga7TVpo2Kf
hRJP1qnho2CQSV7SWW++Dq3CE7f8rMiclhVh3XHz/3lZoFOk6lqcJk36vspYG3YOZAhHLA+NOzi0
Shq8pechz2T2A27UD/iVZL9OGCZjG2jULayeXPZaiDleg2iq4ECNSeCV9VUxr2rh7JZLXY7CIeUz
PDJwJuPHzIbnJqANSA1odPWcYlOyrjZpxMje8dbnOzGN0vsAw8Hnv0GiZGsw4oHx47BzWfnFV+oQ
1HYQpq/Tg5gx5t8qd3HmqGwwwlMrKw6gnHN5WD0/I7wmV4TqJ4Pb7o0Vm1ZWODSCziUxT84JQoFT
3+WaEfcpqF15dRdOuE8dSwJ36IdLp6IKZv5KtbpXA9pZqKxX2aLqTW+yvGiPchqpUy+ijRoe1CL0
MzI96ACCbLc8lA+cGBlMCmYNIeNZXAld/iA0lk26mIFM4mNXE+5qRZIEtVpBqQOuVGuclBymtzG1
isQwP37q/BvFSDYiVNj9uKzkvOK9bIJ4IwF9AZ/h4m6mQJ836/I5Djc5Wy+aakHHvTyUmZ1sPNvm
BvdSRSAhYXoKaaJnKiac2yry+yHNcXgkhQHqjw0NUEDqYkBcuCKldAFVQPCZrpo5RvpGfvon5Tak
DC66QP5IAT9bZcRFRWjOqe5YydJR/ZfDS8g4s+8HBSHRw1HTr1uSla6/00a8lWnVFYOlzncA1jo0
EM+VzpZ3x5Of1vcZJC8fWpQIGR6qOuGD3/O8CXjY7CasI7y4cYCjAW9zcPANaajQ2e9cW4V6YzLW
mV34PE4yUk+E5yUfSbYmwSz8BBm0W7kaydoecskK0qEea1qAHLpjMyX3+nQSVZenvzhLF41SJqgj
txT+NETO00KVzzmINucKwBAx6peXbKlykal9KEw1r6dxCezM/b9noNWJ7syynou93YCSySphU3qM
eFZSjB+PLLXSuJnE1nkBF4XuxUBPJy79LNPwL4+qIhJql8BHa7j4vS35QBJg1uU9TYHUIqhqwL0O
1IIUzmq4Ho2o7wGcRRyCMv7y/Ldsa8zwmRP0ptEM91xSuZozm0HFKbtUkrNQ5zfQDeDjfSax02H0
60pk4GuYG2MiIY7QzfqTyb6CUH2+A6jNbQdMbYzz4BprUO2DWwMKgi/9797xz3kGyiBjp1tLXgXY
4BG+Jq+jbVCMpAIcailyAoXagV8JqIawbxmW5nYPGH5b0sGqpMXBpCJHm7f7+GV4jZQgBobt5tsL
EzgvFUdstiDCJV7HYZMNHMgAbX+HTV0aS6ULZaqtCKCAwhMtnTobJb2AYIcAgUeixN4/QFAIwIUj
FHrucF8TVMTGUbBS50qfta0ApOwgUjaYvpqJkhG4qCXEAAGiO1TLZL/53k0SVu/b25tQsTjUxEr3
9Nb24azactQIgeNv2CtsML1J9QSoBMgnE7Po5MIUBLbvfCHqYSyduTc8+P1AKzDi8wmqmIz+IxKJ
XlZDqretIBqCUMNtYW12SPk36C6bB/m82VpBTpUHxPs5T5DRdFu7mKAMuhZ+U58kLVqTGm7TTIHn
zauqK6RkbPOaBMT6X3NtiELTDWugSdlRsW0dXtY24dG+mgzckdLZUHHli3gVBEdTnhgTDg3l/ot4
0sxCvmSyZMOhcSPV3OB22yKct5NkpQ4pR54THXtuKDaWS2xuD0x8Z9soRoJliEi0SMi92QmCdwOX
yHanZmpr/Tg13KvvMbOC4nD74eWoRl2a5Kkk7g5pWR60gLgvCGAdCk/6iZP2er2XZ1UoiVhkM5I7
UyMd9j4jWFYaFuZacY8cLxAE8a6f1W9VZpoI7eEZP9jJLIV5hA+gkQt2lxoOfGRTO6Ur1HEvqxiM
sZ8jyAUmAdTb3CKrxbsNjRZ9jq0tshpX/7/2YQrwb3LJ01ET74CqFRK5RVJcN663WnEqtfNUWY6n
bFURii7ASA3zNg/Hb3RZ0UjQkO/71+Dn8QtU/HoaOgbwqGLBh5QFOu7hZfZgFGdcJziYuzZyaikP
o6usf47IRYPEQyZE2vjjo3q+rVyuLM6UfwEHJCNm20i6Xpyza+I1t2pySkUGeNBPd78eNX+G5ZKu
36KmeTDd+rBjKsqqMZ3TJDHJRupBOgHhfxBjQ1nP9DmTKHHY/55NiS0koQzNXdTnABa3qYarS+2v
9SGGdpcDVygi3S/O04esiMkEH9PSODXiVL3L1p0zDUsny7MTEmMDDc9dND6M2sjq0j2qSmkkWCmK
WziGTvBsaH0p1fBVqBJIhLHh9HY+kXJcj0BkSfHeo/y0na9yeNleTMLlOWc/xt7s6S75ib8HRe95
zSY+5Qy7k/cCexhs28Ns3g8oaE8q+/S26U8nwwm9pvVnt5oF52rvMHdomtmmN5N0t0mVu6vTaYmA
nutnujox2M6M8jZ3mQ/wLic5vvI+3oC6oAWnaGLb5Y7xbGSNtKxseM/hCieAWlaQ2Ijg3GGf0fXC
8a8mpvEW57pk1ZOeKagLdZ1LD44w+KT/YdKjnao59quh84dD6JgfmkuaYV0hmWgJtS3a05NTsdl0
1uLfwswPjBooVBaSVggJl8RtEji93+vqP+lyCCncBStf8zxr5lbsbq1XRI2mZFUiNLhp8q/rtLXv
avSUeGa99So5rJabPVqCqSFdEVaBk6IxxXAYLwgpjWE7cRp2qNtRRJeiXI8/iql/Nl4o+tyyM/8v
l+pC/NmBXzJ7JRRkRIifM2koTmC5gSOCRHyNsNDKjckURMLb/jBemmcsT7H1/Wanh9FiwYJ4eNIr
fS7KgbvC7eqg5IC8VcR2gOdvJwKI6n+cE6UA/Po/Slxf38XTG+ci55NdeAZS/gT7ZQxlyYFdjBPx
2rUkNycM+/v9tWWqgtAHfh/SdFVoiBkmy7ErUppcNqVuVD9PovHJVQ7arKM3C5stRDRvZnJJ1w1V
vJqgRXuwOJKOeINHTGmlYswO+e9CNazaMln4zIgfgAuUff8Ksey3682T27ZM4fbr7cpjrB4yln7k
Kbuih13Y9W3nCxi54HbPvh8EH2z2gp4kiQ0yvQAoBx7pQkv3tPWIU7xjV5kIgqIPBBEJxj3LrNwP
3CnqCll0+ukU4BXxIcBlkKowzxjSOX0vDIpjXqulPXvObuaMCexadPRVm01TBtQi7+4BBUnHGRcP
+9F8XMvBwBTflDdDQMa7inuKz1rFQjvV77/MuDvgEdoNSLmdIehzCJci/ync1tZ314VdKIwK1qcs
NFdZxPSyt+g10C7es8FvT26f7R4pgRZZppGhzS0wwFJNSgbXRHF6tta853v4qAbT9A11BPEOkSOK
noMZo3iMTEZPOImeyCu6jDNL4kMTL0P8e9N++NfSUcOZhaq9eiNPS2Rb7Za/DFU8ahjsv4GQV/L/
hn+tKkl9eNk/Cdeb1AgywOfObWdsh44ufmpPsurzLTmwg3j+BFYv+iEtD4jF3giDSwrQVI7041cM
CWa3jdDBgBuTauk9IhPbGeUgjfXYDloGdZFopOjLkdVWSgXxxJ8egKZuqRfe1AxXVtb1TSSVvR2R
3sR/prYuYhP9DQbBlAkSFYboQpTNHtLiiPKOjizLLytCDM0fsyFkCN3ILoxKaCMRT0pQV3FI+aNV
lBGNhaK6gFV53e7mJPGx2s7pyb6Sblc6TPwLKMXaydZLq1UmcBmsP8xeIdbRvWUCsJQsMfCV6p1G
6mh+tnt/3869p1SRFlER9HA0OgAlZ6zWiMFwh3Sm8uY0/hRmZhMDR983ox2H1FzTe6ejArauRuyF
Qa53a0UG3HX44sqhXQ6+N6Kiv2M4ItzENjAqT+FBROZiY8xsMtjAxVCuzwdrSzR0mbcCN+CpWF/Q
50hZrcfDHOO/ID8aKKfQpYZDw03LVxsOLgKEb6pooBD9X6IsxP6W7k2EGiMNdnQb5GBBn6H7TIRz
SkdLCEfD6l5ctnlyu+6DTVyBISnRUgcGpAaVJ+PGEhbFj3B11viCPqQu+iuB91yWEs6UbiYYwu4E
ZYEv6OyoIJ1WmDqVEzSnrNyiAz6RNHLQENXDQKLGVWGHI+DhmOBDmwHcGcx8+hUUt0LEzGG2NXlM
HbQoobFLFe2hqVDqEvAVn7NIJztOfNsSszBwR9l1eyU4QPOx/D9uCh/U6rfVFexXo6EJ6ygAk7Rl
yqDb1xrbaQObN8EQZnZCFknRY5+Z7nBfVdLuvirWZ1ZBEObZm1HxDS6Qfq5alJ7fcT1q0CNX7kNh
DKqd2Vys9+vHR1C2c/RIEMBFYi85o2ycTIzQwIVocTx7MDzYbMu0y/23YU1JrwljWyW2k3sJXvC3
jaZHYfDOZAmanee+FEAfO9klpFCz9aU/1KTyHAy2vWH1XUiYI1qvD4AM6c0OBh3Z9Qm6BNgju3kL
4QPDab6KsXkWahwG7xUn33T4PjOl1itTskX1PmHX2h99aPWwIYsk5ICh8q4ZNKM093a5gNOFhpar
Jm3YZpo22s6YLSAAc+m/55yq79fa7TAnxRsXI+QzQUNGgCtGPT1UtmvCMJqqKcW3M6HcO83GmJ00
wqXU/jya+FngnARmXlZPA3bErO1y34eK59gNwxeeSuUgEZ4TtinS5bpz0O5hpHgTikuhj0ebhvn3
/Eaj/e1lejK27YAO+OzpGaH0YAuJmKZ9HjA9kGu1nG8CphblBve8Xyx9AB1GDQ1PwMaMsaIhOgXd
TPhkZkDlW4vRODMa9NpTnORR63D8hFVDIZf73OwsDOLL3tWEfX7aIihI5MOPAWXtaQsKXkVEEdkb
NtEUvkS39mOuwPU99wdn+L1NPXo6JCCma6Os0M49Cg5aXRpLNEW79E5y7hSLg0ckYg++J/fzhhkv
mQbuCn/PAk6GXoPb6wJog9xjnoBjz4J17s3PltdcaW5oIENnSVKc4PhwANwm3qtkp1OI0sfZUqmd
OIc2jYq3uq50b2F3LxT1pdLgyPQitgW4NWJLjoPOXDT9uuLB0OSW0Y8upKs0pcp2S/V9GEosk+m7
B0UuTz4vGmauQq2OzyYLjRXe5KHVkCazdgG+CV6StDdCpTWJ0hIaIfZObjlApgv/zycN/EDFlzti
x82QpojHso6bZS2DyAhlT8buA39781wxHSJlmVsSeMcdsFeOn+yYmsDGHVpOpNLAy3MN4jdqqiJw
gwORkygW3dKXG/zhdd1c8EvaluFRoqkvU7XBhG4izs8im7kl1Oc6v+d6ONb/JQGJ/mUCKTbW1bNN
JkfejFtngmavnKgz7Lp43oHlx33EEYhJGulG85BEeELwV8dNEGRhMRZ411nnc2V4Q3pn9hc43Y4N
UkaozCHArwh2EbGqvBWznCBhjbtZtuYp+lj46KzGZXcuxGZUV0RmSrfAMtezZozl8NvZr8+gvQD7
966xxfklO/GbCJPsYjj+hxWcSaGle5vKkaeCLl0FyRk1BwTpvqKk1hEFvmM7YyhlHxSyTHGIDyiC
EGtLl+zLMOEi+w1IulSMr43JuLPRlYzsTW571a+H4n18ZYmW9Pi0FffTgMQelpx8aGEc0Z/0EfVr
iD6pPCOLgoR/qhDZaMw60UdlAGZhqpmhe5qkNVh17BfHC3Ee9Ge/odt6xdEc7NRtxuBYfSKXbU3U
tXHAU5IdbtxhSWmi/s9yf1RyUB5uPrC+x53ISgfVjdXCR01OCqWliV1Llg1hOhaeo01ugO0hOUyJ
OArtFc1SfefdCkl6GEF8d2iXVQjOj/Yt9za07gI0rPR2Zf9PgR2MsCFYm/M34m+rJbcBc3cp5oE5
DaksLb+8VegLvz2T24Lgu2zxp/vcTt9i55SSgE28cm7AzPfrzumd4ecqe/cNhfSDdYnCN58icIQO
ZqG6VrEw9cG7ZIQFyrP3Vbyi/dSFuvkpGBknwFAVnJQOmfPCoWfZCRrb+GqR8kuwkIbkG6yjT8C9
iEkBgxwzONBa08+lRBj6YNNxL2h8oHIbx9D1qpEYyE+yCFXpfqEHewMpYjyaj3aVNsvx51j6215G
3GoRqVYeGcjeQGFoXuVaRYV+tChBFDkcr50BF8yQg+ojuRelDwe7Sd2xl2YVew/QBYnYZEMmiUMd
I4P6VK80bMS3u4suuyLXpSVE/XQGHxco3wnxDvPhZeP1xXGBY5rOM3xVELGqBwbz06coyLEhFUTO
kPRkBHAIreiDl/2j5A8OKozxBmV2YKFtns4WITjtp2TlE02/WHtO4Gkvk2s4Kxuug6Scq3k0+6LJ
D3KgIKDS+6y9RHieK7W+OL8ADwgWR93Rva2A9ph7G/jCjOcHuFSjR3dbSifrSfVAfMlHo4MxvrFU
V86g0pDq8olPv0pvRidp2nCiz7omFHI3DORMZ7RVfB7coilINyrmBLrEyXG80NrSwuq5khNLSp4c
dejuNBv9VT9/deESWiUfFdQOd1j5uxs43nykTbXZkyjMEB5gTOAilO9eFQolbdd9neT88M5d2jWW
6Wuvd9NP/Z7m9FeJZjyYdQB5MBTaxuWifNT4+kfsKTYFzK9EGz+P1ROq2hljSqLyygoOIiJrvCfy
1PhARrO07jsMWsuE3xlHUCPel+SbU/Cv2ghuptyRdRKjzjN4LyVvjqytr/vSDIRuEIi0GtXI1ddE
onqhlM1jGKaLEIVSMqaKcD7eEdToq89/nzkpmGg7PkdaXG30Q9WbDntzVE8I4SW1s/Khgl5GDLjp
UvAbUFkkNKSFj+g2mLYQvgb32B4A/0ojzKzVmba5CgrGpsOSSyPPvTWzg8McxgOfTZv+mu3bFecD
EJC1QQPc1DRN+uWgvXEsquebTOM8n1Tj10/5RRhzPJzLJW/qanDAO0DQsj/amzexjMIH3lz414wW
EDkFYH2eTbMMHBiEl6zp1UuLNiT2VE7j8rOxKEDLP5vr/dZj64S01EKc6R0ADDEumzlucRpXr3+c
R5cyoC3P0L1MQciXVbiZ0Nh1ygukYJrNQ9tYJ3RK1TGe/Xf03PBp8ANBSmjoXeu2ytdgacgp1j11
PNoQRQQRZVlV7ruym/s0qcj8Al1x0M1jpju3fBcFCUysNRYamBMX+Nhdm3fNsgO5aDvfz+QCdpuz
ONzZZ8lQXDg0zpsVTgBapyu/3XyJ1xUXAQVhDT6cfi+NcO8ugsbpWWMks9lx1QiQ7wwDb/yXq30b
1XsRIXWoNSE6l7/Nle7hzgRXfw5aO6z0dohtg7LQK7UyZnVL3pCf9p4zugywSzbTMu+c+a3lIy5U
bq5xijkPW1KCl2YWIJxUfivZQ1M52xhgwsMoc1N1dOX4K42T68AMA6fw8lAMJI95sLBfkW+7FKU2
hx0dbuTv2qsmaM4R9dej4sSN7DRR0VWW53xGmFOn4cjq/y2GUSjzzLppckno0Ev+8VOJZ0sWIYxU
JkynR5TdUwST/27FbNyB2bmCFLqfFq5m88FvZ/g/YW0dttuy6VacWuBzQXZ5KU2u3//MVlE97+rv
vjfC3cth8bYA2aSoF3rwzxib4CSSnlKF7wyfb/ZBdNjC5ddiyDEt7d9tn9pQ45Pz0yB095yVLRzT
HjiwijhEkkbXmAPqIQzKbQbe3nBSVCoMoMvX1YADuNp/3TI5oCuYtzJGHpF9DWmJM5QuHf2A7vA2
8Y9fmMR60bjY6yHhkT25l7HE7WKBT4HHoj0wdRsvtHK8omUHl3ZMK8ND2n4CVPdt1prRTpZHA0tz
dcGFSgiEUW+20lwYayLRwc17K5kG2BY/NGuiHBcnaL8Xeuatmmdr/l1jFU+jGBkh7QKiKLIYzfwE
gEJTeGQTP8btNB9GW1/M0l0xTuBj7WJCkeVFI78G7kSln6dhmz7YSHfupzCdYEW6t7iBegumZqec
dZuw3Ptuhnh0dUeWWDmkGeY3E+6UuQsfTWVN3CMx+TA8EfygPBjD2qzfeiuFfXARW70weJOwvcFR
kd72pbqx4NlAXun5xhZAiuTC6Um8wk90BDGFVXXyr3eqvrXq0rb/kHi/gSYkl9EOIldweqmBGbN0
PwQKaz5PMBY46uccNf9k2z/fmS50BBDpqWtggEwBjZNf8WaQh2r1lwh8a5SiQ6eR6oYfq8TXsiin
y46dJ2huJUpiA23fX3pNu8tyyt9HQ4hSrZx+mzv9HsIydEHIr4lp9qVwr6cQ8m5ewzGLynEHlKTT
osJ6AxY+bW3PXbjApYx43F/S4fAWMWTa1CHVk5Q+PqYdH2Qu8iUzFJmwgFnxGRDIpkEzGeRVUQYw
zHYOn95m2NUMdlz7NF1VpumSsqYjOmWhBAlQD0RKpFQI/WPg72Fxk7fyIxn0DFWGUfJc4GhFZhOr
7S5cJPIz97ZCJ+flLTIHN7QL6ofdr7J6THTyMNmeniymIenTudg13+W+5I1XaYdeSmlWHr+zzrlN
VNm2IfVeZdIuxvaQL03u1B3lnqGt/NpYjmSsNqaiUNXCcaLHyfV/HKvbGrNO+eiwbus88cnzirLx
XA5XDz5vkVLb9/Np73/1bzX0wJilVuX5ZwbjI32DJSknGUI56nrMfU8oGssU6BZRdnH77pjits7r
m7/f486JOs3VfeltUlysoG2y9L8VGXDKXwvge/FZHiIWb068Gr3uqBl69UmN6XkhtEEJU6o0L8P9
BhQcNscQ0eg/qOXiYhoKKLhHIFIuoIHq7s73L75PV5abR4h1nQCiuFZ60o8CeW6pHzn518OLISd6
1BoZc15TBHDMoNw+/XD8ts1RDzTAT+4TJusVQtzuEg/PUWEeBmF9fEkKYeJfjqAOkC8uiHXr4EkH
/7DRMBwk8lesRpUtRMxauSS1iq5f/1d3LliJ4IKeCTwnjrzCY8DwPb9dTBaBqeqpoC/uW+gueJaz
DJThLhmBeBj6/q1urIXibF0DVw4SDCXODxhd1RArGi+uHgN+215wze5tBe2aplPDz2Av0naSWdTD
0vrNnXwQjXNTS2RJHD9hAk7Jo3+sxjyRE63XMr/6H/nrzUHyxavwYeVn/+ep9xczZFLCdeRV9wFj
z22fJHE5cU6P8DGzEbDz1AExAAnIYNpS7NTOmyB9TSccg9GSOa0bnOgQ3IppRFK/EO8BYgNwof/H
yCENVO8oExnNjJkbDhLNQY/Ls9UQqeSNisyl//Tc4906I5KCfSR/jXZ/A26Oo2JfJRHhVdeqbDFh
kJVftZfCjJgy6JDLwA7BBMQmaWgHJtRj8BS+gV2gZrmWkWbRBERZ7pwIDjpohEFZwQg/QlZEzGFo
EUHGST59zjX3mAeOHm2evb3HSiEzgNRDZz7Rv95P21kXMLmNEFdUQFLn8Yqzx/z7PeT4JyS+UlQG
S8TlOSh1FaiGrlA8c2wDNv8O8A8PY5GgksMBpeh/zLfAEuUGbB8gGGgdX3E4WQul3BuSq+ka5TP8
l2P8j1zMPgzW8FS7v2MVtWXIhTpMpyma0JNYVGSmFx4KwyWBDWUoSYTcJ4g0ckpvHQE+6V4B2o2b
RWzBjPIwNVyF2SjUo5zo9qSzhp4evBB1147a22YbdAnWHqow842qobhct0/uwiFBdY5xz+nyf0iw
Ffvt3GSmc/VVeSKXYVqm8Mc/bzZWs+n6RN+Kdf2DfOBfBBBQokzUbG73arZTLJMkHvl7TTLZqKxT
BhDpBQlpBLpewy2uj1BOTaSKv7PP4ooKi9R/1iBLbXB30VRGPWT/O+BLY29eHP7QBOsJsxwsRqYp
4Z1gtMFy/LPxNlnxSTyWFJi955Bf7sTvHBCJlYRN0kh5ByrtgQrnvEDOEtn52nNWKpFmEq0vJsG0
p6TpQUamNCeGS0EBWWUvq2/6Cs24ZM3MPy5/RgB2E5MRVxfK7/6PvM0VQHsGZO85gDSKJTvqngMg
ee0egGp9LKOh9yjnsyNApQ7eJfhnCqHuXoVwic5cU4XF2JJ/egTs35Hu6HmUKKUczaMKIm3O1Tno
iQ3Wnc/V0VxwI23G2TYNAdUsJZyKs5KpM78dqSzgtoJl0585KH4R5I0cehiiKQze741QgE/uAby5
drrhMg4Hhfz07jGf/SyG2zB94ihWwpWFE0GfJ4gqj5JT8bOpH3uEH+E8OM0kIiti3qcvcVf7t8QE
dMOXQrcmginJTzSij7Jy5B3xkj2M/FbzAej9Aw8qPWasEH2eQlL+2NyEx6hQm0EaJT9xGghHpl9f
EUwD7xooJy+mq6LlivpErNJrQ/sFgOHg/wqAVUMSZElUXgByfuojluY0BHMZOFLCQ/dYIeteEz2i
H/1vYZgS1zDm2F8W2Tvo3R0RmrBRslnphgb3YJD41Bd8W3Zc+ab7Dh7F36oENfWbs4RCKrjy4o+/
7p5nciLPy6S+7EP5lEEPfvb+J66ijP01RAiIZj7hj5xrTIFkuYRuORu+aZWlq0vfu3rDag++3lH/
ytKQhFBUnL7Rxh4wDBk2qhzqi2PvG9TzaGXa0pukqM9sBHahwwXnYNCBUAWf6baFUbHXNMwl/1CL
EHsERbrBlV8stUbdGUtvjRwWCfO4qXJTJ6h0l76/e9VFCYY8RqNtIjKkcbiICXNf0VxAqFn1UETg
c8KO+hv3J2h7zOdCzkD5vrEIhgtz7FkcgdIUnCxi3Tpu2+FHLOKQ9Iro+nUHBFtJ77GrvGIRxYsX
QwUQwfKE5csGlOp6njmXIjXc+5/ZzObqECmj/9KlvnBnkRilwwVvZ75TL6elBW3y6rVRnQLdmcVN
qCkjW/Vn7cotzLmcB3PemqjKPcqfwTQ/xMnVHiDxQQzLi7Zd+BpnG75Op1VVwycD27EfGmXeKDwi
RP1TadVSRBLfriUB+U3gIfknGMcMeqFHX3/+SClO370lwkHiwNgp/zA+t4MQy2RhR635cM8dGGB/
iCNXVoMewEfSpVqT2AIYmeIq5bAlV+fOCJsMnn+z/Af/PV+iuQCMf97mTupwXWF0PQMN5HrYTWD8
9ykuc15GpUdGxgYrDJW2t0t0RIOQWNBxR11z03Hj/1DcXMx+xp2yAQtNhNUi3lDp+94noguuPzDB
SGdxQgIZsmYxgjPqoU5yFq770qmPoUXzUmeCsoX2sVfHDiKCsBurbCCSJOOdky/9kUS6GgTO5onE
8Pdyuh+xS16/PsMYb+vrksBuavldkM7v/9L0v1AjlCCZ5314UozkQMdKu2qo3TtuyKGXBF+dYMZl
LiDefBkon0Q2wy0D8919fiVUzvszSFKF3R3EMJKq5CCmzV76RmSe5Gv28rw8BQw6JSxk62zshzO1
8eeoRP1NQIctXB13AxIjeUd7q6Muo6Ck9Y7SGDMEI5qRiSzP2uK5udq/yae6h/Fy0YkbkiaLQlMb
tvGJymYwrTZ4D4kp8K0/vdY5mMTbyTvjkuUkCtMrzE9hs7HP5qcbCKcU9fBCzLOtohUSus59WKdt
e+Q/CHsev4T+FRtP/0Dt/dTCALrvvUMPofjfCjFQHBWWXaY8ufQQ0Ue8bqxvYI4dJSKU22I1Lvra
+AzY3fnwQsMLQ8OOC6RkpAKOYml0V8UBTpWZFQXbPNQk+BnhRQ0SONH/i9N5oB6j7cvq5oirucTN
EgHto0l4M4HZQk4Cx1HfQ3eyIpqx5wIai3Tb/QmIm18+ucfzqA39LF45ap7PwFf2N3hbkripp6QZ
w5qa0nmQTkrXrvLJFy2JWa0xPHFJ00Yj/3LF0WCMqnOLP3UewEuimD8Iay1wajBRdrD2RWTpv+Ha
mEhoYpQ+g66vYnKr5npWb1EvbIiZXysbXoDQEi4BJ1axpU57AeSYLTT7NP6D5AKZ07n4TLVNFxP5
qAz7snqWTmo2Qk4bw3sFzfV0GFnskBa4Uzulu+yMP+UuIRA8zlFJGF/jKY+sh0+BLb0df12HD6dL
WCkfc7jqXnSYHtuXuyIri5PG/s/Hh5o4jMkeJgoiHztY5Yes/lF+hNL0+vVIYIxkjxnz28LgNEU8
xucvMJdHeBFWPHqDb+sjqTl4lBAjfAEit1onVFT0uAH24ieK3rhNPOJhD3fkDIaICH2lHwt0+GcD
DUd98klCcf2Itz4cdYL5nEetXuz/oj0/BKsAcNUvCYwUZ0mFHTCEwQiUA09fCeurEc2HZLWWq/RA
acOsfSmIqxQYAfSdLIBZrwvuhOlSPyGoZnXac6uqc61G1GokemYy/d7lxQAIrXSIqvAA28zp1aJs
qXfg0Jk1QsTbMU50DA0ia58rLB8Ti6iFtgnQMLprU5mmUjvL/jxUKiQvwm57kizXQNEV5OF0APWB
R5rGdBa6a/0KqPLW+i4YEMps9UijpJbOVMHKjSRA2eGDyMTM++rPQ7kqPdF79TCtErpq7He5AJJs
WhA2saXgPqP739lbbQce/wmYqJNfUuOhwaTEqpaK49wOsKxG/Fv72qhDXWgpsc5Yi4tkc1tT/Ise
WlggfQQf/PCMdvBSeN5F4m+gCne1EquAhdh5FQnz1OKMqXCNNRCIGH0gNyGcLKJrYL+H+d5jZBVy
1I+XFM/qKRZZvZ+MdTRhF2PLkiro+BMj7iXAV4Pay7mCl0ERZGsh3A9W1OscbK2xAoaOvzqEx5HB
O3uHgPpR9CURq64KWOXbZWFyiqfMp6A5t3DUy8Xx92HTyMNhX74Q9dzx2Uvw17Q+JzHVcECEzre9
IwtHf0hz30aUn4i2IKcP/IT1/rvDby5HOGTUQUOW/vUUwK/5fG55dcqF8Wv8kHulj7KZKA3dkawU
WZZfXpi11tb7zSS/h4aiH/DPesot1iDeON18fq7WDl6LcWKcFVMc0MVvCxA+DcoYiLHG4O75aqGD
hWPOhwEyo9pI6XxaRkcxVvHk9Ph6x/U9melJqA5p59TB0HZvvfjq6MUTa7q9WuCk+OPth5jeYXuF
V449zLSbRGpPBnpLIT56nbMUpFnTsgafNGumJbxpc+iF1HnOUnZFqGc/c+gNfl1CVlvP1X6oNwYL
iUbaaOPBvLCK+L70q1K+2b09Di3f3pBmGipd4mfWrSf8lgGdE3hB8w5MjPZISMgQfjVzXvQfmhSU
+G3d+Op1Jq7sbmQoV0SR1AKuaEwyr2TzLNiBUmWITCveWLl8D5tzracGi6Yqf8xdf+CurDcs4igC
8spyyGihwaOnuxtRw9IgCN5DN0+iqcc1R2bHhkvtxDP/9dEKP9ht5N6lpfyZI+jNBBflI+mn6VB3
U8i/av+TjY/mWD4zuraB+w+dtmbz8stXqOb5HnP49wJe1OL3916NO7Iadlq38X3YX3KjaKZkwyx7
okmvM1I39uAPtCJs2jpaiRV+PWe4TPLoIWt6qHOIcOBPzbMXIAy/OplpmR8Wjurs/qvURdKxgg5r
/n4yLcz6B6hdb27XryRxIDVLEBF+KrymQRXB2gzFzo5JvLy1Zca0YSkx9FEM0R0iwbkrjL4JecE+
5ayBHhXrMnoF8gxxviQ74ZwBfHjtv8U3KF6gNVnLBeViy7FDSJlqwCXnHjPrz6hELqkO2vh3QAeJ
s3nwVPsmQyBXJgd6p0lbcMVgStuMU8ChABhSxv2RwNabYi2tgCwTEWaFJYz03DoEVc2fi+3fUieS
Q8FOcfJhVT9QzkbfVIAw0i1907Lix3kUNvHDsDIK0ZkeZEHW5F7+oqxh6p+tXYJquhT3zPCen8bK
tV2Ol3BbrMl63e5wUNMyV7RSeTbSfnkuwqH2So6FQhYnHsuSFEmL0buttXjtD205q/L8gnYPE1fl
rzneTjVxCG7ViiL+PImVr0NIAR+YeJyHcqZPsgX20H8gnQgqm4fEArmSBQpJyvZYqd4Rxmg1FIcJ
bjJjFNuPApo8AssRxLFmvXft2hY925CZ2oLifCmYhuDY1hd4iDGq3SYmJmsTLfJXg22Q8k3yVDo/
K5oiXDHsKSA7m6/fp7gbZOPOZZoXPUhbV9ZUJ/l9pAk6mflXOmXQPia7mPdhe8soi1o7jp3uoj1o
P+CQ5VbAYVD9cWTTHdgCesoG4Hj+McGUh9LxMjUViQ4WWDCqPptZwfNxfejpB9ET6iuKnVkYNSuM
ZH1lprtJ/4eFE3X5BuLjI84ahI6MPtQJcoumI7C6Pe3mbk1errREl0xxOfzFPPw0c5KbYCrNmf1R
oeekY7aCFacEa+62Trl4KptgKdceDNg9y76id28cbktjpFyOQHiO+EagTyrW8tKeJLwcgcH3WAFk
ZdjZ8H6pmkMoaIUC1dpExA62aDkmoOcOfjGirKHTSWQXNpKMiQGZzCyHXNvGPM/AfCFbjC7sYWbH
cY537M/oQqvCmON/I7GPKsBVnwv2mEWfgX9yonOhuUUtLN7HlLBuuH3KARJ7XEFvLgRleqD5rDLO
+KJnveSV4BY/lg8r76GGIwlYpgVErD19Y93tRy3KHzgK6ObfeaRzyZKhrSADjRaD2AMMtitK6ttr
R58vg1b6Akcg92cNMrNaaDZ63r82rG4mMhjzQ8qiOqyP2EApBjgTt5H4ovi0hSLeQbB95KskyWzc
QFSngKLTvNOzHYm3nN4VInain2Xn+7VRCge4D6twSJetPkH6RWXIHAOiSpvuNpc9bFh0IWsa2L4F
gLHId9Y04/q7MObXndznUCUrr4J+AtM/wz8kgXnAPow1JprmIuwlfboAVne4vFdBYlsjurMIFH+T
hRRu8TDie+XIk/gFutuMO/JjgZQSivZGiGx2SoJCgeB7iExyzZRW7JE/vYHgHLA8Vx+83Fw8Z3rZ
o3m5TvqT+hanaMuuwCYESGMcKNz2V8Ncq1Y9vYRUFc7YsbBY1HkvWrAL5zo9mSYUnTAudco/yw8N
y/2WBSTm1IBNYdUJUE7WYIuBHk8aUJ88+G4Ut2ERkJvnsHtPfX08Cgyaxua72wfgetY0dRgFfGsy
9U7WjGqGseAi2hER4J8FNakl8iFSHRbyCwWr3SgSVRqs9sVLclYjkbnH+o+xadEw5OYOCMcLhS2z
qvXdjSrU0MNxzxdCRrFzOGoc6yOt4UZLFFyEsgho3NlBdMDLS35xyoymCJLcjfGMMBmIQ5GKkLd5
DGnDeaTlP6Tsil4TrGfEDx3KAF0NHFPvkwMQVEyRV0YZpe9v5UpHQV1AqfGlSXKthDlyu0gVBui1
4VnffC4f/e6ENQWZtEsWQKkBZhdb8wBxJ4Sk4c8nxRZuPQhKq7sFlUs/NdTZTnepjbn44zDsOOmp
nKsrZgohttK3c5wgjSpA5NEBN7jdstQLZ27r4PfaybIc6+gNUTdK88q2jywRegpSeEPfy8ze/xKz
yKS5SvVQanNXvgA+YDfk9WAULBWni4IaaknF6oWSKqy5qNt2DVVtt4iUWizBadeGK0GYbq0fke6p
yuQ3vj8vu1lIowFmeywZZ0Sr1hsaHUgC8Xpds05zf709/BhBv/c54Is+ug5I/RMzETIIVQ0YTXgd
BjqqJc7OTncLk0Q+dks6jD5oPyVd+JeXNuuV85JVsM6n3ZRhGQ9t7ZUcy/+ZIVMk7K9ReemS4NDb
ZgjgFaPWsk3faLTPxnYxDfKrKPkh+6UcYJ2HABt3D0eJyq2A+utW+aij2DxNbzU5XDdInifHGA8V
yAVZ+bjpbhxE1l2ysggnl7X77p4P5n18CLvpJDjgQikP7Gu0EmohdenFPI3t5zzvw27S9KYhok9V
H5fOIjOWd+Az7/bbg7y0iGydmrW8DMW5I3n/MlhQksMpp0Ng+X28Dco4ZcGMxi2eURJylfi+fgSG
rYaR19NgUa+vCcshcttBcsHEmftEr+YrmBgZCVC0rRcu7fwoYtUo/Wvf8i3PftTeEnGHpbn3di9n
gy3NBTDT7Paim5jnl2NfZm2Ffeai8VLxMWmFPO75w3vkOUfnT0g6RoAyk3huQeTVhm2iyNKxuDNC
wNLw1mkzma+HAuVpbtGpMLQA7E91VJ6Dyv8hgW/Gdy3uTYO22td1sAEHScOWyMoi6Avq4BuasXNA
o/w+fp0mZxJeKz6XP4CCQZNOzKu45hN+0h5ECYn8idjX6PLv2GlKPwEQYfJCJ4F9iBsLL5RD5Dot
YCi099hCB13muj6crBazJ8zCkh4+rgy8PUM/vwCs6QKo+pm/npLEOqtN5CF8i1Qh8V6bivmq7nZD
4bqRvgm/qO3u9zLmChGS5rK4Hp5L3ambomWEW3pdN5hhfrL3A17P1P418kHJMuKfCDTfyMnwbRy8
a5HdcT6jsZVUf6j2GOjJlIzESNBrKtXHi6lKKjya4hePnq2XttVHm7/q97qBljWB9LW0OdLmOOXx
zA+xTUuhWFNSh6FaO7Od4rBR8Tr+Wk+MJ2wIkokI4ZCehvWkdlSH/scxlAvigjehiGUSUrM0Dg2+
96Z1fuc0xhs8PFsRYxtgEnRV0Cm5YZmdRiLJRqavGJ2fqcDcy6bph0r73yULUFjAYcn5y4DXpkis
tgH9jkNgb8A25VeTbFjxU6ReGibyFKaa0XmcDSd5Esratz2JHRmp4aiJoqbxWRWh0XFkmPt4fSMu
Sc2tonFajmaCx88rss0ZH9rrv/0/n2nIILcL+IdL/7tXG3wKtRavkRfa04joWlaW4sB0pUadJVKx
/gIBDg6mKTmdk17BSmUJlMxHiU7gRacbZOUNh9awLHWTNB3iEH5p5APwr4Z9M8P0dwH7P7FhE1sD
cxzCQJ30wRTM00PZyWwdNJwlclonUtoGWh1qyI/8sPS2peif+7KIdWZuIX44X7rR0xVPihkmIS/u
S9kUJ3/xjP6hGdB+yK80B95m+UkRTeDUlQhEMZc0FWdDEvc8Sit4ZVZaamGEl60uKrdcUWZA1Zav
2wz8E/M/4+xeydwqG1fdaWPEkZq9Zh/t0acG4uPWltmRwQaKcUk2gd3TftKZpCTrdi+9Bd2uQMjF
GUWYC7NT5U44LVb/CPTZkowXnCXqwA7k0ySDBRMuFDbSGWw/Xd5CNlPSWn/YkI8tuh6WYwedNTne
gtPNfLwaDQdePeJrwH+4MbpFO+Vd6NpCafgIxAP+CCVZZe0HjRBicuLjGzdNoOBXStvzO6//R7OS
g350nz4Psjij9co5+spcU2bGxfVGw0Ihi04pf1suxPmki3HfPQYzN9ZH0gL31PzCGmavlbCdmNyX
jbiUoL6kjAkkSU20F5DvFSKuybSBaG6t06Ortn35iojoEVntncJKYqcgQ2PvghW48vCg27pyUD1I
aH2m+rhc6beZR7jdfZB2XabOJ+9aehcl34SkYRZTDiL6lJ1N6I8YNZAzoQBLkVjwPZofIKF2zpLl
ih/JtVGqKs1Mb1Xc8TlPPbwEpfCc/ROoYwt8v6iulq62e0o1EVFdmXMMg/ZmWAngpb0774PKRaX/
XMz4j194CULr2gYJ0pXlLkf95U3o3GNKpw7jDEMIgJCmRPkqqcXGqokjnOnaP1ilPZIt3SJy7QST
bXD7HnIqFHugnnA+f0KVN2N58mjs/flrFGyI+fPOhgHgdrTLuish8H6fcQvwxQ5bs9R5fBsRLub/
8ArKdqUp6pUcwPWjbJFM0oCvoRgCuy5/OSgfkon+WNIM5D82m0MCQQ2iF7MPw5e122Fp9oxzhlXb
bs6th06Mz5veTSsHoqYoTWECx+8IpvNVrL0Tfkde2PKsA+47dC0AcKcoPDCVbXfQrPReiF6Ojh3e
7Nnu7jfH4b8g5ru8DQek1Ho8PZgyLlo9Y5lJ9pVusVJOWI0a2BGJfRNqVYcFenYqGK5wzh3RnuyA
T9kOSJfLD442QxgK9JNHxzdixXGu23Tt1xKNU6clnma4j1BDcdQpijoakOsljoGj01veEz6yjgWJ
eiOyTpCDs60JoL705r9vm7cQYEXAnrlZOxb86QTXau5jvyQusl0QNaAWNYIG9e0Tjlsw2KBiEpdE
7KixLLtyKqBeZAnnxK8JHcj/T/hhoKRdLQzGyScaIgpZAnOekc1GfjTWTBoWIm0viRNrKNQ48Y1Q
vHZ/KorawopZZjA3ttQX1aA7jrIAZv5AHnHbDZBT2R+n0oI20LLuNs6KcFhWqL/iXZBNP0GYZzKQ
/4E79Xbz/JsDIIEtosFIcTFxRYrDLiYDSHZid0bjcqlPdSoPen0y+2QygkdkkGxAEbxAfLJjeBqb
EpYX/NQ7/PqBUfDxhIgvbcoHXwt3/srlxKb4M8+m627pL4cNIl4zW22as85c1omUja7UmnJ9XIhJ
LgMcABeY3onPSmSPj1PZFhIDmua/VZeZRRhfAOHmFs17l5k5XYp9c3HDHMYruCJLSidEYP+WZEqO
OzqofgGtbOHQTFwC9JoxViknZPGo/Eej5CCa47maTb8YP/DkCJ0a21dKA2VLPaLykBngj8+DI9Vt
ir0JBJNYzUSq9sDOt4px/EQX1F+JXRcx14kgNhkyuRU0ASme7OvmWhb7LszSXIcJ/Y1jMO94mZMr
gan9knPIteoDWApS8HYSegkJmQkhkLE02rNWu9R+BXbj1BzBMT4idyJw3lFrOVeNjxjmF4eChzFY
ScOyIWIABqlzKFMb8egKyBxXGJtY0rMusRpq7d11L3skdiNh2iTB3/NtKROqidUd8tr+BA/lm9BB
eCQjuhEgK40xA/ItR+y7Aivf/3KDHEa6oTKyuSb8t+x495emNMPZkGynOuqgzTBJBdD6gVIQVl4z
yCAkUqjy2fjA7/dnnwTwnpvYobccAmhdIS5r2HOMh/oxGxR/G3fv/wcwutbXDvYRKYDG4Ssm1ZLy
JmVeZKZK3y4YWBZfay1Kvl3wu8PtZ1Oq6a/u2ynNlVpZdiHC6oaNBwUqMAiBlrk7koe0PRA/VPQr
3fyvI2aY20e/ZLTaTlPR4DGKWHNphBy2hRl3/OIcmDEA6vtNZHUu8PVdIy2Sr3ltqrE+PWtqK4iT
EUQDI1bQ1IDNdMIRfRBbX4G9yHOzG38q6E8pvtYZpRGPFLVXfY20EwK+/7cDyfmkFsY5uIdLf858
m4JCz5ue1qcLtIEe6GyXKTCikM2B+nh833zld/nYLorV9aWUTK1eOmXGOznQVKqzG2ruqbsPLue3
nkyh1BWEWvfVk2wq7ELSJKitpCjau01uObmyiBSXn/1/Apr6xHwYG56ZBv5F80sFGnpYx7SmMaIa
vilG8cmKnFxZ5bLfhkwRcQoV6/rS0JDGhO64t+2GxyS1njPPOtECbZMnU7zkdnficUb03b8iKAOC
ZVpPjtjLjS9jtYv8jtnzfAf3/DZhiX/I9gMZmK3MWo+99zlTFYujKUZ0Fd9Fy5BhcDry2HKuhHeC
2zGQSjbOSyDDOl3c7Bxz2ix9FTh7bz3ck4HpSO3kt6gs/YEHQNamc9mp7Y5Gtm/VztOeKFAorROc
RsxGBvI+NTXhmqdgl0qsWG41KamVzYQAXymfdAVFBgbSmRJSsXA9ZaIRiKFL8shNUCi7YeeyRsOp
XBiuQx4Nc1UtsifY5LGzcALZ83rOqgDkmVhIy3R9O5dGmxAQOXjA9nnS5C4/X5GVJjev+ym/b9UL
uQemxx+0V7dn6mBkIPmUjFPo+u2UMFux4Ii0hhQ8sDBbdqg39jcgrgUru+0f0iYazM7eK9d0f/RU
JrJPbq5G43ejSVzM/9dIOXxGQVbZLJ1wEuda2BSCSs4XZZxpCkTAVU4IeOn8ueVvqXNBnYrXWf5k
GcZ6ur1uGS9Q4Tc/QmxRxDdoEBRwRV2S/DGWOpfmoaCpASOowHgQ1inH3AhvA17XHjlx4H4U7rBE
WbJV/0ZxJ65eK12XQPDPilvfZM1GXiXoD9koiDqIPlWsm3W5B1qr9PaCg4BbZ9diYEzcgObltlxX
Ezw1CZet9ZdzBiBOEp4LAnJfMO3Cq5HKZbky33vN0FUokW8MIwgL/ki13I1SGLhDG1gEXRPTCiGr
5n04qsjHcUEtb6BDwFDuaZUjgVjK4IFMq1ZJ4EiUwkhAzn/3+rr0d2SS163NE3kByFhQs2wmjT3X
jmRr8d5Wo9d6WMJzucFFCNaUmpVt2ibQkNXdHBP7CXv1u/7vPWvdi5u5fKyGMxrDGs2cJbRdfI2m
R4TX2gAGYHVIXnfJ4KcZBvwe10HZUa/QFmpvdYOA5uN0tn3nQLkOLmP14azOgVHrd+DOegtl7qsz
blT8Vr6oaMLTIKCXOohSjHFoaIa04EDHw+4k2uaCK3Ccx1jyRi5/N7HS7mGvff/Ly3yug5vG09Lp
iVQM9xa6OZiuHuP7y11LBV/6JARUG2KeUrrn7DScRaPIGjo6EhFIzOoRaDrF52UlNqVn++Ds/pWg
x1aMul+EiUD2ZNvVAfNHJMTRG3jVmj9xqAqqkKG37yFp427bB3fjDQ6Hg08pUIKzgSR4Wd7ulsXA
tOTd3e+VFScw9s7RLV1hcriwOrK1CVlGUOmZDXCgIPxsULksnXh2xvcbRzw62Yp8/9IvKkLc4KOd
g86f0KBl7WArHutu9c5n+Y0gh+ny9xQADO7fVn0Wj9Unov2I10ECZILh9iGZzKcI+UKnBg2o5KBs
uafdy0kgEYNOACJ6Q+acJa/XMAJt7gir560OfZvNXhwPqHPD+ejZgmSqw2RMewnNLLjhsAwQsPvH
c/VNs3Eyqez6HyeZRyBOYtjGpr4+SOrpg15U0GeEACddVwMAXQYhUxiTfo63JVfYcYj+BzIwTS6K
d5T22ne9xgh5a1GSwC/S6i85YjjxLy2BVHiKSRjrlXqOf7tLBUMJTDRncJxoOc/NhP1n0wDX534f
COi+P4V337K5yT20o2fPGT9ECgXjEsFbO8rNlGuxsdvdBGU2ooIZ2dsa5/sdDfGZX77frUkaG9uL
5JCRBKVUz4wZIcMMxxJ6C2h3Pn091U10WECSlH32xSLq1LchSsqhsyjrtkctshl5suQ5UC27FtTX
V7gqaLr6N8IuXhOUi0QJnIxSUNmQTAc5bqufMlkSd/dO8fLpAz0uvOErOJ5RxBnnRN5dBoGt5GxG
4vum8iZYOCMFF1n0pWUdxlLMCP9BeG+25NmOwnYDftpW5pMCOOiMnX7wHrBWvdU18Ha2P77TIdZo
stuk9fkUYhQzCij0ANkulOevGW8lp/lmpoOi6Y3iJvFrXjZ1oZS2hGQA4RDXYszahBx0ox4sFWdl
dRmS/6hqZXU+dCCZhp7R5wdfIbmuV3/ZdleVFXRRACqOfQ0iXLsUQ2Qp+PDoFo5qsF1ObYh0L+g3
a+LoNh2eOgnlpmpLONwjV9hH7LvTnM22YaKO0kNQake1bScA2h7CqqkqugZc4BkQzsdXmh20pxfl
4yhuKZgse5aH6C5hzLAtnyIvcJAsTeb2T3RxFicMf/Sd5Z53528ORGwYuazoEwFdmK1hPH9u/Rvg
UUb+f6GkkDi6maXMP/pjmnBu5gGw9A2rMmGcL5KoOnt6fHAmgBbYkw+Wla80K/CtxeeOim4bkHde
DUyXVaIwn0snIOi7USal/Dfl4GIDP5m0uzTPZRSEDQTwMbThsSHQ5XpRXkQ7ucgzqmqy+7pCje20
GtNJoXrI6LTkwIB5RwNM5nCubrcJVRFS0PDplvxHN3K/CIek3siOKNNdcW2T85i5I0qbfxk6wK6r
8lAHMNgFq8Y0Boh/eJSLqOs8rE2oUTALBmiRKNdehY2tUeOp7iLu2hjzfgnSNSCatghaZ25Z0E4m
4thvVE7tuFNI4D1XhwzZ3xDENktS8le3ta4G1uja0pCqbXbhox4+G8AwIL/oRBRZp+8hKdxmVJ2P
WPzbxPc2kgZ6uOpyumCOmEMN/TWzRZmSQ09iXlBC4qopVH2MGdsVi3J3S2Xu4dkm5LJxQb6HYmr9
V6UyeAfQigk0aauiJ3g0kExl/U3a/u44DHmziS/Q/FnsI74eQNE/sCkiw0ysb1kacKhc0fPl8e4Y
236k5muOO2g1I4M1mSwK+XjX5hFtNSDYZJ5MUv5ElphSZvLrP6jVqZpnGt8m4HFz0j1JzcZR6tyo
5CNpA3MLGTUiOM/XMxjWZNtC7IvZxVA0P18PYfkilYvy+1s0UB4wWkOZsUQgbqcj4YtJ/1Ycli8y
KaujoSL4nnMrBxKzc5CYdm6cJt8AJVGv3lmfKv6TVXzeybvX6KaHyENwwFCCPC4JP7ctvy3lkkjx
FknvpF4qD26Lr81fMRSLWXe+xDCSywNIfg/yvGdEoVhac56KMYYImrDaA4y/SAdHm7NFz1fOCoWo
a13BVjsrJz1W8DUom248+KmPZxs52OkyE23A+bXWil84brF/z+jD2IEc53aHnKoSR5gdDWoRPrv+
gH/4bSbtSDjSwgyHCJusHNev2/bys8VEEHIXi2EDLYGDMvgSYbuT3PKfwKZuO5KyG6hp0FyVRfpb
UwFLXHL4x/bck5Ibg0ScSYBISYCJxGhnmoAJeF5HDpNBeR6RB3Y0NjElkeQzx0Z0IGJLkb3OvZRj
cKID+qvENY5LI0MFQ+I9dOVrojKqsDPJArxRTRes8RGOxWQEUwbGkMEDedWlGhazvXmeC4Tjzqe+
e44EW10O4d5XfcqCTlS/Ub/KjhjUOwC33daMUWBZIeps5KAw+iFGv9KcO3z8j1hjMI4gMuy/GoOG
Xx5WUCWhS83cn+k+OIUIQQFVHJpfzLNbT3tce4UCV5hu1loyc8Uk0LiD2gS/jzgAxjaJjCNHR1FP
/iV1dbm6haeunOSh2rmqSCKn/rFNOAPj+bzqnvkqZSOJmhlH/UuMbOh/PfoT1zbJAXJr3WjkfSqb
wA0J/gd12zTi28e0w9XAeokrfXCJh+/wpKHi3x6bfEy5c97htHoT5vE3e8bxeSHcT0o7Q83S37yG
E4RBYjMhhe9m8jTN+gzZ7qx+MMITvgbWriRaCnncKAM7Kef5wY9YqIbRaJdxokRDmMcp2/lL7hLm
RG82qEXd4VFbc6ZoDAnwabl/5MAECOSjN3RDS5Rm69sJS4MbYpKbntSLnaVuIUkSbBxqHterokA/
P//w0W1OKGXfFyFDDOM6F5fnUv4EL0ve1yTn/uZTlkloXy7eCSj8FFy+7FeiGPVBdW3lGdJLH1xf
O+RZxvh694/Vz6Cqy3UvA7sfD2F0nJyNidywNz+CTTVxv6CcIxCnpQKzZK1u2K5OL675X44WoedL
w0+DZ1o8b30YXbiK4MDMiNUL6Vozru88BuCD3KY+owbGoTw0vjlGyNdB2Q6HKtwz6KvmWWZ/jU/T
jtH7hk021IImn+WWrlmVU20Yy/VkVitkBhv+Vi4psr6U0Oim40cLOfqNykNoq6WDlwYjSYwtNVmw
VVMuV+kz6/bNkyH/Ak0SvFQuNE4Fy8UednCB4/5JzQv2uUpm/vxuCn2uRMs3XgyGKOdOxLf5C7OD
0qE8VLrwbp+9WZhsAVvChyaZeHaM3jfqr4CcAQyUVsLta+fkKLzg3D3Dz/M4Q6brPLchpQMcX1GZ
9jzfA0t49fqsUZBTkKmZ3/UmdJUFUZkG/ZlIzLE7iuy/xcz5OFNANThxKqKjoEla7t9Yxuz0C1ZU
zlpuVlGEOXfC2xxmWpuScwrdYbCHkGRBvtK14/cm7dp9FshkAv3lzKllUVh+DO/15DgLZ9MpRQTU
GwuOOSq4A6cn80m0+68/fugEhK5hjQWyGMqrJCqqQwn+twHXgU2fD8LHFD8tmoTO3F4m1wy1S0Ys
znFvuu1tn6a+c7D29TBZ/V2Hw0FG/4xg+Ii1AY+ft/7GniBEOVSDv7rhDnULJ8tK+xUppAaN4ggz
Or7JDmEUa2T4YFJMfAErkVssGJqzfHeuGUN+EdbK6ke4xGXwPAa0dOtPKHRkovXEKjcBWOifwU7v
jkfBuL4b5bOPz9Vsg1K0gkrOO1rxcGoRDAmFCLKFDaChLyvw7Aa7srNPI4TbDgur48rlEgXHJe+i
xxqmB9i2u7h+rA7/ssIqM6IRnbt/mMGB9o2mbJ0n1Kpu2GgO7gRZ1Kn/9la8j+wu7d2SWUW4zimQ
VH/88w0GN0JcjMwX4vSH1ppSSDs/w/NlYYDeNYwEnsPypC/2jHJQR/1yAD7iCD1I+4otJBM7Fegr
lZE9uQjrwDfo+JKmh4G/7KvpzdM1jDkHBdQlCP7I/+tlfeq6u7+zuCssh1Xc5lthglQpuLkVJNq/
hjrhAxWYXR5nfAsa+0zKBNfQV77HS4XL5AURWY/CVpEdN+5PSLDaE+OB44uWFUIFQ87swZ22vcwL
nqJaZI7J2bJs8Y2pymomRRVFdlU105LRl3a4ktjxa6UoLvyCi/Sia6MAkDwLzUaNg9TzSNJUrgqc
s8GY7oPAbbCvyg84SirYNN8TpjueADRcGCstXepTUi/TJlwyuu7BaoZKOi9F7vVFN5RU88YaCRY2
FYXlrQLixvlBNaBnK+rfJDCU0Vu/MOiGlfdv6pyz8LH5s+bGQssFfvP7tZUIsCCRbdW2ez2Q421C
x8qP2kL0ZuXLg0e4P2tcWevryY9fSYHQJu7/POsgPipoEtyDuyQGlANfr075pYCvZVVDZDOv6OCd
8gtoC3u6wKw8ySYApdUfZRThF9rxSX+BZbi2pF32C34q1FwrDxtUD6NRwN1+nF6EAAhQGBVfqOnr
sgHYAWhxdSSKK4x1+iLWvFO+NR1kr2RwHOLpMW1eXrCAVHDzKLM9lMWy9TMx/rdhumi544R+w5+j
vq5qGYbPzHIVc/hPUPh0KHLrBdVZEWydHGwBAj6zWuVbsFt6S3uRUY2HaUBSN2ACwR7xD9tlc+wH
Wg6V/edhVifZKv9fvDdKMKH2gP+9TmVuyqla0oEh8oxyD+1v/Za9leC1XDhZyUAgZ1baKPY/tjiG
/kBeaqUZKwqwvPGQtPIH6Qp+DvFLkXJuwGya6cN0FQHVROwnNZGfghnTLgdQSNWsNxPdpbxvAkuv
fJnVO7MPuxSnJAFgHRVMzG5TU4s+i1rIkEBFizZmAJb+4dgqacyjHWkYayqqQy7UTUIyI7uklPrT
9BMFfcwOqbyLgb9Cn/SZsPZdiuXtvSiHPpAFu3qZMdh7TNygORIbhKGyz9wXcdVSXf5aGC9OjbsG
24jjV5N7d/6qA6xuaKiZs+Boe+qa/MHAphhT0RsfLAyPG1zMfkJ1U38iM2D3WXl+87XdWbFPKj6q
swLi3gp2hdr6DHQ4eKZYPD080AEvvggzcH+Ld3161I9W3E537LNQp1q1/Dt6w+XFdemBimT1+aVf
/ECDiv5+D7w9rl4CNR5t0VwPQVeicGUu3+fW2J89NWUCDe6eyOqlPinvpeKXEYLW2LRz4jJP3VyT
n67IPEySrOhiyBKd9/K7jN50UzydDeX+p0E726ZNMTgHEs4w6zo3BIFIU7glqchVrX47XuQS8nUa
Bq4bLIuVY8pAeMlCxtwcQUmSSj2NhTWR7S0LW4y31VXMhl3j4Q46iIN3ktlDWCc2g2evFb1Q0Y7O
0+pZ1q/f4Lz1AW4ArX2/2+jekmlHBZGtWBND5RVVruR3ELwguZF3Hc9t4Knige0QiR0RRZ8j4e4D
4bZdRq9tHWu3cLK3xQKus/WZP0B0qXGqv+FwZe7Umz0zz3P8mzwCkjj9JwfDwLm3c3qAlHDq1hds
nruVQNVoauu0/EafAEtsWb2YFBfHUtGF6TeJ6FgD9W5M9xBXBJZFoEJRdx61SahPpNdsAZQfHZWg
kRHy60i+TmiUFJbtdUczHNPapBiKhMymDah+ZY+l2TPxYxmmPzw/aYBu3PLEfH0pGx5Le6LueG8Z
/P05XSNGufKrq9H7ODHEBHgMr2qkKlRnIJsdiRDONGXBqu0+25cTifpUFpS9o7G+2N4YB0FYTrGH
v03xe2QfHTbOVXwlkpxmC3W5vwnVj9BKcYxHaiHuruK65ak68xv5ThZmTMe8NUd8S6zvmeuTPyrY
C+zYbrAyi0R4Asr9uyD6T2y/JmJ/c72Lbwz5lz2BLWsnytTH0XnvNXFc0TDzxWQHvNt102BgqN11
K0NEYnqYQKf/nTvKBnbG0lXYBpPMsihrBdmIlwxvt7LdeabVUfENgRPs91/+Mo3I+WG6+7QDR7fK
V7p6mV0/ExTB8tFczEGnZdEuSYVGJcIZSyfM7fr+5ktswcTYnRl3mTi/P0smoG4ZG3cpOSVPuK67
1NPQToOmKQDM7TE5ip8/wdNalfsEMEGn9cdQ92eO0S0oVQk0C5064dzPq62/0GBdQMEGuVl6T80k
xg28jTrw34mCqfIthSFwOD0q0gQXnvrnTmb/1asqHvJO9ZJ8w41aZBIxUp6EN+DYsWD6m1RtztEY
T3PVbCOt/cQxyb7LgFXaphibtDGdpEiB8ApZ06O5+XPpb5TibjztXEgzZKBCkX1O++vNvjmSVsx9
3bSYHjKX7vueuOKQ5bA0v2GLJB9l4F0lOaLh1aO0HjyzhtNb8fNUfhgio7V6stcjABcGdywtXNzK
g3himxiY+E24yxO8pR1gG+EJYWtA68kdsBRFUEbuIx1+cKiW7bgKge3oH/MXOVNPXzATcEvFFk8m
FllrY5OwYeVCPuAJWLBhpkfmxeuaFWb8pG7wanIIrWXnytEx9uqtw67CWItSro+5PDEMRXeram4R
WhtJMGQFDlKS88yU6ZXGjdZZKRALBq9M4Rj6vf0UQcmjdhU9XQc5bjNQcpj4ff/Ssk4Vs929GsE7
TLuY3x3Il18xDRE8NmilKcfSUlQQyD8v0P9c1a+DWX21Yj3130NTkizgUqtMs6g6vKc/AEoMESkM
PSXoRbjbSg46Q3Upci0WmFhTBc6DrdCsruZoxzXgc4asDdEcGyr17XmzQedbSjbxNJLD0yP1bqI7
FdXmlsDKm+91c8jI2VjdAAYd3Z0UMhRD5DdmeqYUc/z8yGfMXBQT/EjJiSvyvbqSLX8GUtZCdXKR
+/zXXBuNSMVx83YiRuRUQAzK6JMfLB1IN1y6U8g5eVxcIrZYoErxLxmPANHu4UI10nHE0vjSI7/x
Xran7qL+qVUqb+vzlNTqrwe/6vqs++9b314/3iR9n4vjzXvkaXBcKtB3Vz13f+AekBMDIpKyLYXA
h4qCcv9bXljDr9Wigg1d4ygNYzUPrCwGcbL5cryyMoBwpU0p1pG4wmfkJnmfV8VZL8e5i7yQ8ruj
uxkA+09Bof7jm10rxeulvEo7cbMzv4G7Z45s3Jg0VOaVK0hBQBeZ9/5jvPXZWrkGSxUstCyG0B+6
pb2pUXl02iarr3QdpU1tQpfNFo/DhvqebXSDMnbhlO9xzXzh204mAU3sWFUGtO1LyRtX0+OoJ56K
X1pZu10kKPz6kvcR70Lj5P0GlsIXlRMOCLptokg6B5+sM/ECyZiz69Im9sFl6BDwuE/3BvdY3f0/
7pBpRMgBSVxMGnO+KnwQ9wSVaz1zX9A4prdkP1b+Hoqs55h6lzUJ1Wsh6+1iZROTOAl0We7qoJJB
DC1iLBZY7QxNdKNRgVwEL3v6+TUTI4ltIwFrx8/mtcS/jgeHb3jb2Rw2krkKY8Rux1Mzb6d0ZdAB
pmDvFT/yEtHaOLlQU7k8Ng/C3z2YWtKOSI14eRGaDU5zM92VVndGwmFltVAjQsEMUPMipU5r8FoG
VoFwEs40uVUlA+d0zyGRqryUnLTHSf3nDARPultlk7tCFeQQTSsz1pDu5CV+WsPY1hbHmJF1OKje
RWiNF+xu92KHhYs8Bgdwxix9bvgqrHgM9I/94cSWat5Dd+3lzSWXnlI7zZYUu2uZ0PUsWjNAQxo1
T98UqocP5dRAgalhHOSI88fYg7SwmaS0Zju1PhkMou3V3FeX2HYAPAfJSzkxutPcRt4GxQxpdCoe
ncwkzxO/74BiRp9WY7GXJN+l/Guomzu77DJGmtCWeMxWU0bxSo13oIIOd6qF4ixKQ+DmSba49lzH
xxLmvObqR9OlH4WjWjxOUlpn5SImi7M+W/x2QOcP59u71cbJx/3+cc4nGffOKf8CoFhaeERaOCnN
MNCfiS1AibV0xUKzvOf6M3rp/4imKEsojA/KgbXY5mveJzsrChn7BDKSS574pr7NL/j04f7WYkIM
UMhze+FWn4I9kp64wEsQdAyXoBSHkUM5kZ8JmUMYj1l+8RrbmGyQxNlPgI6jpLrqBy/pvEiPuuW3
7bLA9YqtmpooPay7kY7Ht8bSneVu6kF5QYPOiTlaf1mgPk+EIyrSZxNWa5OTb8yjKKx9n1e28F9g
3XKos+m3j8zxoHr2eV1O4bU4OTlKcEVE6FReMeIjwWM0j21TvvnIg+/UibYNTjvlSsDMZdOJxTjW
VV34K4o2/x169B6Nin4LiWe43egMEzEjTiCyGMys5Ze+kfnqri3aHgjjIwW6vQP5Ah1zj5qyTnV4
MVdkEXeuddS8Sp7Hhkjc+dc3WfV7SeUKP+/mMAW1m0rksM978Z5u6bATrULz+EfuKHf4YjUySXNJ
uFhEW4dY3GdospwyRTUvZjMu2/tuqVYrYWEf7tkjwdKcMRdAtUguZzZ1oMzsUpBNOjiKbAiEyRuQ
Od0IO/ADSAbeL+pTHpo0LrWgcsPeIGDC4H0QKAdRl2O1sxe/uOpY3GcTEr+0dUFKqqODFxxXjFjT
iXOjM1m/6DypTlmtF8unDDtcwTWNp7VsUSlbAfx7Nm5QLGzRGDLQevgaA8fjKDe8LqklPlcH7NT4
PxR1D8Cg0MLlU3uHtauTMJrB7Jla5vmYtT1kfFhbxv6wT2DNXnAGeQMs3621IosCFxodZu69ggYS
N1UaVJ8puYX9DrOw9KlTnL/3IKkR7DtKnax+MfcpsHbDrjEXGHjMv+FKnqXM+sihVES4t2HwmYgK
HXOWi1dSb6OXqDmOz8MlPWyoEFBKMqX/rgoNDj3Uq7y3Q9xvlLy8ZhG8D0ANn40FnbB3PW0r8upO
gl2nAO00W1oK/Ih4ihMEj35N+7LHL+p/x9UQGt38qhgKbgZbI9io+JhyBHIO3gIXYUGfFGMKCrsV
PJ3vCMZKmOFTDCM6DEdg/0SrIWLeO5KITqPRhf2AJokETj/KLB9m1YeYDS4h9uB5ixc9v8qOn2SD
+1EPB7KwLZG5AZ2lHgqOHA2fbg7UhJH+pRd7Ae6VsGZXFi+2S16dTQPislYXEYmV13smvYVDvM22
GstQ8glWTyjptUYs7r5O6Jrjx9bEWdhpG4DarsB/z6a4JxPT90xoniyWKq65kdox0ZuGUgDszBpv
+2tioeWSJLy2f5/XSkpBE+X/zdEMfzTH1ycx+OMmAraJG3ay0dSFpE6+JBC98BwHMbMWi2tt6X3x
A8UY7U33XSROuRkBntp/bFSmJGEX3esMNwpvj+I2dMO3+XjCK9+tCxwNSjQUqqFDQdaukwT2I8vj
ZIxUFvUKqPsLnQmWCMRGx/SUaG+g9Q6z8HEJqtkRr6+LAp2vi9V+VM1gyZ/ON9/HisJuGmlpuWAe
c03dxSZXwqoBhS1IoZFdPpxxgQ0c1WAaddwpoqnNzW/DUMvEXEzeMJ1DabdcyoLRfEbvrzFFXplO
/rD9V06HsDouIXMFQ9nWSOPBrejewJV5uCPabR/jwXMlYcGdiOVWRqLKSODlEDDgjxywvUMLXYtz
L76GfBNe7DDiBh0hqJeMxbycgabF5qBA3PkWffYtsWVIaWLEm0S2WKO9PjqhvOnTB1NspQSykWjl
4PEEVmqbb8+p4ukB0/QTOjG98d8QBOOU4Bn+PGuj3//Y8N5s1onASI0OcIy9oQXt5CxuDdJcyOJW
xI2C7XHxVOiayBPwbYuNy2kMFMcu9zRKHJcyveqRNVyD3NOZnsd2HN5o7vt9HPdcZDq2cHPDFHas
VQ+TmXGEJfxz5tCcqE0qRBuwV6V/HqBsljZH73U1AgVHA6J0IbJTvODCikzO1wlHe2iWCxUs0153
cXRicQ9ZdtvbMhb4K+hD7s49+xX19SAQrrdYZzzggGhhVZIn/y02/aFRMvC3hjsOI1TrxRc+1g86
uGXChqewMdaIp77ykkG5ziB/LCYomC21LwA=

`protect end_protected

-- ********************************************************************/ 
-- Microsemi Corporation Proprietary and Confidential 
-- Copyright 2020 Microsemi Corporation.  All rights reserved.
--
-- ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN 
-- ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED 
-- IN ADVANCE IN WRITING.  
--  
-- Revision Information:        1.0
-- Date:                                    01/22/2021 
-- Description:  AXI4 Streaming Template for synchronous operation
-- This template assume entire system and AXI4 Streaming Bus use the same clock
-- Cross-clock domain handling or back pressure features are NOT supported
--      ** AXI4 Streaming Interface **
--      ACLK            All signals are synchronous to this clock
--      ARESETN         Asynchronous active low reset
--      TDATA           Frame data is transmitted on this bus
--      TVALID          Indicates that the source is ready to send data
--      TREADY          Indicates that the sink is ready to accept data
--      TLAST           Indicates End-of-Frame
--      TID             Needed for switch
--      TDEST           Needed for switch
--      TUSER           Reserved for SOF etc
--
--      ** AXI4 Lite Interface (Configuration) **
--      ** Not Defined ** 
--      
--      Questions / Open Action Items:
--      AXI4 Lite interface needs to be defined for control signals
--
-- Limitations:
--  TID, TDEST, TKEEP, TSTRB not supported              
--
-- Recommendations:
--              
-- Update History:
--              12/07 - Interface defined
--              12/10 - Initial version
--              01/04 - Update for sync interface
--      01/22 - Update for TUSER support                                
-- SVN Revision Information:
-- SVN $Revision: $
-- SVN $Date: $
-- Resolved SARs
-- SAR      Date     Who   Description
-- *********************************************************************/ 
--=================================================================================================
-- Libraries
--=================================================================================================
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.NUMERIC_STD.all;
--=================================================================================================
-- AXI4S_MSTR entity declaration
--=================================================================================================
-- Takes native video interface data and converts to AXI4S
entity axi4s_initiator_gamma is
  generic(
-- Generic List
    G_PIXELS     : integer               := 1;
    -- Specifies the R, G, B pixel data width
    G_DATA_WIDTH : integer range 8 to 96 := 8
    );
  port (
-- Port List 
    RESETN_I : in std_logic;

    -- System clock
    SYS_CLK_I : in std_logic;

    DATA_I : in std_logic_vector(3*G_PIXELS*G_DATA_WIDTH-1 downto 0);

    -- Specifies the input data is valid or not
    DATA_VALID_I : in std_logic;

    EOF_I : in std_logic;

    TUSER_O : out std_logic_vector(3 downto 0);

    TSTRB_O : out std_logic_vector(G_DATA_WIDTH/8 - 1 downto 0);

    TKEEP_O : out std_logic_vector(G_DATA_WIDTH/8 - 1 downto 0);

    -- Data input
    TDATA_O : out std_logic_vector(3*G_PIXELS*G_DATA_WIDTH-1 downto 0);

    TLAST_O : out std_logic;

    -- Specifies the valid control signal
    TVALID_O : out std_logic

    );
end axi4s_initiator_gamma;
--=================================================================================================
-- Architecture body
--=================================================================================================
architecture axi4s_initiator_gamma of axi4s_initiator_gamma is
--=================================================================================================
-- Component declarations
--=================================================================================================
--NA--
--=================================================================================================
-- Signal declarations
--=================================================================================================
  signal s_tvalid_fe       : std_logic;
  signal s_data_valid_dly1 : std_logic;
  signal s_eof_dly1        : std_logic;
  signal s_data_dly1       : std_logic_vector(3*G_PIXELS*G_DATA_WIDTH-1 downto 0);
begin
--=================================================================================================
-- Top level port assignments
--=================================================================================================
  TDATA_O             <= s_data_dly1;
  TVALID_O            <= s_data_valid_dly1;
  TLAST_O             <= s_tvalid_fe;
  TUSER_O(0)          <= s_eof_dly1;
  TUSER_O(3 downto 1) <= (others => '0');
  TSTRB_O             <= (others => '1');
  TKEEP_O             <= (others => '1');
--=================================================================================================
-- Asynchronous blocks
--=================================================================================================
  s_tvalid_fe         <= s_data_valid_dly1 and not(DATA_VALID_I);
--=================================================================================================
-- Synchronous blocks
--=================================================================================================
--------------------------------------------------------------------------
-- Name       : SIGNAL_DELAY
-- Description: Process to delay signal and find rising edge
--------------------------------------------------------------------------
  SIGNAL_DELAY :
  process(SYS_CLK_I, RESETN_I)
  begin
    if (RESETN_I = '0') then
      s_eof_dly1        <= '0';
      s_data_valid_dly1 <= '0';
      s_data_dly1       <= (others => '0');
    elsif rising_edge(SYS_CLK_I) then
      s_data_dly1       <= DATA_I;
      s_data_valid_dly1 <= DATA_VALID_I;
      s_eof_dly1        <= EOF_I;
    end if;
  end process;
--=================================================================================================
-- Component Instantiations
--=================================================================================================
--NA--
end axi4s_initiator_gamma;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.NUMERIC_STD.all;
--=================================================================================================
-- AXI4S_SLAVE entity declaration
--=================================================================================================
-- Takes AXI4S and converts to native video interface data
entity axi4s_target_gamma is
  generic(
-- Generic List
    G_PIXELS     : integer               := 1;
    -- Specifies the R, G, B pixel data width
    G_DATA_WIDTH : integer range 8 to 96 := 8
    );
  port (
-- Port List 
    -- Data input
    TDATA_I : in std_logic_vector(3*G_PIXELS*G_DATA_WIDTH-1 downto 0);

    -- Specifies the valid control signal
    TVALID_I : in std_logic;

    TUSER_I : in std_logic_vector(3 downto 0);

    TREADY_O : out std_logic;

    EOF_O : out std_logic;

    -- R, G, B Data Output
    DATA_O : out std_logic_vector(3*G_PIXELS*G_DATA_WIDTH-1 downto 0);

    -- Specifies the output data is valid or not
    DATA_VALID_O : out std_logic

    );
end axi4s_target_gamma;
--=================================================================================================
-- Architecture body
--=================================================================================================
architecture axi4s_target_gamma of axi4s_target_gamma is
--=================================================================================================
-- Component declarations
--=================================================================================================
--NA--
--=================================================================================================
-- Signal declarations
--=================================================================================================     
--NA--
begin
--=================================================================================================
-- Top level port assignments
--=================================================================================================
  DATA_O       <= TDATA_I;
  DATA_VALID_O <= TVALID_I;
  EOF_O        <= TUSER_I(0);
  TREADY_O     <= '1';
--=================================================================================================
-- Component Instantiations
--=================================================================================================
--NA--
end axi4s_target_gamma;