/*****************************************************************************************************************************
 --
 --    File Name    : mipicsi2rxdecoderPF.v 

 --    Description  : This is the top level module of MIPI CSI-2 RX interface.


 -- Targeted device : MICROCHIP-SoC                     
 -- Author          : India Solutions Team

 -- SVN Revision Information:
 -- SVN $Revision: TBD
 -- SVN $Date: TBD
 --
 --
 --
 -- COPYRIGHT 2022 BY MICROCHIP 
 -- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS 
 -- FROM MICROCHIP CORP.  IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM 
 -- MICROCHIP FOR USE OF THIS FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND 
 -- NO BACK-UP OF THE FILE SHOULD BE MADE. 
 -- 

 --******************************************************************************************************************************/

module mipicsi2rxdecoderPF
#(
    parameter g_DATAWIDTH         = 10,     // Width of input/output data 
    parameter g_LANE_WIDTH        = 4,     // No of MIPI Lanes -->  1 indicates : 1 LANE,2: 2 LANES,4: 4 LANES,8: 8 LANES
    parameter g_NUM_OF_PIXELS     = 1,     // Number of pixels to output -->	1 indicates : 1Pixel,4: 4Pixels
    parameter g_INPUT_DATA_INVERT = 0,     // Choose to invert the incoming input data -- 1: implies invert the incoming data,// 0: do not invert the incoming data
    parameter g_FIFO_SIZE         = 12,    // Fifo Address width in Byte2pixel conversion module
    parameter g_NO_OF_VC          = 1,     // Virtual channel 1 : 1VC , 2: 2VC , 3: 3VC , 4: 4VC Enable upto 4 VCs
    parameter g_FORMAT		      = 0      // 0= Native, 1= AXI4 Stream
    //parameter g_CORE_EN_DIS       = 1      // 0= Native, 1= AXI4 Stream
  )
  (
  // Input Ports                    
    input                                       CAM_CLOCK_I,                // Clock from sensor (Byte Clock)
    input                                       PARALLEL_CLOCK_I,           // Pixel Clock
    input                                       RESET_N_I,                  // System Reset
	  input [7 : 0]                               L0_HS_DATA_I,               // HS Image Data from Lane 0
    input [7 : 0]                               L1_HS_DATA_I,               // HS Image Data from Lane 1
    input [7 : 0]                               L2_HS_DATA_I,               // HS Image Data from Lane 2
    input [7 : 0]                               L3_HS_DATA_I,               // HS Image Data from Lane 3
    input [7 : 0]                               L4_HS_DATA_I,               // HS Image Data from Lane 4
    input [7 : 0]                               L5_HS_DATA_I,               // HS Image Data from Lane 5
    input [7 : 0]                               L6_HS_DATA_I,               // HS Image Data from Lane 6
    input [7 : 0]                               L7_HS_DATA_I,		            // HS Image Data from Lane 7	
    input                                       L0_LP_DATA_N_I,             // LP signals from Lane 0
    input                                       L1_LP_DATA_N_I,             // LP signals from Lane 1
    input                                       L2_LP_DATA_N_I,             // LP signals from Lane 2
    input                                       L3_LP_DATA_N_I,             // LP signals from Lane 3
    input                                       L4_LP_DATA_N_I,             // LP signals from Lane 4	
    input                                       L5_LP_DATA_N_I,             // LP signals from Lane 5
    input                                       L6_LP_DATA_N_I,             // LP signals from Lane 6
    input                                       L7_LP_DATA_N_I,	            // LP signals from Lane 7    				   
    input                                       L0_LP_DATA_I,               // LP signals from Lane 0
    input                                       L1_LP_DATA_I,               // LP signals from Lane 1
    input                                       L2_LP_DATA_I,               // LP signals from Lane 2
    input                                       L3_LP_DATA_I,               // LP signals from Lane 3
    input                                       L4_LP_DATA_I,               // LP signals from Lane 4
    input                                       L5_LP_DATA_I,               // LP signals from Lane 5
    input                                       L6_LP_DATA_I,               // LP signals from Lane 6
    input                                       L7_LP_DATA_I,               // LP signals from Lane 7
    input				                        CAM_PLL_LOCK_I,             // Camera PLL Lock status
    input				                        TRAINING_DONE_I,            // De skew signal
    
  // Output Ports
    output				                        FRAME_VALID_O,              // Frame Valid Output
    output				                        FRAME_START_O,              // Frame start pulse
    output                                      FRAME_END_O,

    output				                        LINE_VALID_O,               // Line Valid Output
    output                                      LINE_START_O,               // Line start pulse
    output                                      LINE_END_O,                 // Line end pulse
    output [g_NUM_OF_PIXELS*g_DATAWIDTH-1 : 0]  DATA_O,                     // Output Data VC0
    output [7:0]			                    VIRTUAL_CHANNEL_O,          // Virtual Channel Number (2-bits)
    output [7:0]			                    DATA_TYPE_O,                // MIPI Data Type
    output                                      ECC_ERROR_O,                // MIPI Packet Error Correction Code(ECC) status
    output                                      CRC_ERROR_O,                // MIPI Packet Error Correction Code(ECC) status
    output [15:0]			                    WORD_COUNT_O,               // Output Horizontal Resolution in bytes
    output                                      EBD_VALID_O,                // Embedded data Valid
    output                                      MIPI_INTERRUPT_O,           // MIPI Interrupt
// AXI 4 Lite Ports
    input  	                                    ACLK_I,                     // clock
    input  	                                    ARESETN_I,                  // This active-low reset    

  // AXI 4 Wrire Address Channel  
    input  	                                    AWVALID_I,                  // AXI4-Lite write address valid. This signal indicates that valid write address and control information are available.
    output  	                                AWREADY_O,                  // AXI4-Lite write address ready. This signal indicates that the target is ready to accept an address and associated control signals.
    input      [31:0]                           AWADDR_I,                   // AXI4-Lite write address.
   
  // AXI 4 write data channel
    input       [31:0]                          WDATA_I,                   // AXI4-Lite write data.
    input  	                                    WVALID_I,                  // AXI4-Lite write valid.
    output   	                                WREADY_O,                  // AXI4-Lite Write ready.
  
  // AXI 4 write response channel
    output     [1:0]                            BRESP_O,                   // AXI4-Lite write response.
    output  	                                BVALID_O,                  // AXI4-Lite write response valid.
    input  	                                    BREADY_I,                  // AXI4-Lite response ready.
  
  // AXI 4 read address channel
   input  [31:0]                                ARADDR_I,                  // AXI4-Lite read address. The read address gives the address of the first transfer in a read burst transaction.  
   input  	                                    ARVALID_I,                 // AXI4-Lite read address valid. This signal indicates that the channel is signaling valid read address and control information. 
   output    	                                ARREADY_O,                 // AXI4-Lite response ready. This signal indicates that the slave is ready to accept an address and associated control signals.
  
  // AXI 4 read data and response channel
   input  	                                    RREADY_I,                  // AXI4 Lite Read Ready I 
   output     [31:0]                            RDATA_O,                   // AXI4-Lite read data.
   output     [1:0]                             RRESP_O,                   // AXI4-Lite read response.
   output    	                                RVALID_O,                  // AXI4-Lite read valid. This signal indicates that the channel is signaling the required read data.

// AXI 4 Stream out ports
    output [g_NUM_OF_PIXELS*g_DATAWIDTH-1 : 0]  TDATA_O,                   // AXI Interface ports
    output [g_DATAWIDTH/8 - 1 : 0]	            TSTRB_O,
    output [g_DATAWIDTH/8 - 1 : 0]	            TKEEP_O,
    output				                        TVALID_O,
    output				                        TLAST_O,
    output [3 : 0]			                    TUSER_O 
  );

//-------------------------------------------------
// parameters  
//-------------------------------------------------
   localparam				       ST_SOT_IDLE   = 2'd0;
   localparam				       ST_SOT        = 2'd1;
   localparam				       ST_SOT_ERROR  = 2'd2;
   localparam				       ST_SOT_DETECT = 2'd3;


//`include "memory_map_mipi.v"
//localparam ADDR_DECODER_WIDTH = 8;
//localparam INTERRUPT_REG_WIDTH = 8;


//Read Only
localparam IP_VER = 32'h0;
//localparam IP_VER_WIDTH = 24;

//Read Only
localparam LANE_CONFIG = 32'h8;
//localparam LANE_CONFIG_WIDTH = 8;

//Read Only
localparam DATA_WIDTH = 32'hC;
//localparam DATA_WIDTH_WIDTH = 8;

//Read Only
localparam NO_OF_PIXELS = 32'h10;
//localparam NO_OF_PIXELS_WIDTH = 3;

//Read Only
localparam NO_OF_VC = 32'h14;
//localparam NO_OF_VC_WIDTH = 8;

//Read Only
localparam INPUT_DATA_INVERT = 32'h18;
//localparam INPUT_DATA_INVERT_WIDTH = 1;

//Read Only
localparam FIFO_SIZE = 32'h1C;
//localparam FIFO_SIZE_WIDTH = 4;

//Read Only
localparam FRAME_RESOLUTION = 32'h20;
//localparam FRAME_RESOLUTION_WIDTH = 32;

//Read Only
localparam MIPI_CLK_STATUS = 32'h30;
//localparam MIPI_CLK_STATUS_WIDTH = 1;

//Read Only
localparam MIPI_CAM_LANES_CONFIG = 32'h60;
//localparam MIPI_CAM_LANES_CONFIG_WIDTH = 4;

//Read Only
localparam MIPI_CAM_DATA_TYPE = 32'h5C;
//localparam MIPI_CAM_DATA_TYPE_WIDTH = 8;

//Read Only
localparam WORD_COUNT = 32'h58;
//localparam WORD_COUNT_WIDTH = 16;







//Read Write
localparam CTRL_REG = 32'h4;
//localparam CTRL_REG_WIDTH = 2;

//Read Write 
localparam GLBL_INT_EN = 32'h24;
//localparam GLBL_INT_EN_WIDTH = 1;

//Read Write 
localparam INT_STATUS = 32'h28;
//localparam INT_STATUS_WIDTH = 8;

//Read Write 
localparam INT_EN = 32'h2C;
//localparam INT_EN_WIDTH = 8;
//-------------------------------------------------
// Nets Declaration
//-------------------------------------------------
   wire 	                                mem_wr_valid_w;
   wire [31:0]                              mem_wr_addr_w;
   wire [31:0]                              mem_wr_data_w;
   wire [31:0]  	                        mem_rd_addr_w;
   wire [31:0]  	                        mem_rd_data_w;
   wire				                        glbl_int_en_w;
   wire [7:0]              int_status_clr_w;
   wire [31:0]                              IP_VERSION_w;    
   wire                                     mipi_en;
   wire                                     mipi_rstn;
   wire [7:0]                  int_en_w;
   wire [7:0]			                    LANE_CONFIG_w;   
	 wire [7:0]			                    DATAWIDTH_w;           
   wire [2:0]			                    NUM_OF_PIXELS_w;          
   wire				                        INP_DATA_INVERT_w;          
   wire [3:0]			                    FIFO_SIZE_w;               
   wire [31:0]			                    FRAME_RESL_w;               // Frame resolution [31:16]  - height, [15:0] - width 
   wire [7:0]           status_reg_w;
   wire                                     CAM_PLL_LOCK_w;       
   wire [7:0]			                    ISR_w;                      // Interrupt status register output
   wire					                    soft_reset_w;
   wire					                    reset_w;
   wire					                    sot_ready;
	 wire					                sot_done;
   wire					                    SOT_SIGNAL;
	 wire                                   L0_lp_data_stretch;
   wire [g_NUM_OF_PIXELS*g_DATAWIDTH-1 : 0] axi_data;
   wire					                    sof_axi;
   wire					                    frame_valid_axi;
   wire					                    line_valid_axi;
   wire [1:0]			                    VIRTUAL_CHANNEL_w;         // Virtual Channel Number (2-bits)

//-------------------------------------------------
// Regs Declaration
//-------------------------------------------------  
   reg					                  core_enable_r;
   reg					                  sot_error;
   reg					                  sot_r0_cclk;
   reg					                  sot_r0_pclk;
   reg					                  sot_r1_pclk;
   reg					                  sot_error_q;
	 reg [3:0]                      wait_cnt;
	 reg [15:0]                     L0_lp_data_shift;
   reg                            L0_lp_data_pclk1;
   reg                            L0_lp_data_pclk2;
   reg [1:0]				              sot_state;
   reg [7:0]				              r_isr; //Interrupt register to store corresponding interrupt
   reg                            GL_IPT_EN_reg;
   reg					                  r_int_dly1;
   reg					                  r_int_dly2;
   reg					                  r_int_dly3;
   reg					                  r_int_dly4;
   reg [3:0]			                MIPI_CAM_LANES_CONFIG_r;    // Camera configured Lanes

//Address values of the registers
//Address values of the registers






//-------------------------------------------------
// AXI 4 Lite Instantiation
//-------------------------------------------------
  axi4lite_adapter_mipi_csi_rx  AXI4_LITE_ADAPTER_MIPI
  (
    .aclk         ( ACLK_I         ),    
    .aresetn      ( ARESETN_I      ), 
    .awvalid      ( AWVALID_I      ), 
    .awready      ( AWREADY_O      ), 
    .awaddr       ( AWADDR_I       ),  
    .wdata        ( WDATA_I        ),   
    .wvalid       ( WVALID_I       ),  
    .wready       ( WREADY_O       ),  
    .bresp        ( BRESP_O        ),   
    .bvalid       ( BVALID_O       ),  
    .bready       ( BREADY_I       ),  
    .araddr       ( ARADDR_I       ),  
    .arvalid      ( ARVALID_I      ), 
    .arready      ( ARREADY_O      ), 
    .rready       ( RREADY_I       ),  
    .rdata        ( RDATA_O        ),   
    .rresp        ( RRESP_O        ),   
    .rvalid       ( RVALID_O       ),  
    .mem_wr_valid ( mem_wr_valid_w ),
    .mem_wr_addr  ( mem_wr_addr_w  ), 
    .mem_wr_data  ( mem_wr_data_w  ), 
    .mem_rd_addr  ( mem_rd_addr_w  ), 
    .mem_rd_data  ( mem_rd_data_w  )
  );     

//-------------------------------------------------
// AXI 4 Lite WRITE REG
//-------------------------------------------------
  write_reg_mipi_csi_rx #(
    .CTRL_REG      ( CTRL_REG      ),
    .GLBL_INT_EN   ( GLBL_INT_EN   ),
	.INT_STATUS    ( INT_STATUS    ),
    .INT_EN        ( INT_EN        )
	//.g_CORE_EN_DIS ( g_CORE_EN_DIS )

	)WRITE_REG_MIPI_CSI2_RX
  (
    .aclk           ( ACLK_I              ),
    .aresetn        ( ARESETN_I           ),
    .mem_wr_valid   ( mem_wr_valid_w      ),
    .mem_wr_addr    ( mem_wr_addr_w       ),
    .mem_wr_data    ( mem_wr_data_w       ),
    .ctrl_reg       ( {mipi_rstn,mipi_en} ),
    .glbl_int_en    ( glbl_int_en_w       ),
    .int_en         ( int_en_w            ),
    .int_status_clr ( int_status_clr_w    )
  );



read_reg_mipi_csi_rx #(
.IP_VER                ( IP_VER                ),	
.CTRL_REG              ( CTRL_REG              ),
.LANE_CONFIG           ( LANE_CONFIG           ),
.DATA_WIDTH            ( DATA_WIDTH            ),
.NO_OF_PIXELS          ( NO_OF_PIXELS          ),
.NO_OF_VC              ( NO_OF_VC              ),
.INPUT_DATA_INVERT     ( INPUT_DATA_INVERT     ),
.FIFO_SIZE             ( FIFO_SIZE             ),
.FRAME_RESOLUTION      ( FRAME_RESOLUTION      ),
.GLBL_INT_EN           ( GLBL_INT_EN           ),
.INT_STATUS            ( INT_STATUS            ),
.INT_EN                ( INT_EN                ),
.MIPI_CLK_STATUS       ( MIPI_CLK_STATUS       ),
.WORD_COUNT            ( WORD_COUNT            ),
.MIPI_CAM_DATA_TYPE    ( MIPI_CAM_DATA_TYPE    ),
.MIPI_CAM_LANES_CONFIG ( MIPI_CAM_LANES_CONFIG )

) READ_REG_MIPI_CSI2_RX
(
  .aclk                  ( ACLK_I                  ),
  .aresetn               ( ARESETN_I               ),
	.mem_rd_addr           ( mem_rd_addr_w           ),
  .mem_rd_data           ( mem_rd_data_w           ),
	.ip_ver                ( IP_VERSION_w            ),
  .ctrl_reg              ( {{1'b0},mipi_en}        ),
  .lane_config           ( LANE_CONFIG_w           ),
  .data_width            ( DATAWIDTH_w             ),
  .no_of_pixels          ( NUM_OF_PIXELS_w         ),
  .no_of_vc              ( VIRTUAL_CHANNEL_O       ),
  .input_data_invert     ( INP_DATA_INVERT_w       ),
  .fifo_size             ( FIFO_SIZE_w             ),
  .frame_resolution      ( FRAME_RESL_w            ),
  .glbl_int_en           ( glbl_int_en_w           ),
  .int_status            ( status_reg_w            ),
  .int_en                ( int_en_w                ),
  .mipi_clk_status       ( CAM_PLL_LOCK_w          ),
  .mipi_cam_lanes_config ( MIPI_CAM_LANES_CONFIG_r ),
  .mipi_cam_data_type    ( DATA_TYPE_O             ),
  .word_count            ( WORD_COUNT_O            )
);

interrupt_controller_mipi_csi_rx INTERRUPT_CONTROLLER_MIPI 
(
   .rstn_i               ( ARESETN_I                  ),
   .sys_clk_i            ( ACLK_I                     ),
   .interrupt_event_i    ( ISR_w                      ),
   .interrupt_en_i       ( int_en_w                   ),
   .interrupt_clear_i    ( int_status_clr_w           ),
   .global_interrupt_en_i( (glbl_int_en_w && mipi_en) ),
   .status_reg_o         ( status_reg_w               ),
   .interrupt_o          ( MIPI_INTERRUPT_O           ),
   .interrupt_overflow_o ()
);

`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="author-a", author_info="author-a-details"
`pragma protect encrypt_agent="encryptP1735.pl", encrypt_agent_info="Synplify encryption scripts"

`pragma protect key_keyowner="Synplicity", key_keyname="SYNP05_001", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_block
GYRUuJIG3IHx61F/vIHuNuuGKluyKZ8/4eop9h06s+OHzChr9u0NGaFAu51EE3VOsgfTvfUx+rpP
Qyz70mCWlByl5+4PkrmJa0L30YMm0dt1ADB1NzTEqQacsDbyvi33PEbttzhsAmKYHjAh92z3qDu/
n4H+fC0RmpLpcG6E4ffTNwGdC2RCy/DpAeRqrUzEFuey5C+jTql5txsiJnLO/KXPRtt7ZUBK2VgN
gM23IH4rpmlyrPMPBup3PMvwtBRQSfzaitqofwOgmu2aEf/fCmG/txSCzbSeIxVmyYgC7PR32DHc
8LuSRw8CcWM9bpVsL9L8RZCaptiOfFQtiRST+A==

`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_block
crYgiFcXWtheV5SIZyIhPjuyIWvVb8J/1ga5GgJwWLvOShQRVehL+URlZIIGEObC5SAzsiM/Ntr/
FY2GStiKjxJlIPloyzfucVNHui9TksPHIPYkrl1q0CRLR85RMIa7JOlPLB03tAyBKtvO2rSBdvfE
IB5AYPDsD3FYdsMSEX4=

`pragma protect key_keyowner="Microsemi Corporation", key_keyname="MSC-IP-KEY-RSA", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=960)
`pragma protect key_block
XIpATPiOjWHXgxm7lKnCNp2SA/5x2Dr6IRZ+qzDAC6YKJImoe+RhwB9xjIGRzDg8Iol1gRreScEr
/1jbHWlPfDsH3c2TRFkoR4gkEmu3O6sL3qN2dYSOTr/2lVg64ZU70bngaSnyMo1PR9quPWOvM8gq
2NK0uASdAW4y9GnViP3JG0ohB9EBkzXGvhvYOc+Dg6R/GyFvOyvsdQ5pIgzhU7uFx+3oarZ0FmYY
7K5FtY+BKcOgnhmxbeWy9F7HkstYBFz/8DjYmVAASVvpXn1sjYG2ecpaWQ4oVb3QE1f4/GpeC/98
yDbygHULx46O4HBHDA4IJSsfcUJRn7URd+pPzVwEp9U3pm10FA+bpnuQF25uudSQTl45YknE34hB
11WOVNaFnSc5xXR90TMtQc7qM8Umx8LAcAQM7/R7Bn5wELc88ypIJ3P6hLgxgGTYQaXsBTX+5tdu
X9CVNrwfauCo/i1Y4EB3DK8CNeoA18DU88d+I2JzwztsRUzzHrx7/SniQoQSb/xwGZ21Gsfdc3bg
Cgrg/SfDAvxoO3CjfCKBv162XbgUIhbjfZhVff6CYjvMCWBNrThwqLmyWGZ6JIqIgbZUgJxnpnLF
jHQPCxoOKFM3qpK9Dr5ROLRveZRAW4aPheOwOh2e6ZwI6Q0CZJjwRftIPjqvZUd3Mond8x6vhNlH
jq1DlA9xhX5srRzSXlRamwaeB3RyOU3rz4N4HHKI556Chbsup7j7MegnLBfx/NFxeOLo67u+jKE8
tRjrKS05ZvOTekglEwtfkeXVAViCgc+FRO0ubufmtTFqVmI78QEB7iLiDhBMbmN4SOsgMtfu0MD2
HC1zQkxu6yB07Skt3Vje1FQwpBo3rBx6ASLO+kUfaDlaORya5F//yYLqmqNHhkEh/L3Qr6Iaw46C
TrdWfv0ohWo5PbAo7mlROqV/yXcIXe/Zq5isZ55aiWfVg++ECDy4FKCCj9Ay85YjXPAmUgkK9xkm
gIXANXu6KBA6wQsiHF6VQP1TAU3YCzyjEzCWVPhSXk3JnN3va4iZXUuxEqDCBjn0Oh319QjG5hkX
FHUCR5tCdzWq47HEVB6kKXsOOn3Ss0I1IQoEBTWAOCNIjuzJggbNibBjNCxF740zyo9DT2wZ0VCG
/wiYb1/tyLatbTuXSnxF/PSdLmshcx5a4PzES8AJGU2y6zloUShcgc+iyoutPqFiYHQ+Pyt1vpBO
GEDx9sgcorHRENv4IyOTW4CyGyfZnYkTgkoCse4wYvjXNaQnPuWNLSMuVIUNf8rt

`pragma protect data_keyowner="ip-vendor-a", data_keyname="fpga-ip", data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=305632)
`pragma protect data_block
iBB63lDE2DGMlfVQYs6WtrvlPByK0gBKm4pvN07LgoUV80q0RwSoIPX8VSbOH8msgwUDWJtrWn80
Z8FEQzAeOAnbSzItigOMLM1Xtyyiw+gRmMyhxbK4+7hIMGJ48uQfGwJrdB0zMk/R/+k8Xiha3KkX
uUyQA6GqtAFov9XSjL+HO2vmneP6+eGwnmJnEFjj3WXClVS1zbsIMcuYMQeJUCa6Zqr8vgfFBk1+
ePd1zp3WmDW5M7mtfe+vaxwij/H0AY1FKzdWhH0hj1as/9nTW6ZVmaEQS0bEuO3O/IPG3gKQmK1l
TI25kIvW3DT5duxCh/KPKJ9A/77gVZ5yEQZIY+D5DPzzwEXX3vIXQ+R8v5D3Z3/NRiWU6lmshcuE
r420qM+a1oK/m4XrMZCXwyWmGIkER2ptujxM2dagVyPfAcyXoKQYnPlxNS8Hq3XoE/RnzGOpT8DL
fVKFa28/O3DcBSMqC8cIGUWu202lYgdIhFqgufn8fc1/3crzyWSogEoUU3BGTQEPQn/IeJl7vR61
J86OGk2c1fYr+0ZXz/nWnR0j+4vRA9vwE8idJTm5LAuGv0EJETaOW7VRXXKL26vdwPoHt7NFeX3r
DZhIMe30p7ZbbIqOggBLSSIqyQh2P9LACTxYK3UFzEc37sicm07LCqzZ7yyCavwNom4/uNFcLvZb
fZ3pkc7V2qNVzUYnV3JTacvDRwCbcdxuBEV3Rs9DMKPNUNbCwrmhGrK+NpBQcpWhZ9YODnRiK2us
9YwpHQQbXwjeg10VCRq7u5yeFAR0x+Ik8YH42yATphZNGHw1XSuwK0M7HZB+/hLFZAWW+K7VjJGo
k8iSoqUyj7GKeIY4ZVL1Gh1DQxLGBj2idfMsbtMtZvHWs0EcFWDk7zQyXdc8eSR4S6IR/TNurbhS
pV7uEHu/iWYMu6FNFtN2SHUdBp7gP0pAXHoHPVoB25+I2FreWb3gVD4ZTkfGRlqFT6k63KwwmEXE
TJVHtbdMz25q9vI5S+Hw1xQQF/UoCaiiNRrSQeAPws6VFiJkerUzYFKOZv1sOUGrmNSOwz5QHzeY
j7nXyyg2KaypUlARkQfRYoLv9gG3CtwW/MTZ8Wcyg51/Gu4MoRhSdjKXbIo6hyqhzsCtfy5bCdFK
zIzx7TX3dR4b76fIVr7vxX6lzR05irIcEnbBDoXTzewzoh1Iqxi9TAMudFWdksR82p+tlhMzAJ76
LLMnaAp+va07tPJsbbUA21p+3tuVadXSVi1rh0Q393mHudVbwQK7+kFge8iiKC+ir44bUNng1XDF
tN2Vqg91fXxB5V/GaBZiLAsaX22npFa5P+8EVXvctxWfYhk5lWdQ5y+ouW/CXy/TUddNxzyPKCQB
KLw0iL/rxHTXT+SsP+mfCEGjwa3TIbRc6K5L5Pn3eYiyvu9qMq/qE9E2CgXJbQREhNNRHjEDIE4b
hl6XJ6ouEC58V3gZvIiebtnJMwYMhh6Qph4yug9nMd0D40FXqClVsgW1G0EdHnR0XvUI4uuwh5/0
VUubsiHlFtBtJrWbinjbb1DwTxZsG/MCovxDSMNLKt/Q1KL4pdr++j0PjPvgzimS4q7keKY8Ms8Z
NoF+1yLw+mRoCk4p7rszvUFolcsQVCUvZdMMPN3DGmlyxNNHyVkSB1UTDvASBEd7bMZVQmMdFX/B
K/+1EAeqk0Hn9xU80vs8u4ItECZZpsfIr/pnnQtwtAhMlymqtDa2De39b8pAd2sic/BtuXji0fBx
otfs4+Dn5+j/oFJc1a7TxAdsG7/1MFOK3CI87SA+DEXhFvHf6itsh42sp0rwApttC1/gEXDGOwKZ
PLAcL0BARuOorCkS0vlD6Q6A/9++jX8je9TYMm5RUAd8A7fOSbo8mymgfyKI9ZOsd2glzUfr8nv+
hGNTqTGiIV8KHcQUwPsGe3u05axWRPLyd3OIXubpdOLI0gArNMMP7ejhXcApDjNMLqsHQb3/Fp9e
BWFkyaoF+eOROT5YRArGssVaSnFp+DlWiyFFb68sg7LKuaRdviMehXc1+Gm1Ld/5uaIVlgJ/UVqH
ALfiGhiRKqm/erGEhbRN4wGBuc0yjakWEfJ6ubTa52lAyarbFdUIYjr1nThAWWT781OB36HsHNpf
BciSA+dhy3PEFDJ/dSWg/UmVz94SWWPpAtKEci5xRHtODkr+wcb+OIP4X59sZf0P9XBWc5+oHrM6
m4HLGw//JTWTsKVk6R68EZoTFyZt9tAMiVC63XRp4xao5mS1y1sXP2lF+g/ILUL/iafwMsCwu1A/
SKi+6/3IkFwkm3K3VVeoM+oxxXb+sePpTJg5xJGz+5JimLH1Rkn/bt81ZUsZN/mgBd+f/wfvI1Xb
UlKPDTu+WnK1uP0bCSXatZ+3+NzxQ+wTzEgeMqK6LoGcaaxzznnlbf2eUpRM+f50h8NK0FPgdrD1
UnE9K86WMroW5UvF61ZbRItNPWyDKBOooBFWi9/cxDOxrSuPievvIBr8ajVKOlfnrMXphWP40wKv
/uw29RgzMYSTjNlconmPpeEVzoyUI1eZznXh41autTKD9IdgYTfWU1nNeOWkhJZc5v/U3AVAV//J
rcWhaUBdOMDV4ptvr+24bTjcvw056HUZLg1eIordrIXSWby7E9aI/xrZBmfFPkFokUUBKunyQkdp
EslQn0tCGQo6YLdyjZknml113/rFmmZsBKLk7i9h1QC90wWoO2lMmFjPJFQP4+i4oVAQbvEPVgoO
hQU8DgLCYN5mA0uan7MVa8cQY0YvDcnmYHzef264PA/ng1wL/v7UWfNQUb7DpO3cfe+ykn66mAif
LReacS8nLudWBI4YzEE6QXYB2pQVB/y4PPxofn4pF7Lhr1W1DQlIZSntTbbSK6664optf4kYouEe
lDaxY07d5ffyWchUOH4C7NGXQMLSuOUJhBZXbpetZRvlxLNmZwD+sI4EpnasXGDxp+lOc0YwKUma
HrNVeHo8OWZwlSY6hehfZIsFQx0c+KJHwOkPEqYUwmHfwY2t0imL/6YFjybLUzGC2s6FF7LgOruq
WRqUbBPh1RTmds5Z6m8J8vpZRZ9Z+78hHmw1IJROU8LYf15q9Y0nPg6CacJcY/+103U/MB3qJJdb
oLKeDaMm7YZm5zCeBoPhMR5AcTnkrr1LYA0UUrNve+Kitc6eWVJNzDoqlve4r6UqFK70O7vGUrPj
8wIdWaz+NdW5usZCpRuWDXPpJRQv992CnWa5Tprq//HA8F6EbLwmXhTVG9m7L0tT6D/5DSWFnZli
bW9iv9sEclaS6DSKpK7ntG6xp72lDJOx8gF3pcvxjdgmYwB9z1AW1/FM84ARWcgp4c91/hv3JH61
Jls6CyMluMVn1oahk2ETu37N3pGtwf8LTOP2ULlCyu6az6nJSdWs2Vn2l3CPr5g8Y7Fhjz3cvrNU
Z+gbNnU4295Ax5+sKuCmO91wH5lhrqoD1HLubSOLVXBwpom8ZNLizGg/YKkZ8i/ba1qiGPujLibG
DSSAi946fn2vaQSDPrBgEd5LnW9w7X6MYPnUVT12Zd8AH6TW0MIXg4QA3nLOqGuVCiE6eVl+IU57
InYJid1Tcirlf5Dv157dyQYe1YYDQdKFXLHYXvAGEgRnL4p+gokdiD9wqATXEKKIEC76XBOPrEcO
lWIBz5xpNBIG8tPVDA9gn0A4NQmyWwbsW0UCVKvmJLDZoDyhAKAu384zH+MrkXKQdT6Nxp6QpuoQ
WZiH1wV2SuemylXPbb4VrVjUf3OtDYnTxad69gBpTxx+cPMcFELTqMA/tw6WBrgcwq+3HS3SGMSJ
+tsxmbX9TP25DwuJiUGTjU5sVzTEOmmWKiu1CxG60DiYUNAsE6U8JMa3ESKX1r6RbgARI2JWeUCl
sGbxwUdvGJs9Yjs2ItIYJQtK/uzSF4uIUsH3w9IOMaxgEo8Pw8w7jfuHH6hxKSXHGLCYgJXSM51W
mrr41CkWfDWyLj0l20b9fzxlU9dSj99H0TGvbt7+lgdXj0iZi0rhBNuYnkiUb08dJKoRro72/FM7
cqe5wNkTb30MB4HoGQdnsbK0SUI7527JqHh+j1D2wAeQW+F4vgsidp891UF5sJM660NwCaZbhdiK
19iWDj4utmg6DrnFETILgn54eCDNA9UpJHE2J/VBLeqhvxKC58UzeA9Fq+lneh1deHTDaERsSmkH
Y7qiWCzcki3J3lZ11AbV3UqudB/z0CEjlXkLL4+uIPqtzmhx+XOnaqsHnVSvqayzgJRfdTuKaOTc
f7dhCpUzMJvUw3ZfVKvSewUeycqMUNU9OwVPVDor2UhEE1v0OWyyvTQ0Mj382WK7Ja0Efv+Hhwxb
9cwNadzE9EPkamsyqSXCKi8vFwDUj+ZHibJ92qDrIj+6fDY/jM2kKyXCRtdimFBgmiF9wFXQggPU
xuoVPJ0XIjmgtoJLL7xaHw/sLDiUqefQDP3Z685PPTK1URRwPhjq95Mg4d6XqHDYMyP2fXeP8k8y
h5D2hM6kvprz7GGjy2dk6vI8fOSbLutdGdStObbie8b2GRNYDW1hckO5qAMtMfHZkxpS253vygUk
+Oe71nNhTiP3/m/U0u+QnnkNrcKbi+eYMgB4KcL0NXVZcJZoIBS2RX2VbpsKGdedpZhvOZt+zVjS
ZP4ZCFYjn4astLXIfyG7h8RWGO9rQiCSz3J7XjHH8gElUmPxuZhcJrrcrWinPvH9Mqjmq3qD5SL6
fUR8vvpeQl3vQbXVUF7SBESlr2S+A37QnE/WLP4exmk1xOCdAc9GfXu23HQwqU8hUPXpciDxk8iq
C0CPLQ4+TLdCL4XsbNkUD0Z5EHCuLCubhfqABvLrfx+EJKgn5gfe0K+QgjDHd44I6nCCfWCsYuCk
Z+DmfMcGUiS9AGvWpae/EBKnvphp2zOvSoWTl6C+sGtQjwWpRESJVVzRNbHipD6xXzkzixZ/0mQ4
Gk5nge1y43WrueyMdsHR9VYpitbzhfy6x3lXgB+kKZpukOMJo92b1EV0FtAEniiqlbOraCfyB8uw
XmpsymzK2qZ313Z+BSrLQYeTeTfqCNrNe9atu2quTJNEBOzbwvkjfjLgK3uUj7WVW/97vB8u+JKN
C3ZGEWbuekIBI0LGOwsUQC6ksCtKZaTU1uPnm3LIEs1G0HZJ2DRXq4F9w6XqU3c29shQ5lLxTyIy
dktKL1piIQCH6AHgmyU94FHekCX+LZ/EuKUzqT/lCRj2oqZI7nXIw5kNoRT711FMyFulGn10yc8d
fNJsjmjU4/pk2c1jnUJXK0igilfAH+/7tjrQK8DyE+xlmB/pVRlOpbshN03jUpA0FxIE/Nn9nd5F
+7bym3OMQ00TmVA1tYWMYKM1K+f0AmL6G+J0R0GUm5xFxvTMKRXyEr22ze3lVpOGBWCCAzaif2Zi
ARhyTMweDwBV3PEn1wZrPyB/059TI6jsicIyQ7fRcLQjRYW4V05/NyTWdYt2VsW6hubZMy9wB2Mc
nUCm2AC/pM65oGcRqDNRZCKgNV/Qk+LQYO5VE6xVVpLVRhyk5qC76+GkYNnrqgqfQyR3ogEuEGYy
Ymt54IQWJ3S/QEP3D41j8JVcxwwnTswvu8vuaXF/3+bXkIyNMybs8InZPoeXvLuU74mSrXC2mwLz
VvAxm39XkomtNmg60dfw6Y1NfaGFF43F0ev7J769cSwa5qfn0i/+314wfHTC7vbyWGUtz4VQArcf
y1G4cGsIuNwCJ7zrXgmo/yYknq/pOrPTD5QPGdfrrQj5N69xY1BTh+fVAw0VmgEPrLPRYDfzSU7L
TxOFpuS3wjixkrqycNfOd/yHXR5EoxyxbzDTU5aOjbpddqAVAOM41KNSItfrC3za1OR5sgEHFhr0
8vRGw3TZ14EepoZJfvqYnUn78suHSKZt1ZIdwn0X2+okVzGGamhgBe3I1TXK0TjmxuEXf/oR2DKl
bVHt9mzswVq54xbQEyXegdP9sfDR8kmBcgwQaB7vSNr2WiuFCtUb4lWVd3HaQ5xIoWQv5Cyj8PrT
fjsaNImo5M5b2sXlX0s5KsW9ac6G3zHXZFgccRKzLQn04QjGRereS9UHeEn9BCT7Zuab2l4sFhL9
EkV7C7uU3T5xycnxW2aaodPXpYgcAYsLkr4iEv08/q8xSxHW3HqtI8Blxk5qa/q7aakpHGFBFmDg
tTUxxJsByGBuWnBL3mv8Ci2mA4wI38mspg9c1neMpUyE8BZJQsJe+rY7202Jc8JQ9tfuPJDEDEe7
lLNMSm19kyrXwpTb1suuOUa3HTAQ/giKbYftlZXrwI4EC1x9PWYzjZhvKg+0d4uBCPif654QtF/h
5CzJiJZPSxies8+GgWal/7LXjClAAaMftoPcMNPZ1pgnhZ3Ls92lkuNfRct6TtErllJh9ykhtT8x
c7/aPdvS6pss+26kAOmnbfWRRfX5Fdwptu1SO0RvyanX9E9vkg4ZN7Kmll78ld0OEaWjqQGwfaQw
6cCwqy0w1Dk/SkwabKut3TNwcWdHb3u499hUZ4j/IElRjmmKKKtNxmwkQtAfHFCywAu0jZVY0CGM
NHNO8PwCcT81gku0DcfZG2K5UzKPLrtDltjD5quajxv8a1Vhim5QJRo+BQIthBy5ucpI2MiCfuff
kEoRXIYZYCMp1sbJpRbiNb4PkIjH7wTQlmzYyBCJ+BFPwqWI4KqdwwRMHnz1yWPE3HEC+6M+A9Lo
uL2MTgUAy4huC4n3pkyTk7bsdxkU8NBdnh39TNkbi9l1zyMlBpqHPi6E7KJWMIzVGp/2RQHqhyC8
D9b9TnnRCE6WLNedQj8OjsnXxM3tucY/tvSvWG9OrlB/uiNQyBIiKyrNfN08grATXIuDQTEbddyv
RXApDf2TURUa+fOI8FJPMyHtKpcATVkjDT6NyAyFbC5C/inLTvRaVip1/gJ60PcAL5iRry+du/BT
2J1gzt9R/7thDFVwII5gsf/1Uif8XesvUjWjR4bAZhLUVYgFHAsJbDURqNNLD19c4fqmf6DGqKNe
4O4su6RQowVI0818aX8EFQOxebyC4M9GQRX8omvbLMinjDPOFJAMSUbFQFhCuACZwV1wMUp60K1m
nZ/3LfFR1SpsL3zqPPiNzMz2b5pVliC87/hU6FwV8khSZyi4xQ46xL9auI/qE8zatRduzx7gbems
GRenIH6viBTidmoiZcR4UfTNJ89SHjY6rvDY7bStdxaIVoa0Ck9vV8pK+dffFh5Sf3j8fO1N8blR
0L1PBNhf/hO1IZ3r2QUvXOirQlz2osh2bo4Rz6q1lRi6VUw7DM0BMk/U6IujeiajxN5C7o/Qa5IY
6eJddSGyGdgFGbxi9wmsBZ1b0wCO5RpaMlSXytZr5N+RJqrU6dMF/rBdnQsE9gvGcPS9MtcvZbPu
e4ynlTgJNU+4cRRlLvtMeGI1D3DvYOmboB/4bDsQAw6PupgC3/BkesX5Et/nU5g0WB+JtOu2CCdZ
8s55WylX7gDhfm/Mxq+pT9ihhnVB975hKlAlCKtkwmQgw4f1Dbn3ry9sUqRDzVYk3+tIvWbGzumD
SdzvQA2w80K7rAAwl5gjQqoL6pcNdERihiIH7EUtA7LiDECWUtM/ds4Lw6721chcmbf9tKgZei0U
G0BrBC96JgnUjCFilb0m2XzDFbgM9R49Lo/81byXpyZs5cfAU9e7RoXIywzqLG9cp8d1ECVv7ChZ
jc0bhOcp4LeiqkBfCmRxrohsCCYnOCtXFL+3tJmabNewHx3FMHcerKcNyV9Hfeao3czjJQqoiABc
Lf1MFi1OBjghcJsZvNr8e7ylGQ14whidvSkqrWXQTW8yyBrPZgYfYmsX4yrVv0IVaVx0o3bf3cUA
cMZtKKjM+tIeKvGLgO3A3wXTJuxMD8fufPm0ghL4dmq5zJqlNny1f6+3eLLCjF0brxJonjjH4Tyr
UBMmLO9XGNzCpYtCTvFZvDRJgbgLEPFUGLc1K1iXGiN4d2lPQN7sy5VAcDV9bGcG2WPgaa1+M4m7
hkKLnW+i6zNlcuBnnyIgSHWkN/oRh77tTwbgAoUbEiMUPrEV0pK+M7vHQOcxn5++SkRENBGRqaOF
hUGpSASrEXDsk38s/6dNlIRuCKaII+8/P3tIl4LIw9ZflHeJCdrTIFRRyC8RkYPKLq+SfXl/VmMP
HKLIr9d0cr1L5q7pfykJAiQtt2elSuqQ/lI29M08bjgYidatSkH1b2rDsVnF7xYerH/2+yWVsWa9
kCYop5bMY7otBcsoUb1UGjKuguLwJntLVlFfeqrhnWqv8DtpQggU5ruUW3kiYsFfuovyR0s3JxtP
RD9dZOe8hbc+vJWKjSfNUssZzvQg2kGts6q1ROWg8rdog4ahLGF+qB1qXVYONAYCgjGMgZPqMcq0
athu2NxJDijmztQ9CVLPnD93/sgbD3N7UUSmjRo6BLuGE7WbRflwsW9+xtyvZZS57UPToGz+n2jW
71AOSffio68jia8ApVgsLBWAt/IolUAYD+2/hPzlWc/Qo+u0xx1unWsPhOmwCQrbjn2P/5wG+ul+
KtG+TxSJvz0ezm20aa1m8M+NQrzJki2pZVXy0sSrB9SO1SUvY6CmkccMrKwVIpTWgsTQ75FZvzV5
JtPbygP3W1h4Q09D+4AfDEAp7FFy7P1ehz4uMHdutsLtyUPdpLqUk5mnU74a1iyJjTAINy9miTnA
vc8EilEBXlA4R9fyvz/lzJI3zItgebRj8jOkRHfqBgJN9hpvR9dui0vzODncv3yby8UAWvtbU/Z0
yTjlM8MPZU1daJKHM81VHGCdaK0maa8ZEcab3nCZNaGup5TtJXuXU21bWw4sMIr1CZvuEzn1+lQq
/GHb7l83A/uD8d+86ddMTo7aaS8GKrjeK13OiwBnNei3iWicKqgTf70c6dzEFlZIBb5mZlsmmQJB
bZdngNVYH+2pzcu9EfhN1HtVxMiEd75ItamcDM4/XfFnBz7ZZDbZdVtusx03Qu81oO7IpS5mJ6XB
Y4NBR3rsIBrCXIf1ROzFVXvxNXb2TN1OwVsgpXrWvOuil+awYkNzgF+eJJwrLOVuNWJG8BRyVpjY
bO8UtJ3FhPTZ8dUPf5y9wCjj6QEs40JOuEfjaCcN7k/qB7j8zcD7KL9AZtQOqPiemUPemqpssC1E
QfarzcDu9sdHpmA0X+h7qVnAdzTkLY7Xo8bhNUuNizRj4EdvI8tlJox8zLncqgattK+D8aEQAkbZ
tRkcoBzBdV4JK0f66xT8Wj/UprnAlVLmZADEoEOGz7GY011DlxRveWN8zfBeq53HX/qP08RcnqdQ
UunRNU5TkG2duCdYw2/ToP8Ww9AKL6imw2pIe2d2cFn4ZEWktEg6WxdGpo3KiJMceZdsX5Nhp/3I
gOA/Ni/jQ1lyFDW7isY/AfVtjUlUNUsd/erE0PD+8OmrmMSGMKmfHT8zdCqGZXTybLmiIrz673eL
lYhUCxxPWuSh1E2rSCfoo8rKYdIBzld2YKeQqmTF0HapomojUBwVIJqw/OoB2SyKKsZkoIkVYts+
OgV6PuWrqnE0+tdvtkh+W9geEOxfVizAUDflMHvCZplOERg/88+9V+qgqAYUpdARZIzMAJfiaA+z
8jGDM69kyDP8AYLnZ1U2e/Jr47Q4lHeQQ8TzUc8Fu8TbSsWeHPcENAmj1qmF/ruOX5mdvsCaJ4tW
gaRjh9yD4QCX1R3QpaurAFRIY8dCHIhKwD5HPSwwl70ow9EmIq2J9M+R/YAmcEkbc5VwdE3DGtNi
t6EhEoMm8cf2BZH5HLBPj0CHWIxBecA5zsaYLorxTOqP6VRLUTzP5aQOiex9uLzdKCdu/7Rxc2fl
xzfElLUzzfgQV8h8G61sRNR/4Q9f80ctYzqAQCjRVrSvjSVtLd8pBytF+lSQWv/IVdmBCgBbyvwm
oq4Y0WoxQdX/olbbrGmcWRCw/aFSz6YkhE8sAh38LYZGdyjX7e3rCxbNP+JoGNSM3aZHPL9K3ady
vie7rI4QEcWeyve/6xYiB1UH1qOULtTuzg8AqLYavzxKD6lSa1+MiFvNW3Gg0W3ZhkbcYH0j+P//
3HlDbQdZR3aqJcbkRJmjhYl9PkU777k+zqGmY29jdUEMpynuBEp0+jz48u/0hZV7La65dvGASZFZ
wSV7rMf8EvXX3z74M7cfesvumlSZLmAYqYx6RxtM7Daeibb52O93Q1fPl9+cnc5T/Dazih4axl5V
f5WC0gWcVZxrQJWgcw4F6axrLo1Y3HQS8+vUiqlExHyHgT5uZgTLRqHqZi0A68qufdT/47rWPsAF
QfJpR+J0U+gDRQEWUr0oigO3R2azT4aOdnvL8R58+GuaLXgegDKQmBo9vHrXtRKfRn/2+TgY7PZ+
lw/k/PDbYJJsYRbHmc385dfWlEJj1MQ0umH7QmRadC3CpYU9TGSWC7c8scz3prLbtJlhKrr9aXME
Jy25Xkc2KskBmc06CdqDsblc6gLd96GwaG8Pf+8+orp1Gr3dW157XQ0v1fwjTNz76FxMM5BQhE1h
U6Of8Z01ScST8IjChywZ0m+MkBuEwDkMjdgTokBRTJjHap6jE1mp0dke33yb4LPdIbXoEJz0jGRL
EzoK/s7dk6HL0ZL/Cxc7jzBjyhFx4tlcR1Q8fVBMWbzhQgn+dvQETgNmRo2jvqPDfO+Bx8WTel8n
C74zuNWe5MP+444pUzMNvvG/LkiMH9fk9iO8DDy74CjREQd3MY5DQBuCZzHF2P8lh1YAuL1cpGlc
9blJt7aMBlznw+EQrF2CvQFOn4zb790LCazBjPdGKv3a52PU8UrESLxl+176iUMvG2X2c2k69/Hp
ta+iHRzAlOxH098eZbh4z3m4bpmmJHh1aqIr0TT0egpYqdNJ0VRWU1lVfzQL909FdqDvF4cd+1KH
+mmMt2+9qUpBR66Rv5NSD4vtQ07AHxsh3qejhIVh/3FzB5lIR6bXfKBKmm2Ip84YKp7CmuJDBHeu
BrJLxVexQgGlZIwQC1HIO1EGHdpKS7dztGub9blf/drEiIhoSnqW7TpG+z3Jbm6nFP2vYdH7KFJi
lJE7Y635oomDXbvzvjKiRiLRkcUMkvbqXF5WNZoSqtkYWK1twwUIr26nvF1IY1Akdk30sjQfyWVi
jctRYWdHsz6nl2T1TrrCYgM/KmX6jK4+HqEQhCbpTanKO9ury5nJby8pauP79EXIUIHaiHz7dThP
lFci5qTJD+I25QiXTYaKXLYS7f1pP11/oIv9+eNztdvXcR8ZY92xAyhRGGmxbinMiViovjd6/50n
33AnBBFAguMaq9BZDa5zgad038OKqgxhpHMyxUvixuMRgCF2DIF50rSSOUdS+GApIdfIYjr0N1w2
GtL+l1fuVQ85o7lUa45Wiwf3sHRbT7ere01MDs3geJJU1xj+ItK1i2dW+mlgssVjFPVRqp+kr0Fj
mz3cgfZIgacsh9ytPEv9nDx0CBXGuYWAnBPj4ZQav+SwPxjWSh7N2c/isE9HnCeteKJrwFitRRdL
GCtwedwiUFAi8SbXzrrmZWbl2CcrKztZLMiN+9La8p/TB+3xW7EFonp6KNQygSWC2F8Pot/4aa78
nOqPevvTEiXfDg+3wkUwfMxULnFxl8JKFgYJ8Ij4tOIb0SbGA6rKrOi0SAS/tfkqMrFVvtI1An/w
aGNLRVdImE74LcivI+npWzr53Orxm/9jipzM64p4OUYGeU/cjik59LWoRHqha4OZKtrHJ5j2UJ3/
uNgh9tB8LaDXEfesyGmM9WGPbzQxi7QKSorZc6a/d8CNw8oyH9fb81QHOO7bx5c8flJmng/zGidH
EfHRhDWcUPO9+FvLirsYubjEuqC2EQAoXhG+DKy08XVCqdjvI3yCEkKD3ZfwKg2f95WMC3jGzwE4
dLYgq2R+M70dLtaKD/k3EjSDMG88QigbyA6Cm55quirUcLY24TsjXme6x/jfYY4jP3F4LAYUBLkU
zo3VaA7KmriBLMxY6pCZaQE6vAWM3fr63konw4HK2UENsVgVazyqPyscBzThGt0pAEcAM92Ywe3F
7AzM256ASUe51K1rzN1IC3gWNd8lAzOEnPXz7FkZRKILmR1T96jaHBSWQLtPWY7f2hUWmkH6euNm
cYuP+mrKYIklF1AzKYF/V+UGbtWF1DdtrtLwAizMoa7/kP0Yn98UzkbqNC8Fme7lyb66V1EfW+/s
58ry8CwZ5MSiuwUPzUMjTOpfyrTbG5TF0ASrlkVxB22vUbb2yaI1UIflVDaWi42m7xL3P3l19XAD
AnL3R6dl7+ofrDIC8EpC84nGBsMoyJnqaGsPKcukXEB29FgUqjcR1MHwMWVD9qe17E9K1e00M4kk
1J85I2TwiVL05AvjozBnifbw+rdgGGsHWd9Vp2LdcufRj2ujsRrTbAhJxQuCR/g37pQgn3GJ/j4v
BChvqHr7tW2PDBJuy8MyXPK+pxXXcBntegUoQM7DfeYnghXyGl1X+khPS/v0oqzestYRU4UToiS0
FPj1sQbQUvH7eWjiDVytfR4yeSNdzQ8d5TVrawriGpAby6yzxnF8qI2AAHiCMC1K5nj1YmnDZDBE
eRXhA8gWqfJ4XUjO//9W5IPfZjBksL67ISZDhrnTf8epXMc9sN+w8+KpRuXsEmndRbWK+OXFii5N
jnG8Bgw/UHtZgwG/lA4TZrXg9Jy6IVLb1VvoUK1gq3VQdbQThYHXsmp86mbxDMsYgZbC3qY+Iqe3
s8LvdJGHhKzM7g4dgXLmScmgGSQ50/hTiBsbb/y8ceBF3jObW/WqI5aYBLVzQBqEhYV5n3k0oMUS
BGI1qi8XwtqFL5z9cKiXyGX75PwUBd2qGVI7or8M4thqInwbHJ17N7Tml/GAv84vv/5kXgnBPNpH
98zrgI1P+LMfOu9EzxCZzR2+Znfqa1SvxHyot7x90Xq1AEXXXrMaXJ1Gb+MP0wp6I8WxI6SvjgGJ
GelbXXmEiUUOLBMxvL0aIrWLQRbV83xV3q9XDSEUzeyQ370xQpXG0xZ3yBmoeJzEMLqwwT9UTBoE
yljQCojIn3/lwRCv+tiVz3Mu9mb4FQUr5bIUb585JTkUd3eZWnCnFfsqaJQurrv2kSz5rYTwSu8Y
PTDI32tJdEJUfDO7O4Gn+RADj12Cipo68N5srvZMcqEhTBNO73A2OxR9mVwSVFrAYkG8igQtyHO+
ASLbNuOTn4SIqa8z7xLziDEMBjb88Qtn1uzQSXPU0enhN4V/8nWOdzMfPjYOCQh2BGGV87heDTYV
NHtJJfkcriEZcn1iQvzcynEj7DnI7MgSPp18ZjV5GYDIXoLOyhJSLmSGeGuOmJNah0W4xdnlilzc
iuOwMSYPoXUqkrOQBtdO3kwNiCgqRop1BZtAzCcL+PXEseQQiInkosOTddlHPF5/ikO8W+YfaUTR
TvPKkWpzDfU6FvLVLx/JYsEvZfM5XgIbhxwiGFAFXLm9uOorvK7MYZy4rsDdpXTjfDp2Ynvbl+Kt
DpKPHNXLobDmAN8vMH5wEsSxpWltMA8m2U4Nd2TBSghOEf8/yXhGDsj6z5zJCK3uf0gEawxMJoCH
E5WOKQ4pwgCsP3GVAG3S4SBBXDplbIYkNByYPTesOI3IwD5wp1syti9R+snSGB+PZPPNCGbYkVAY
4f583Hz1HgTNaK16JHVuM0gOf7gCuCfvwTwubuVKduuEMXx9LdXZ3Dbg9kRWq7TYtjmjpuKGAEKr
NH7dqLPEU7wv0uRuFEyjt47QJ+dlcNiBfKHl7ZNfsluzfrRrZCnfcfq7r6UAKdx/l3Ak+0V1uzDX
qQZBknZyKBjNLzj2AfoAdt49Fg5NzkmVpb32yuQwaZAiRw0CKYz4tc2oqWN+X36vE5zkmnf378OL
NiZVj8SH8+0Yygi29Ap1ReqUil07pvKS0H5RhGulmmlzUP/CNecEkN/b5KhvIgnS2bNhmrOn/HwQ
YlyMqzbNAEdTDZ9vBnlMsib/5EXjCinEorHvB7SV3pEnCkf9Ads56QMAbfGRSl2dRd7YPmaU1sSn
doKxaNN0hTfPOVjPple0vG1TwxFvhFRLmG4EWWfTKYvV0GWHktiMdrrAMSpRY1hIy5Af67mPCOo6
Gp6kPASlUBZVtE2hzQPXeTI901fPl26otP1EG6QY3ElLbtWUvppbvSRA9LNwoT6SzNBFW7hc9DND
Gb5jYjr06ZkyZl8NILR3RFL7RCA2n5K6ckt3syCqxBof6Dk5VH38AsETMmUKDIp0fnKdb8V7MGJs
pU5T7w/w5ialyjival4+xxzr9G4KQbkmid81gwAZ7tJaQdsbM6ywed6IHDHPl8SNOTb0jsquCxpM
Hw3lZKPmO8DkK3pc+r1bX9iWss17SMdDTNJKFUANsU8Pf9euDJB31Rf3a24goDbW3k9/iFFaAHse
dBKBLYFXQ/0dJPuNuEgD2kDveb5IgNfSSTs2WZnjP33r2EoC95LGvy9Mp4c4WjvMwvkV3hycI1fw
Arn6bNNhHB+xRCc4THlrB3irH25kuBSj4M3AFkDrNp4yrQZiOVoZQS2IQgVHfjnA2GLlaRAknJrz
9YXy6NWbnGyimXt7ZyGxZJEjN8T7t6q1qsi8y6oRrDxnjLE7dNBpldqvjbLXLWySNwavwn5Mjr6f
CxBm8tNomxvthQudMTMMTDKYPgIzysgQHxm/JshCHM3Lan9l8V1/CVnSj6ugQ8ONyUTSFN2zdWkG
Y/iN+iJFf9dygdU76uFWFpXdqp6bE1dJWwKMfDaSlhrv+d2z6KvqeBIAreKmBvgUtYEdbWc8BXqj
IfH0nrM7cSvI19f2WLJR/ylIzT8lVDivdQrNEZLrkUNMBtyjzDc8dGhMg544rwzEzhiwIU+ywHN/
ZU9Zny/fGNwrAZsw34qHxXbz0TU3LGZqbecQZpI1QNDjvx4VtxDO8G3VZfcvU6raT2iR1PFXPhvB
4NgCMIoAgh+v0BRox0Ao+77V/lmWVKW+InAF6NYkf2ENqLCcSt7s3U3NiW2T32I/EYMiHxSJ2KG3
IUbYRMWPuiOQC6V4l6t1XcExtFrPM3yuRhMHkAkH56TaXulALx1lGSbQ6zzO9Y99oPrgjwG3jY7K
zpHOEphmuGd9m/y4tenPBGr05jzFuvO1LGcQd2ly9YK304Rv4T+QZ+qFbSKsTHfqV6LYtIUl3VFn
ylupQZeXJPi39qimg3qwEWtHiBZpxOB7kVc/nIHncIiSfuNgCv+cDpXPtTduDsxBAPWtdS325dUy
LelhQAWgmEOLMNLHRMDlccg2xgDs12DB7x3MmpZdqDo2Q/NgmMNVSiJF/IwdLaITe7WcRODNIAVv
icCON7M3Hia6mULGpR5rAX44rnwW0pIpNt/xjvrWuPFiANdiBD4mMJFyvxJvAAHVoAwmny94xdiK
e85HhM/gb+xceAOsk8qdAWqAXanYkxC8+ZWjwemR9lB4CQxtl8P54DRoJqrhC/PDLcxJaqtEulp9
jjxspIAN9+dhAGiLv3W+TkNB+V7MB3vWHM/k0MHv/6pjeEypw2pGUPeVR4nA0VSZWV+HuWP5j6zn
OBlsQwtyYPW88UT6tfWuigToLi2hc5D7AYimVTIW367XHfKjZMrDdxLaUJRpGqbORpHPNWjkYokw
HQVpg6fX8k5JCxggn6NZCiSGhUkICHiCGEXvgcfF0ZxTpsVBboMMsWqGyPEffcHVapnj2XtHPWOj
dYP95nsy+3V6NC3fH79BusHLOd5mVroF6iGkGtkAtwgSfw3wOG/WQ9dYBvyZ5aTrMPB0sE8a3LOB
+SsnirFI9rYM3oxktWn5tItdUqRi2KrieGPwZ4MnWDTDjEK5oGSZzrBxq2fdBbxOpZddfinTpZjQ
c9uUuoPL+TL7OffiXu5cPXdfK0tjiXw5XnaoPgyt7dGWV1LrsNM8OJTw0s+vy8vr//odvFn8B8Iy
XZm+P9Losouo3eOPYDxJmgC+ig2OJn+j5kwtfjCXXVNU9NsZr7f4b0tlM+GKXZr4WenF69kkGqdO
PWgbgrUeczTbhKtaorp9yHLdXQ87mXxMrgVFTrbaOdRYi/cnPMtXfeHmIZcpW54GQks9rrBztiU3
0kki9qpkf5Uc0cBlaEv7M1fuhFT70KLotr8VDkuAB9m4hROcD9DsNfyFJrJSVKzF8WnfHCOeMZuC
25BrfoIgLyulMnrBOlwaoibE/V1HfbD8QDEZeq/6mf09XV6W7NNygn/Hb4kKs9rg1yGfQrdVBm3d
/Jwd+eGdci0CdIEe5VzPwwXH7aLiM+AhFzPmqUZSUjMFPR53L+FIz8uahvmAKZwGz2Tkb6LNw1Z8
Z1u0ItLeh+vhtZBP5adZSkraZDS28sb4xwg5H+utFpsVUXcvmDzn68u07aGqjzSauo+744Ev6oxv
BPplmWxCis91QFyaWopYE5F7P5Hq4rVANH5WTMAJe0l0V5q/jz6LmF1VSQ1fk4P6SMy+YiWi0Gb0
9cecHmFPevhcl2p79P3gTASANcmETFcbPMgQoEhAfl7hs8K2clTGel+1HKzSZ8aciqyeh4ioWMqL
WUd/jkWvH2+XNmq8iBpSUWeGpnO+RVSCkJtWAiI5snJtXpJ4/FHcrD+5gzqs/tGzSC91Ej2fNN+4
HKGgsxDrQJ3fgOSyVuuOwavudu/JrWpK3WakOiKUoKbAFSrc9Y3x2od95V/OCgNYXXYuBAJfF0yz
/6yhCWcOFKN9wTvKcXxisHgK3cjt2IlZN6iC8bTonPOnI4bHMpECJ/ybAdNVsI8jqWR7UqSJjXr+
j5hgNtZ4tUaQXQESPEKqithSvRBjsxH7k4vYXpz4LTc1CHDLCcd6SgzRdy6/G5ry3FMwrmXwKPaj
zWUWL1grbJW+F3FbdXCg+vW8313PiRPTUe88HzeAgf6n/XRdkzpGF5A0ubjyYNOg42huzg/fE9z9
71yOjI+RslOcERIQ8qtCw7oQW5V6nHCQb3ko1UKOYYPLUwjce8XGBCHfuRwbfAy2kuOp+npHrWfO
YLhpuLhZCj79Gb4HsOT2FNVr2VhL5H+EPrwbzmJL0sQwoFpVzgRA39A8IYSs/y3SUbAj/oLim3x9
YPgzkKtLrGedXqxtUr5UStmXyoFwerjAZo8cfStuohBsNfXwr6ybyPiBNlvJBeQzLAOLAJdRz76D
ytk2cf7GSjbimh2iVnV9+KBvC+JP/D2oT8yvbZGbkks9TlqSjCTgPlmEbpOFj9+gxP2QJZR20zMs
EsetYIteFqY54BCEPwhyLHuD4IidgDsZiOM186jXm4o3kLoNllZ+fojTkO9483+poe+KbgHCffyR
W75rR4Is+WfFdQBkUMoJabdrLgYLL56FrTK01NZBk8ZkRf1z0NVjtswrJQf5hp6Me2pU+1qCeUTR
3MmR5yUwZbAhNQ9e/trUr8LeZC4MLRuWlPpl9TPceYWBb6qdHfmJk8U4eTJsYhVlCMnGiNqNEACY
w3qnsrp4gzO+WUsIEGlxDdzFoGG5TZROZEryLsuXmcWbbtLnIuO8wgxHJym3pdJjwc6HJ+3VokDB
d4nM4WV3N+wADbt0dj+D9TZhir3RBlMBRJ3um4F3655Aanygi8eHSaWfHi+K/5kPHGyu/B/DiLDJ
2+dV7vvdWmI6FzWtMhcxTBJusumiOBtUDjnjdMlnrtotN2sdUEssov0SLz0sUMQOiWN8nyml4wk2
u8T1uQqS9UWNMmCv6+66mgbv9IUCn5nBftFXJoq9CsYplm77yZQlkE6u/8AaSp3/6gwQsMxcBaD3
fzb5NgUgzq8DYrUqZZ/YWbuRc96FUoQiUAMmXVX9V5ZXDz7wBAgPJz+T7WdKUhsOW+GpIkGejGYR
fnKmiFIXkiIKnfzQvbojZYYq0dHQuC9C3scYpVqxDD8hCDqjfhtuiSu36iLXo18d6ghhHgC6cSAF
0oxKQaa19ApbB0WOZRAYWppTNdG7H1UiM4qd3unDGEyZN2BtuHMy8FUzPpWlfOMJNF8DCZKwbUw2
EKCllQXCz7LBLVSc4PqT32BDNl7nh3Kr2CQ4gPLOEwxDboa8YzHdOnUT5K9X0QoiGfhe5onJiZ1i
lhr+pp3crHoqr9P7raF6ksG+gsLE9X8Z6/c3ONY/0APeF1QJPXm5ST5MrxaDhaonVLvhQzsCkyUb
eomYWRZXzd/S/itqpLcHNWC442NudFHMCov3kI68b1Ik0JFVvDd7Mn61fmmtMa4Y1F7GFlhg+cOj
q2jTT1WNT4+qVJ2QdupFKIS43UYKXU6kPqpdzYaq1x3ca2yftWqRl4Dt6WmbbfvPkZUyRW8CF1Oh
rWUPyaZMzWTYlmSCkpXPOuJMaEnDoMUo8YdBRw6PiP2/gKGe3xrZOEgFTRylwZ1LjuD9UQVQ16Hs
pJik38djbykXzvG6k8/QqOjdQun6fm7oQTYazq0WSP8kGPuHWBaOinRN/elPc7gjlEQeejUiQIod
W0qao8uslQ+W4dy2Nti3zr2hAWU1WB7HO3ZPFKDZjN7sokeFetyvqs7B2Q1BhNwkVB0aPa+b5kFA
MZhERwscZnCNTgYniXfT9Wtedv8Q89JrqfRhxauREa3iSBtF3mLVjV4A+Nu40iv5Xm3xFIDkIeIU
muYQmYBzVYu/BVWXcW1SR3cWVbQOrijdEvFihJglOGbT5bugsitWWcfkKU8LM4E0h3mbTzQybMFV
lnBHETtSE26tOtpVkbcHvUh+zJfE+8CKBCleiFNL4l0WckBcQ6dBS/jsMr5ixcSoDS10wFYLbzte
SYZGuXqtoTphVA4Ei3hu8NmEipChbaAlRVhsr5l1xRU8YKgGlHzfWIm0/ufG2+VSVabGyf7sIp9+
UsNUVHfSQ7uueizErEkuHCPtW595BGRou1zQsyKLgXnX/jsYE+jyeEAUtx3aGenZuLET/G4k0N92
IWn4vTSWfQ+Yn4r14IkazA0btTDWpY7QKu3FHgthZMA5NK1YWlYJZBkObvD1Mb2HK3qTHmEfa/2T
atjnc9p61IxSb2QkNvuo557cZoslhvL9vZmmQWTkf+qYdAb0szvi0vlZC4RS6TMW6WknJJ7Mz+0i
zfZWtGD+EVevQIVAlK+26yjZZ2/jgLcoFROCs6UgPbYC+YC0CWFJeeQiIrgI3offzb4l8pUVE4Oy
R6uKuXN0fGim3XfZ2ircKYcsqYz0CMQLxb8bCQbx8cTnuhIjK507+J3lEWUt7rMobY9XnHriZdLs
UheWYWVFkirqcNRDtLVYPOhqtJIbVpz8v/jYtjn0UZIKNhfOSBdehlfgbjS3GGI6qsGNcOPa5ZcK
djB67srbSAcsIQQmkl5m3/7QLv5YB6d72BvDYZ9XOFE+18oWlgt3X5eE+Cqtz61lAo7f6KqoRjd4
0j78umszL4E/5gnX0YvLRGG67eh4GxP0P4sdl0LMbwbPFJm0aXDdtDvmZHcyeeq7TK3PRloqYYHH
AUE/v+dA2M7CaW+0GGul0Qnw3jqJp9n1+v88xhT545FYgciokq3vR9YodkbUye1CN2/5NQxurb+c
KQteB+EkUS79tkKLro1rkZc1D4WA+93gIB07tPO3lN5KOebR+73wbveAZUBbMpAopDKMw+GPFMex
7cFzOI1hV+T7TCmGudI7065zx6WL+TDahlaJh90tAk6BdntmmDLu/dIaf4BkeZ5RQMZJEvzwSRp5
GYhbAgFohGg8buQaXToK2Wgv7UMrSRPHUCxk5D5/SXcj42xsICV3jH5E0KgdXbyQxOUbtqc0N2r8
4zKldQVLNcCv/PJWoG+B/crTSKry4RtauzbiGyFouZqS8i9SaHUX0pZVjSg/FwOohf6iG6xA7rtI
unkzgmweuiL/DG3PLeE+B4a2CfT11shcljVq5vYmFSpztPyd9MG+VbeOB72pZSeWbU7PNdMb88en
pId2Z9opl9BMquJx/0ZIDb5DDw3UrLzTi0XukjoV2s/0iMRKsiWi5TrP5+v1Qc3zE5QaMkBUzdas
Wo3fbGXrudGQ97cWJzgTQTqnm5ajz5jbr75GUT14/K3ihyzOlza/4GhNOc7H8l7nt6R6OyH0Ifw1
oR92Wb1m2yrWGO5/To4sXRHR5/juhgCEUPLr+HYMPyIEd5TmoCXCkt0eO1zC4MTvbnFK9tyFdWGD
g5TMsa04egGwUrWlDGZY+3O8p67AaxNjPUC2/nYobQ0iTvxd2Eqf1nkshaCxy9DtrveARXYtTYGT
REKZv0zM43XdV2oAqdhKMv1Gr+qvPe5MeuZ5RxjS39jmRoSP4FyT/ZnCRzG9HOA0d8/Pl7vqiR55
hu0tPQKmpdGLwJXC2gsmqcz1BH9dIXFXzNSMD938H30ZAMTtA/udZ9QaXp1bDmk9Z1mkpXmJgEey
eUwTIBslt7cDaijme2bqRJVOf6D26XCBdkbEWmw/CDxLCoQ1YX0XXAGDDhFF3ZlGnDdVd6+Pu1DT
FddVgwhjfH7QxiYRRpTBhL2q/o+JCxplu83n10f/6vRGYWyQgUIMqwS1qpkmwTNXIRNYw4iPkVsM
eO0flEj/hr4DgivZktI0VBSQwZjbkm1g+MIxMdbbLLMMrHGeggapnJVUzAFCvJ4q+N8CIUCkqwff
ANQl99ncFEmOuzWxkV0yNwLl649fCkUsaant+WdZAo8QKxpZK5PksQO/gG4gO+OTDJV42qDJpuOM
5aP7BpT7NBHVU4Yx2sbqMr7jCusHyUMMO4YeMIwp3O5V1zsbNiBKYkF7ddhSnJNedzCd/MYs/ppI
DI8ez/PiZ6rMpoVqVqGXS356rQbgSLMx56Hic/WiWAnH+RWJgTyin5+WBm9LhlOWkyvso0Nc29PH
nquoj1l14oIsHWGXNb30qF0v27J4/ELGsZSUiWrr41fxNEOXvQlTPdcjrjAelAEfpJd3IZbtyOhZ
kCKtc4GjN3jYbp3es9r4O9n2lTY4p+Mx1OhdqeYmC8cXT2T47TLVxUAKAtNCKURe+yRe6JQhdqvQ
I60AOQn+ApQWckGCzrOyN57wN8gXuLR8Yan+HKo0TJeGU557pW85K2UkBwUJ3TH2fLitOal/k+bG
xFtE6uUDSl7B5Q22tFMt83W+ALrMCK91Onj0a15hrsSmUHckBkV8dlnLj8JiuWlnSvVLJ0Z4GIOK
6YCmXa9qXBHIxtvNcHISAw49QLrgvJU7cWCl3S4ToxuYa2F/IgNNxz/Xkb/9TiFQnXvKDyrthNtl
bEz0zQjUzvgov+gmC42ZzH1ogxoC6sGUqMDRFJiuiV0EquNa2JvcTDEf5LwZmnxQUQrPhgXNMtRv
aop5kt5BIs0TLuzNobggbzc1jDN1gxpBEskNPq6p3Az13ILQERiS0YPJXwVC7jzQKtdXBFJcexYP
r7zAaWzsG+ZCoXlCbqHPe4uqqr0hLWUfHIr3OF9zlPxik6q9JJwrtDLHyG1+hhnmcdNyxe+Ez3VA
q2XFraCXSp2kettLBhiFVQ3HhUU9rPHEhhZxiDQ2BKqxuRq1g3lmlDeB11f5h0+K4a41hwgonbJD
IEqdd+e12TfQWouD17iOiKsiYMMy8E6DO+s7Gh6uDmItNajfj81PQh7LFuaszxPw5cffA4la9Pzf
nD4cUF6V7P2+/953VEJpHHn0gmTV1EKSav2KMrIxhh7SblQOCLHwjgIqI9cDQFwzb/TiBrgHRvrH
7IVGrmd9SBMRmCrZgsu3+B7Gigp4NXXGNxPS74fcU0gIfbXqd0uZ5DJUCfRTooMCkP2J9s7Uvri0
w1HBtuvqcymrkix/pj31BkAVCIWdD59eMCE/1acQMT9cPZmZbIsHcWQptjHL5v5fQlncmyqPdN5H
XBzqUsZj//fVJiwa4n9lmvHsFHI71VBZdF6cRscxYsQFtStNRuzJImcvbNGjL6evIyFfU83CqNIO
ExDB3+FWWufNGqRbcj2yySbCdGICDxV1os+WfW/IMShntO6XLeRmCPPnfvF8+3qxhKPFCvAr5INb
0GCgHz9Zbq9N2RzDMiPV16xyK9u2R2yerF6zuMg9MDabRaoW8bIayPFROXEH8QdNeuXFaB5dD+4C
8xCgj+Ibv8XZvBxdGs3iR9Sv0ZmqTXUNnH98yOGhV8hL2NU3/dQ7dpAeOtIMEVjDpdMxd93HPqvS
nzM29i1a6kpGQ6sj77AiYQ8xsXPv2EwqZ2SdDHl0ymSBfL4QS4CQWZwn8KDLOx5gZFe0d5miufgS
PDRIqkw/YVrveBp4/QDsLULOxmR1kzHhTjNOvC8V/cm+6YHni5Y1MNAfiND7MbrDw4bbylmIrSjH
gkwBNpfekF4fCBFQtt9WTZdLYS66k2lJnfk2f7WhVrD9Jr5im36qmsyr6OItwgy1Ou03yqH4NrC0
dPjKHvfA+Zg/c8AXOy8UokWTxnr98PWvG0/Dn4kabDKn+fm72XM36kOafxddzd4qEqxsZtWYy6kJ
ngHaqw7b5eAx3lUvDGNGJCRQ6jqh2O+BRVKTmHkohrVrPK856xSD4x5Jt71oELrKHaO+oF0Kh6lr
htH6LQM0LmuV19OoUVWBfAZKWc3HSrNYorExjuy0+NjY6v4VQ/iiUuZEnDnE7XnYgTl5bGad1Jbf
7j54kjo9bEcHOsrQf5dvY/K+cFm4utHKFSuhbMyOdCB1mnemGoT5dpLHElG0UO9o3iq6GziXTAGi
oZ1Hkq260vnRmPYMERGX7o78uu1w2N964Hiuc7TxJFttLBBwdvjc9ciuP1aJ6wYYeAy7TmwTr1SF
E+GrsDw423f5YAL1CyWMyTpF5xLx+oIyprKSOStLWbTRMgY/jy7LhrRYehhm0gYQlYFJRUGbnSFe
i7+TclCZV6wQD1yFEAQOadxp8yqRad6bDINvlCeIdFn1Dd2CBnkWbSUbINvQto5FvxzR0YDchsnJ
RaOiEBrQq0e2/7zXdye7vEe5/8/89UQ/UEdBR9Jyq3SB5SlxKE0hv/9jcavUAZh6DM4GjG2DSPgN
qKxOp1MbGX/lT9RpgpFuaAZjHUaz5SUWK4mnHdk94Fl6x1FmsNBSbwrL+VbaSfTWu7e3tEfHwlBp
U4Fk8VKGCWhWNlUzOFWhg4RkoO0km+RCHyFWO2c4YbnfL3+kh54fuYfbhPnCokSPx2PPIsDT+8Ne
7QsLWe7Xg4VBk975EnJBzPi1R+hh2xCo3Jw0gjwhjWUsc6kE5xVlFwhbiLrcyeBK+kVautIGfpnb
mn9djGbbfqgkpaBWen0M8yrWAh5Z0r8fuq4iiV4jqkmyRqMYpHvwopo+IpAUmlR+vk1sOezbtaQh
RU7jRYz41c/3E1o905bsVTHohoeNdfp/178BDtoBkV8sOt73x41YLQwhX64nbZMps7m7wfi97eYX
8wPCQeSYjMDBOJ4oJvdbTnD2UNrtyoNIRmI+5d8sB69t5LUQaJWtYTzvgl/Z1vdWLdQ8BT96LWCq
iAbualquPGKxVppXCCPSsYvY9elnUEqlkhDGse40pUDnSTgZo3ftCOFU2H2th051KQ4Hn4WKYnV6
11jfNYzsTbHw41JjDJxTXuvbRIILBoBO5q1/w4jRYLKP5VTkewmkhd1uEfHkg6a9fFtiF5sj7bRb
lq5WhHTJImJAEZYhSk5S/cPY7REJ+E4Abs/AdrNe+wYWaVroSWCwX0tyMeElaqyRVERMZNOpvhg5
QbYFTlackn3FY43SsHRBvNxak7aeHleTn256yE2IKiclpCuNaVI6xxZteMRitKSG5aElkI2JOW3a
IfcEqqG8JSf9Go1q2e3bzOwUTVesvL524dGUmSuBMX2XgEseZkM/m42CqKYG3pr30q93OaE4SaSq
K7udNxhH4wUD/yqtJ+sCyu/BqxZZ4+X9aRxCy4NGXu7cqJH0Knq3qBf9T+Leu39RllXKYSZFPerM
CJWbKHSerYckxWucpyFbVX6ZgxXRnW7nM/45nReu6mXT69xbMftvKUcPthAYoTc10kJa3yLNsqvg
84MAf1Ih2bi+frbPDWyzmX2MxuNfVsf+0UwBAnEt57oNLQD4mZ+uMxwIOqWKr5GFjfMBN66ZWZ1J
RaH7z5nmfk0eY48bAb74Raq9Vp93BvqXl7n4T3+9ap7GMdOS0988E4PHzNFkbg/uh6NIphHJ4uT2
AJrYdePGOkkRF+DW015X37cWhGytOWHIOnjOg1yUtMLhVaqgePQ/Ys1uIHE7W0iprLHfqUDa5erD
wa62Qr0Jtx9+iqKgMO3RNf/5NKNSKsrmdikZ40n/e/+i8RbJuDid+muQho3nk5tQuDHeHfWkzopW
/ZBLqiAbWm5yVZK2yvfOt+vc7JZkTsUTY5o36851wz7X7hIgadjFsS+mbzdz98cNyRS+q26vJAm5
7uWSAzcf7FS2pQYllcNOSCzJw+jyvObZ39dp4aOG0IDF1iAKeDIKpjgS2CZkhcILGYT24qeZ/CPm
oBkMjzzPrh+ZchMa5Yhx+bY6OO85FqWuzom4krNe1XEEfTtr5ZhakmJf9NclmlOyZr6Sx9hRZNLg
WBkBDLo4dguq03O+Mc22XhEoAhtuDlLAo8oJVLf0aGYP3DnJ++DWNSG3WPsOqkrNpG3RdY5Jtdgw
ONW3581lIEsYf6I2UTo243dAZvupS+TAcx55fW/9ULnLfJmtZc+EFzEAKQ7lhxcrGUzWyBlDpRH9
TYMutEOiZQe9Zd6XQgIyKAbvhbGf/PaF98rvnYK5MLeHOj/KxS3XJeZAEsU7ZOKrd2ycHj9QIoay
LhsATw/Z4qeL4jYMQ33jWo5bj134JmEzeJ68+LQFYXojtVuzSlsBA7X2WVgJvj1vpqaj2RvpvBtE
hj+EKvzvp/PtKSA8LfleZOKPSayUE3k26uV1W1MDWbFWyQaY7RgZEFnpnf/PPfGKjxT4ciMS2gmD
wGXWjxLDkgu1XS616d5aSMkXogjGauddErAdqrk+WEW4kE+/O+wskoFML9h6uDGVr+F3VBo4hOTo
95lScGd9bqOEX+bTZUvnnlP1YvqIZGbbpQZ/+ZQ7cg8xMSC+h9D+gnJCZ9ZEch8LuxW9Rp7snf5s
KQCe9t4ZSiJUT35ll0Hsy0C/3i8y9vCclOFxpoFMAbygQmaDM7KL0fsIlpAqYTXUbtYQHuqsooM+
8pLZWakaS36qBrPXsz3JE0WIWAMAgkfnoYA4l5hndw2kZUmtajeuCJOHxTpyF7Am/sTMoqKdeTiA
0/RZdDuyrLbJOO/WEkGFuoJHlcLvx8S0d0l7dA2Fdcp3bVtYmxud34ImFqRZY4XCtW4A15f8meB1
B3bkygZsMIna0ZjkvzD0aVq9JD1eUxcc0uyWGIEurSKhFDjoFbmz7qSDkt0OeaeFp8/Ah15JRk7h
tbBt8onhvkbjLsA8BnSZUjGHkYtgVLbjVuCVicOxPrKqqinaP6JsqXPO0bZJiKm5SO3kl7DnvAB9
GrdGAGSVpxxNytaaiqByIeUpFa+pPDblhuDXb6gXUQP38aIXRx9CHmm39iIvBVx6MNHZPn2ast5D
GFsYled3fCspRuZwsWNZygzYVXt/EkOzYzRc9G72hRQPtY1fQf3zcn90X05cmG6J8HmxYozggQj+
qiWdyTpROm+YkcDmxm/PJ/W3HxtBJoKDBXcg0Ta2hDsES+QX8B6HlI+eRT5lGnmodv6+pm4/6+qW
ERf1oK2/55h3b390A5z2rLBojAHTWK+cd5THXkCSlVOyq8moX0XnAv9ws02+LnOuE6uODyLF0kZU
lkD2IVQGecjmolg/nDCC3H5WnMcA0jeai+pSFUcMJyA8u2UttOgAAmGp+xUQooImniWtOQin+c6u
FHQ/U0SWt/1lq2saSIDJDoBT6Ad9/YcSwIg/fQbS1CBVe7MdDahtSQiGF4c02L8R+gQJ7dXqfA6I
l80spp59ShaytMQpIOovjemJzbFC+lDkV9oKak1F+b8BmghUoM0KjAKnmBhGnlUOo0oRlznZhufx
dUr4JsryVdkKb+W56wog6Ptdtn0TDMDQ3xjBPF/iIQZ6uoZVx5HarrYRfNTCMR/nziO6X6u9Pyje
SG2h4IeInC3ZUjplAd8hibluDwvVtG5tUvrN9WOpKc8PQ1GB16BiCsDf2LcKoJs2flH7JLP2xKKc
bnrcw4bUBFf1zgpU+fKi62wqTng7eCDB/HCiNHoGyUOHdeVNBE9BnzkQxg3uVvknHHu6/YqwwP8s
yW0UbtixYaQ6YC3BoPzlJR+GWME34vBwcri+B1xqCqWui+0UzEvXlB6auFVIl+1+pY2zGfSa6g26
RMBJ8Z5YfIMobeZ1Z6I8YIfJlQxJIjE4qz0fazJodyRNiBvCjCLEQI7e2XbzIK7ngQJKEF1eBTez
zT4VHVsH4wXSvWkSDMhng3GeXS/b3xVr2FTo4Ri5crOCo5sVUxKoiuis172zm5IoJcYg+q5EOKqa
wHH8uPYVgeBSOpRFIRcxtbdcrXE8FcsahG0GGKbuQkWJeLoZ98jgQlkcgAyfTVRSHKOuYGjMWBvi
aM6JB4SflX0mZ0L+tO1jWvrXNMcfGoPPOwOE2s/oKqKRVT3YXu8337QiKJUALcZqVvoPKyF0Nzsu
qiykeNiMF435oA7/SCLI9bwkzy2Ksys1gbMyAa0Vasl6vJg557XFXAqdL2bkil6wYceUddSvq25K
OIrpEyHynBUHVsHbirELKKiF5lz2MNn3XLF5Fuaq4Z1HrgLucljRGrdu6E50F5GsxWLKPPOejXGF
9qqcy9c8MFm4TvZjtkiWfDVxdLMLTNp3ns5dYA4hw62yzrgBM68i5ZtI6aKOkpLnEWXwE6Ij1qmb
F8XAdsh5l6x9GQDdfx3cd2sGL4pCQe0VS7ZNS3aYm3+M5T1EwTsZjgWPicJ+vAnU0OubGd9QmhgH
6GhTIyswBgXeoDC6pVfgmY3aUPC4kUIAiUBTh1hty/YEUndhY5jxzzBK3PEy2ELTN+SUbd5q+Xrp
Xi0nAemXfvFZspibGenPPxJq4jZoLoTvJIEh7+y6mq2tZUDskojsZKh+b3HE6YaoY4c32ZP/rUYU
Js3gMHRi+iOltDHoCuJYP+p8chn3akpEI3RoMtXeXi0AMzxSMjwlEGGs1JwvIXgAXK0l7XiQTp8H
FosAa848dnw6wQqxuPq1KP4tR+gM9mJ1sVmdi16ho0aWdnFoSRDo83g9mHuBpLWKQXoKPOOwMfsA
1QBdAqCts8RcAgdJFVXBgrjWr7foXAexFM0JYOxRBrIWfS2VW4rwYoGrqu+Wd92X+oQyNnOzSXuV
0TZFjsPbFEu60lV6tom8D3p9crgrW7V6XVG/pJm3IEEYsLUQoGbIKn8wR0tqSG1w5B6twVw41fut
HJOBX/ubqivuFS3zvl6mxyXmr6EGzkSWkokvnvbWjXn1M5ebdEYsjgpTEyeo4GpL0HcUD2B6AmtJ
piEGR9dHdX6slKqboxYQEN4xB+q9cawewM8nSAIAwdeJSkI0L1kWHjCDVEsUhKncl4ZVDf48/KHf
YNb7jqgrSAo9Hld6ECecLxXRQHu9r9zTDDRq1pTf782kKj/3+kvi0VX20tSoiE+Fg/Lrxm/PIO1M
jxYmWA7aYqCKKFTr0mwOCFjt7+WxXWPhBf5KII1nAC2BVXcW53v49HGSe7KRL/Qm3NpXAVnluJYu
dhQrMNJeU+RIDCxT9qckt+uxDKYC76Mo5WMAys9bGlglwH2d9tGaRyZXWRayDblgP/enYqhUN3qc
cyLy9Kz8g5bHZXLq+RsaKcwEjj34ho+RJpsXyFsaIVd88tK5AmqdZCSIr65trZYgqUxih55CAAXn
nUN2tD1GU/7A6LiSwGmbTFdXv6U5Z71LiqXnzaZdJGwKFGfbLITXZNbBzVHuIj1qKFghZnaDdtsz
CJCBk232N/tIRopnC2s/IE+2YMxe08PUcMQG16zaBHpBferCUvFGHJwIWOYx61fIrjByRPvH/R5k
IkdHCAUQosoqU3esHA3pXO7E80Uro1+HfvwXw7k06UTQEpXnRskGYNIfl3XY/9JHiAUeYte8L5EL
nQvx6wktVWcc9WmEjsQ2lUiwzF5ttOJF1FNMBZnmgJXPXTdVBoI3mbg/R+ky+3X7AyzsUx8xYAVv
+e0YQSt6m2pUZRwbwnZhjh3uD7xK1bR4JDdCMIxiW7W241/nAo19NB+4vRi2rKc/sXh5XVeqh7Jc
F2zJ/lYHCB7qA9tpzsAyh3tGIutDrnfB2WFo4MydEF1ju7ArJDTPV2lCcGdwOXMnAHBIb/z+Upbo
z35ycIiX3WmFik6L0VaFL0qdeFTwrRqMm+Retn2pc5S0D1I1utEizMp7rqaXmYPqUKqShdFJqMl5
r9lEFCaUHQ1r5OuVMx+gteO6FDOJ7lcB8eTanTraHVBDARoZl18Ju1FY6c0rgcfiVJ05c4X88WY2
swy22DA8zPioIOT3KEUAP7K9wDa+IvQLP+p64CUsR06qi6R+CVkib/9hT4x8vd83LlxDp2jYeQ9v
qMNPE9jOWNybf2X7neC2F6hISHiu0Pl/EvQgPfBshthnmVDvYmndZobjP89pMc6MJby/W6IaBTVI
260myXlYS8A9jTG7fhNWoKqnUKXqnmjvLO7OFrmrwuf9+PGFiwuMETvrEwlVL9dskyNSomkK/E6N
5BZh3KHIM/LB0yqJJsRTyJ0LS5AGNtCd5KV+0IpbEHlUjSZtnyAJtgsWBa0Yq4VTIxev/Pqzs4gD
j2uCiUOIZ6YW5Ofet9u9v1EPfekDOA9ZGUMM1nK5cuLt7M+xa2ochjb2ukKQ25ZCNFNPwIwEwWcm
NZzPoEhAJkS+MEreTFHUm9er0ijK9dBikD5D/yWWjIcvnLKcez8FSm6ERIZy/00e2nE0RpdmjsGl
QAUqmvAEXYCmALsfM8L4ZMyNFIRjxnE7Oc+PuirDaOXMXxCBEwh+7Uk7sKyMJXfqTegYaJYwNqmT
eDK3rm+nYYBAndGuAt8EDF1VH3exPilf4uzTAdg2OTpqWblm4t/9wOXX/3dvYVYkBnnZxkvbP6wv
2wrSLPV0ZVr9rYZi37dSGg3Dq9x84vlOQUpBw5r4bkCQX1GH8iPQwD9dDE6NWmBHox2S/yFvDSnB
VMj/Vwk+wy8F7jG4Qod3egbSET5SLdKFR4lvdxT20UZA3umuac7UeaPARFH8wPzXRAai/cpHeOCj
lY+SOi148uBbPeSlkgQCF1q+UNTd825japHzIOQlVtUIRwEpi2ixLqhKcaOcPgduYIExoPHtSVpC
tI/PQLwd1m3oFN4sD4L1piu7SSgVwWDDaC3XV6YhANZgHkY4yL1TUeWdiKxhiGeOa1EWqKrNgKRz
bzFE1b3m+VsLg/9if4AXO7lpWz66RkawsYxGv54u3hENi6hrAK8jqC1FJazSlJ/QF7AULgLCz1JR
cROg4S2b19HesBZWttdtQ3+MhYqoss3mLpS+AGZCP6e3MJilp08VJd3CMcBkNJGCVZxLEYt+ALiq
bZbL2g5YlaLTr8U+G5FElZAPLQF0CjHSCazZWs27tiBC4g+Id/DUYcN46VgCsWMpAEwookwuPFB4
UVrirDIDUpZwdr5rMs6ncEHQeZC+ln8JyxF/xbvuuaeGGzegHQWuMEuKXyPeIyM11YPwgimMdlig
bUk04V15SF6RejyWFMQcvO4yMG4o74Nag5bqcxAfY6/YvvXOCb91+bmmwyLVW4ufmR9sz2QAg+R+
kXjDBH72FVJXo9m1h8/xRCVcwOgfH1Q2624nqziL3KaAcSWP28jIqjpIQKh+b8q/v6AAfvR0cj39
vg9dHxajA7U3j3mwCu2DrB+XdjvyWVu0K4/QTL2KOKL+JmAUcobKFw9MiwMFoqtqldTGgBVQaZG/
Z1/s66kci7uon80yjENXcNdwaMps+hYO4KTzQFN1gxaRo2kx27gtjVt4r65iYzvd8MLY8ckoa0Hs
5hdvNswitA6FRrMJcJQ9s4R30DZ89uQ9STlM3cq5UErHUriRCC3MkKt60j4MRRTuXbY1cO2eCzLy
Mt+OGKgLEJY1KwuR9xrLJHV6R0vHilBaAMgdAgMkFk+spYaFdhnaG8VzTl/0vgRkzvVxRG1q53Um
/oVgaEC6vHKcr9+Qd5nRAeD1mhfpU9lV0/4t1dgDtxfg5OW0wvl0JwdTBfI/dR3sUj84u+9MJf2n
gtSUfigt/M/buDhuEgk360oxjF1UUx84IkdZLdXPKIWHIb7QghJmEnuIdnYE0Nhrke0+AB9io6Fi
QcVG+AlOyPjY5XiGFLxF/Bc2Ij1qJLTi68szqdQkJwJu5GIl9fTZ8CjCrBdNK2sWn5kPPBZrvf94
t0SG5jbUsyK50VuUfVPRdEh/a9t4tBGC25EJp0RzoUq7/6gLTrdL21L89zDr6xOE/sGfUtkhG0N1
Uv/hpNLzXHkQdLX2ypf0dM14/UY3KmNzBDabOPntUtiUIYua27j0efQk7HKsh/gp8H/ktQomgFCU
HnqK8V68PMPBVMNyfZPMChELBlp03A99uuT1Oysi93Eqh+S5kyT5OGtvPRAUeLrKbt6anB3yRHpV
+yCG14Jp/S1U1ZTEYH5fxYszSXijLD7/7lxXK9uK8snJgsR102RpKoUEGABfvGSVz4Lc78upVwjj
5QOUSRXM25E4hPVxfpPEHtASYH4nPmX6kX3ujqjxtf6fxCTjScQpYS0r4j8dtnganK8NIXX3fC6H
htJDLRydpit66/sbiPD/YBk4wk0mcH8biBXIVOOuhPxNkTbKcsTLEjBQ8nz3PK5KKZyjJSEFUjvy
+YJcl2Hp/p91NLJZlvuRptArF26Juu6mO7OWd8pMu1DO+4YzYjQYwBzJsz00auMWiPzX0xVviqxU
iPKRs6+12/+OxcZG+9LasYniYxTv2UhJZ6EVyxLpXPnGiXvRVNAhkztqqENqOt2OyRUaOTK1lpP7
TCwbX5+hiwQmp8/Ux+nYcJJ0jC29sHve2r3WMz7kNi0NSJYai9ElnRNFwWZcd3FrKI91VbMVVAv/
/L1daSEjzWe2Pyt4T0CpZf3dhuH7WnrW7+MCEePL4XdPNDy3B5HYYnNg8iEbfEPru5lIKiLm1yD3
SY0VrAeRdONxcqjuuClXUQGZ1KFECoIxtUJQoYJ46KTDXeeU2spYL83FRaRSIcQTkMG0CSSq0Lxf
Hv3fqnHJVViLf+B28twjxd6+OBprLcjrELCCBYf7nvdIK9hXMyBYsCNYIPErCs8IF8Ni1sv1pu2j
mVm9lrlNp10uynCBM4eDCzgyypuJm1ZEE8+nhptP6bfPMbXGwjmhOiJ54gZTJJ6xAp3cxR4ENE04
xMaJ9HBDH4ByNwiI1t3sR4Q0nDqa2+2w1LZpE4ZEzhiJrMypsbJP9MRuqpYYQisbjH0kIvc7eA1q
SUtypvX+UEX8TlLJRJX0niSWIn8mAvnQhsCFmNC6SATH6f/sgdb/j1hff34wDRsfwu6HVMO1znLy
fiulSg7sYsORw+D+nOjfudk5N3lKkIuX268JZPNlS6z9xqGIGqAnfLMSMLyeqNBNU+ZIh1myl7Ea
75ILIZp0jOF/ijZMcydFEQsA9nUjsOZGNo69sKAZHqfqswc6tLetUZhZ2ozBMTry+mGAHhgv9Bf6
+a2sU8sMXWOVJAdkFIrcpYqJ8ZRMOrx9X8tttzN5y93MJuyUadtRQ0IAIUp2Jn7BIuOodkD3ZLIo
5jGDL7JkM86uGcg2L9S/XqE9vjMiRJWshoKnY2Ebu7hK3rsGA2X09XnsGxfQWFIxsY4uYjr2XSs+
ajWBm06WCSyisAxu2jyaP0Eyq4QGMlN7UcS/L6mAA0+g1Qwpmx41FwT/H1ubIzg2UYRG+IO3rLJ5
LKYE4Kp6Xo074GLfwszNKI3UROuTuJiEplLijQTXOekl+VJShgJWw1MvKEAYBntprpcu9RRpSlat
8mNgbBaLrSYiBPRypgSYNK89YSEVa5ImqUN/uEaksbRU4TxG5PRFLFS3LjY9xN2Yi41hrz8CDKF+
+ZhQkZfy/VfAJ5/90cDe1M9MwW/L+18ul2KVwUMIB3qsnsOWKZIZ0FLkIlHMnjaYXCgUMP9LP10a
VoeOI8hYyUSq1m0qhHMAbqCpV+CW9CnET68oY0euho7NFqzHoMK1aPP+ntb03jY/EBXaKempAGH5
Z+1GSEt1o5dK9s7MZCOJx8QUDdZDd4YIidpWYny3Z2BL7wRvcO3p/iBeZYhhQII0FrcQMPnwe8gx
JY+4psoufzdyd3fvptabs9VfnTxp4Zb2PrZOJ1hA9sP89aFBCN2CuqjfO4IVMpnmJ2TEM8xG+2Vp
guwv0zLw0rNwEIVNOzLp9WUWpS+rno//Vz50ndSUAKkHCgzLKpOjymTBbPNtHPfT0Sx3MaCXyE24
dgj1orQLRhMn6VywVVR9MHnW17Juk4NOH0aSr1unrhXkD28iKHIax9FbxQCkg4YCEzfGvHqAQo5B
3vAz2o2z/3f7mKPNcgWX7MmhPU95ZTPJZqIyHOwhXbzkQE8o0YXPxSJaGuWNnC/lS/B/aEcDn8gb
kRrrTTSc57PkLbVXl+TrP4L6NWG1HU2Pa5cXyc+o4A/vuzHFyFXCHjUaDiPN/muNd9xEvum4fwFg
RZ6PvRf2cNM7+NVz/M2d/ITO4SJMheHUibdW3f86rsFMvAhDirUkxKHMRtXQr5P/EhEWxhD4KyrK
RrvfXAUNUwauGopaytBnDbO1scH8vkeVqhjIv1ZSmtOFzp/A6CDSf5Qq6Uns8jO9dkARh/3kMsGC
poGmGNy4Ol35oAR7HBb4nC9YTf3hJxySTPEeX/2SPkp0JABwJBfZq5ZxXw7hzXRdxnHvZiTwv8Eb
aK3YN83Nyg344vaf+9K2RM81amgD40hcEkizUD8/I/UZ6aZtJjWNPacBNA5Weh2bYIej2PVvBVdu
IC26puJx5dChxTupUdmUUzYAouCOxNBDp5o0RrJTH1jUt5XZqNZGqfJmP+1jfBFWd4ZmhDAEKNMi
XTABFY+0tP/jKTsogMgN0cb0qwDrs3l31LrEGXfR+cQFy+ngGcsVlb915qz0oaaue5h40fWt72cW
tDVo+OtIQVj2B04u53BFT8kPi5I9FahrvWonqPj0pOOIAe38c+0fmf7BOmN+dz2hReDMXRS6x5vF
goJ1D0FSlISEIqTq+7LKI/43hRKhff3d8OHSDdUMDhwzRz18On7j3PPr/hgIkvt9v5hlNvi1NTcm
lUuQECtOH7zGVO5zYTPzlGGFgKMSh/yc1tNqb4MDM6ws/zSh71c6+18NAhPsFaEskKNBiVG7XIlr
2kN6N27D1kB7LONY2srGVvETZDQoEtMCoNqaHxVNWszl6RhIWb9IOi7pprWT7pXD5iX49isDwYwt
zkTPXzO3eCqmmiQEzFr+nfML9rwZByvtDRtJo7kSMF3FZqhvuSjg5AABU9ZGlbsdzrzC4S5goUG2
Z0wiYUdgm6r7+Of+oMoz1IlFsWDKABPAHOXcmBAI41u6pEzDLdUPgx1S42cLHTfsBe7M3+i4dGFy
aAqPCXDh7XolCWTYMaleTPwJK4HlhkO2QMw2U9VsDfJcrqwKoYDWiX34i1Cw44Lq+ByBCR0NTE2a
uwL7eZ41JkpfP9va8n2wBp0uiaLeFEk3EZwUBSly7wnOFeVGZmyd66mABA7V0l1jTnJrGvOV317K
6FmTYSUz7+r1r42BZPP7tLhXwLajndG1ZPIgiSjSo0VAcJjaYesTpuihXIQgnfbf3QRjax1N1Orz
oxIilN8lRU/ZA94xn2LrvNNW3bo1kNYR2wnu+84JWt8IMWNKumP/yKkOlfTkXAmej1JtOL7akJuX
TyDJI2UPMlBLn25W67tXAgF8zdqjxKwafQgtf525SoCL2nzPEDbMov9q7MiN3IOMh/9xyxii5RTJ
18kVScJ5wFdZTNoOVvAtaD9MfAV8AcYHUgveFLqeaHn/7GEV6wirOGiz2GA2y8KwEBGP6uYXo6o2
f8C0Q+dP0xhWEnZjkmPH4I4hmjA35bGJJuC8sZKWaNRpb2t7Mt7u3qpg+V30WBeTqAI1JngP9lk6
YDCDZZxaTFkdZMaI/b09wm/gcMfSIWFuCgQNyrv8HU4/rqusjayU+CgNgZwT8pIV29CEHRnIIw5V
N7llmnhCYO2DrGO17i7t3W8EpprxTd3QRyh9SxfLOPJ/WTjeMJXkScVK+NpLtl5ob7aAHrieZwy3
2kRlfQQenihhlrDR+Azq1UxO+OtLCw8+Aa3qYGjAFtJ9Oi5f9SfbMfhW/x2dODkw9jCGO6LOekLP
Po0VsheCvwhAK3Y17jj3l0WVdxgYlwSCDXzyGrs6+EZbABwQCPXKN4sJiP0eGdJ0HGo6PDAn9Tn1
l57/bnzh+qC89ZnqEUU3c8aCzTxo4Dh31RNse6+RHEvFZiEnUaELSTuoZqFyCMAyMVXa65WcxlCV
YPiPXOnveDvhjuL/vql705mjv0eo3ev+QvG4tUO427Zf+g5M12qJkDkJzrFhCu6V1oajQKihzJeJ
TtFJIFsrRwjz7wO+99bEitjPqihjbC1VnVR1jULh+LjmjyF8ZoC3hMRcG5XObM0V4Og53lfV7t1K
dzsX9IVQ5FifgSO5zjR0ISdgt58g4xTZ2w8TiBiH3fBxH1lnIzdJ+Zri01vU47rSR6y1fOyDSUEe
rxRbpL3N85/rM9g53WOEAdq205/PE5n/XwMRwu2lH8hGDRh8ekdfO8+B4q64XNJbPodBeoIoLRwh
/RZPMxBpgrjtxVSgPKoYwiHZOOJbWSTWWOaU3oQlKJWNsNVmuZI23nLf7psSxXmw7UntvgrKIlOE
QmGIk7bEillwNHlh82DZ1MjNx93iXhoCwWEoUZNoJg/PJKJLj/YdrXgMaKF7Sjduj6VMCbvbGzeT
Z4Qr4C49wcQShj4W3lX+TQa92Vqn5xdXmeH7btI4qUNaK+OCc60XTLT2SDj3ENoewoxA0Zn9zgyy
E9u3Az5x2hNGMaTvS977GuWT4SX3yUmtE0js7xga/hlMR7Y6VPluIImMRLuvS5dmSSmYB3p3z356
AzJunWptq60tHTvlbLYLas+dS3Xul02qmYG+N5o7rIRJm9X423JjWwpck3G4boZV+xiVKW5mDccs
E3pEIM2F0KsstUvxW9VDI+/nCtnQzt5XZVITMH92/Phu13IASv+XzR9Y2y1dNi3RrPHcbSFn7Zys
k5mzRmUcxAKorjtgeT2Eq3cZs97bYxzkZWuF3Nbj+JTxZrL65+Ci1tM9lG69pKb+t1uD07nNXEY/
Th8NzZn3j6cv97qdIHpw9CNmS1tF78+7JT6QHxVSzjqACXje8GH6qDeGbmhbrrMi3FTw/QXbr54+
CwmAHpG+aostb3o4YSLbkeE2Knbjj7G/dwE+kZgHGC+F3aQ+Se5EZxJT4Uu7QdXwik3T+IWml7N9
Wa2KUfzb/rrOnMGD001kIFUch0t8bFElJqQZEVSxF6f/ghLg/gAzzXVPVgFwyQaiPOTSrkV5RcVn
8eTSqLtuvGdMxxR8ZbbT+31pCQJJj0z/6I9FkIgUEJXu0MukD4b8QXlf5L+nRNlJhCT+b1TBo6mX
cJAoULC69qMVDdSQ5ssYiYuJgdjG34tDo1mJNzUJ3xOEalAJXapgfzBvIsve7O+ZLXsZ5WFOPCUK
rJoQIM4MpHgebsY8XVHTH5lFU6bN4UDBj7WmL9OiVTDfktV8811DU9CYBe2QlAdh/zcOY168S+58
3APd7jT0Rc9/42z1LIKwgCUanHKbJMYEHzf9wwE8MM1QNdWgDml4GKZjul7gx6ZPx2N7VjnhoSgo
atp66rpKMechUzwrBrvDJzcB+QUClpbKGudQuStCsnOXK1Ee7HWiCDgSlFa/IB3xNPz1dFY6a/Wq
sN07wC27adIJKDat4ByIOYZEyeh3EXKfQ+4jMC/WQra3OYSpz5HG6E5+6syTFpEjfmEUfvII/98S
LkjxFCAAhRlJ9uqawf+++ym1NR7OXSC7MzRJpveRkhABly5oWAS5eCmfv21fzSrDIyzeugxym4O1
IRBCDIqbcor5kXsJzD6+2JAswKSWOpUgh+gb8QHu932354ty2uRyglNqltWaL4g6vc5CDe9lXYUC
NFXXILpa99k/A45YTlKI+HvtFAxH95RTcro02S9cYhkQUDjlSOrWpn+HW4k6I6VmkRTSpILPaAtd
afJrPFTnS6k26HYfJEMJwfVmsLihVcRkjki1Y1ByGCQWvIMLrBzUVQOM0uABHzqqZ6rbhm1UJr+z
3y9NbAj6h7G8AO9UDP5BQeGTEr9BJ3lApgqatvRDXFPPBxqiJun5VaCiz3WDl6KHvzvYPPIiS61s
MFXY5LVlSRCP5upUS8Tqw5A9cfugLxHQhsDby8WLB9MW5vN0iz3joEs8lunPfKX0P5zUTHGolt2b
A1Old/HAqvFPnQZyH/3kHKzA0M14nM6LXQTQ/8pSFaa7gQp1KE7DMBTwR/meBe8M3HSvh7agEIcU
mHMeZJCckAtAJerV3ipBP7waH0gjCoTh/+Km7rjtlMax8wx7lBc5pXcZy+n4rpegqMLAVM6ff7RY
U1M6GJQKc3+Le8/qEvykJMrV3BQOFG0x5tUdLI8jYKsHqfqL9tioU0fcdQk41YHr1D355+j/45Nv
8ywQikvEVh5VX3697aZRbSukmy4IcYqUx0ZFzJEFhgPBudgjjI02IFT/ljv8sVlU9qOH9V8lyvjm
V64gygLxwSGuHTLlTxoLgdEIFunv62nzNaOAszJuUkySz8kfSYlEn3Jk4wcGt55AgCBpIcPRKWxc
wRpz8ftdmuNk3xp9r1OkWFCiGnW9dwMm6TsX/Ogh8WBCdSAfO9X8Z+nUzmuWxHPunRUA6fbvaVbp
ipvRAN32qu2HUd6uP9t5+bkSva+vs4NPT9S04eXzDZQmgmp4Ba9H7lM2xKJO+xyWx9L2GXChni/8
KWNZGSE80IHpgrr0+bY5htq4E240ucJJmk98w8cmYWR80cZd47MPl0GLSi+QNNftNe+S3LMFiEor
ShNLIzusgiWIvBUNaEcAtl3Qj2iupzFFfCRurDG6sE2OEVn1b0t/UOHaqw4DiRxJy9Ywz6gr07Ra
DClnD63+gkgJwoLP9blrwLnXzWj/Q4s6MRACGIQACMbORfoFr6TgX88TlHRJhGY4oLU1qOLLmWf2
uRR7VHvp7RN7oJUap83H0JNCNMK6m3gLV6U61o7TnXTDVJZllM/q4w2s32Vfa2BalKZCjL4iM0ji
mcMx8kHp5H1O+cGuBVcihjIqknsekKe907nCg3Ux8FTCjefWYZGnk39Me10GVFUwVIb8QIT+hUtY
VnKthVSiQ1lsfzFazdc/YnVSwN3AoFyh1LZByzQCS3lnPAGws6FxzbOJaVXEF6VvuwzYWGCoQ3kz
F3r9+mC6RiCcgP/34u6pLzMeIOw6UbGRZ5WwW2Nvfh9+J0kH9TDSfTa96DJPtXIwl1qiCHkNqu/y
IAVAtNF48ri5VXeJGONstsUkJW5K2AnS/Xqu3b5jCYp/ptiL/WpoW264gmb0a/7clNKjgCjPEtz7
TWQ04b3HGvmOpQob/isOBe14QppKJurbrX2nENkHZMKQ50AfHx7rPSg+zO2X1woVGeDDgcTt0dp8
5nIOF7/kew1CiqSAMpkjK+IzS/C9BBnzkVuJU9ErioGzq0ofP8eqnzWEYpLv6pPubCy8MH7f4z56
T4xwJYnt7T97YaOaVwHqKRy8YhScvkWOXb6n4F5v1KW8LxUsUlh0WHvx6pFwJWtA1rjiZxtQB1Ro
uKPGSQUys+bWFv2R9wpg8q9iDlf6lbdV0tLyIrV2Q9XH/QHp2xsFeBROdXK22sC1DkKzaG0qGdu9
0mfIOSvcIO7oFttX7w7KURU155KvKV9BYmoPE3+GFUz0ma8x8xOeYU6osMMfAVHxqhkakWKFsfUE
gyyF72tWHvKOVfj1RmSltYx2zomJkxzAPjuKPphBensczYBey9hXIV9767gTap+0Uw6KMNxBNnqD
5H/slqLVcrgjDt4GlAxorLzxVxlxYtI/cas7iNaWh308QCIq1K+SeTqpFxtunPZI/LGJS/PmvXf8
fxNiDoikyqF/RAhMMwjWHpwmqWu94eV6XxFvPOAzfdypMRyEN138q2gfm3dSE10n6TNl3vKjYF2M
juELUBZmH5o9J0R7h7MPXl6AEHxRWzFC7fDbDBGnH23rGJ4ki68VqJ1xe1BlnWBpRd9Vq0wZJxTJ
jIioG/m13tqHuL2fovffY3eChkXOatTHcxS8ndDo50VjaYo5V07IPhatNwbvlIMsf3AaUXc7Dhck
EGEAKp3d0tqh22avWtlGR632/xi1u9slf36ZEoBXGeILOSrpZ6of7B1b1XO2I32jQ3WA1zk1AZ+N
GOGd06ocuUbJ8e+3mcbPvgKoaMCwI4JywGXDGZK9wNKp5L2xjFKdQ6b8oC69HBS0lD3E14IbRZi2
PcgVYvFkfKZ1C/iguFx6zovIXouFdnUaUIEr+bKkqCrNn+gcEvFTZblILwn5MDiHVVQjHw47wWwh
3Tkb/i6xw+4Xv9xpq1yzIwdvC3m6TTwvysMv/9sbjP3nvLUdhD4QKW+Ldv+g8Hs946GtSkrTms5q
1uShxPJLHurK+JdNUTo3Dvjl9h9nA9SkUducZtZRKYezJJebXFV5Qa+L+88QV4vF2tltxrXouewq
btKyGDrlphU0Bj46oMjJC+VeSYz6AgUZzZqFAR/GI5BGsAjK9EN0nlsRN4IEsXzOmNxexIiRoR2Y
mKXn3xX6+ljXfxyyQHjieP4t015Yn7fUTUIPsXTTdcNNCfuZx7/n16E6dYC/vZOWASoCe0zDp3Ai
/PPixFMN5WHll0s+oVWFi368jNSKs2SZnzPrmO019qG0+AYNhCXc76ANlovuzKEUwOg5DM2oCaMu
1gkW1tkgDMiNDyzr1MRraSh+M0II0UNnFXpvFLnJ+Fj2smOBdZnUX0XjUTV+toIfjX5b6FUcS3Va
GuwDJh4DJflBDyls97C/eJpkoR8lPfhwNVYtvdusVQGC2dSVLuA7wCEDwERAWJVEnXLV/ZOlu1Ov
mr6VGj8Q7Nf2fUJXH4pBszoXv5x+M4mghVHUTj1GGr+TljQxfkPn7FrDT5jUJzqWeSc+3i/yENIO
u58MDd7VynMs/TXQMehMFysa/D1NdTmtC7/SobMWyjkxUifCs9YfvCNwJbTpt8RHD8rpDIvinzlY
kVVJxOZuWDeHNtJ7doJaf9OkvHBfpNW9esi20erL9c1wOEvMqU5/MD39hllS4liK1wx0khqS5Glr
IsYi0VHcEh99gEzMRjhaRWDah5oAop/XbRoMfFvHQDkNzM0A8eIPcHADqyU2HH3T9ZTTNnQG5tkh
g4IwYY+oMOEAtkq8QRjtqPuisWJP00rfwz5K8hPRGUIqI6/GzMyln+KN6hiMf2snDY6g0dP9gi7X
H3YEu+VpvB1d6+pxOdBsT2E0du2FkzNLNjdhdHBhCmSQHflnfslVsJ8+sKDjE+/U/JX/othugEol
9K4f74bC/h0/t4N28bwTtq9n+avo07KZRwJpTlnSZnNyXdw6Y9MSqf5pOFQxlXbjh9ndQMzuZ9Z6
g2h6DgreDU6XrqCLpltt0FNukgDMHqhIlBKAoWfHXlQPOMToa6hPp+C5hb8i4ZBJMRE+uxnRlCIU
w3TnsTRx5hxz/eORe9TlNidkqYGkmQBxmfZruqh2CiTlmyS/xcZcGKnysQJjXJDBJrAMmYIV+AoQ
937410T3NN9nIDZidFsjM7PORg3G+d//sNuNLvo5W/k/BqeBfqOjSnZEneOKttbBODcl7Xhq1uGU
HVOzsoz6VCKVh8KHKlXupAhvYmguU161342waINQVo6TOydwDOHv/yIgVY2KOF9c2k2Q8G6VvR6s
BhUheyOI6d1q2BeE5Wxpq8dSj8eJmBhzC9rMHtKWSyES/WLyUnVh1SHDM5iMm05frhixO5RT638f
7uvO4uUu/QTOivAVEhX3fFzD6iQJCKaFoow02VIgPW64cuicoUyuwsNDZDESCxK4UeNoQ+ZV04Wg
6e+q+fnfIsgswd/nFKWxIQacSBLZkOlk9FE6/y8QANg16LtYD5AMTXqeEIRo2KaeIpiCePqlOYPm
QulkisaccfyLDurvOBIKaIrNeiEUGUsZax4jSH2ajlm9WUf+SwoJx4tznPCv3WqSxuQgIRMu5/32
xfkTmvWpOlQuCmQ5org9Fa5ZL1XCeB8sXLCrEkmhYmDBuVoHXsvhtCmOqHlBydV2545El4mupA2f
o1nAeShl9rCcgMeQft23QpeqTchugE2UacxvhMazs4a8BdlRk8zmayCxSLtp9nrvQlMqsiracGWa
8dCIpXUxv6A8zO6NyUqnbmeMhWYgoXlBoHMnw0PjXEWMhD91lWBLTT2Rfesjwuga8dkjJIJGoXcl
CiD6thys18cyWA/KE52wT9tWzr9H3lJYZ1FtXAndsucEYLsuJ5rYVpmeX8pextXp6dKhksQZ3uzx
G7WTffxK4Uj8sWQvJ2N0rhuPYm9wLH+pMtZ4PTt+Wdln5uV+R7ktThzIfqM3Ulc13HuJEBISPfpV
4bDdV77DvFv0TBrlHCfJ4kdAe10mMHnIc7f0slquRaIv46Lq+rPNjtHpLATDokvU+FacSYAY7kUv
M2fJoq0CBqEzfJ/ntah5EDclwWflyMmGIUGNIDrifSoE7SHnQv8SDJbZuzn+cq/waoX40/LEim7E
cl6/zGR7jvvEX1gXsAatPDcEhDgB8iyRcYSyiOpx2Okm8yAvAnTE6NVcDMa6/qtUlWqcEbndJ4bb
bw4/BGvLx4eLGRIa4Qqo2ond3o1vZiEJLjq+wHrXOImErlSjVG3C5Ir6No8aeTExtIjCMs0fl3VS
KdMmSCxBeZyw+yu99T1xTKy3pkkaYaCIrk8Qg9Vtg0PAQb10w76WIkkmT5eGyPAsrekF4ezSmoyC
W5z7sThJbr/6qjF6zYRpMLDeUYeX4nXOrtrw2cnE2HryTA9yDOEDQfRuR3mTB7vmSkc+RxdODC72
t2qfmFCoY3YTermLAzOhgYw5/XV5suW6/sg7bwsQo27PWwio5MnnwGiR97vbL+gqIDOGmo6rMNlU
LoW6c4fYBMxQUrAGFASWbP5DjurCWk7FkL0HcvYvtrZkmIYhWLkGkkZ4To1/CVefUsXuDv7r7ZdI
I/MUleEQUgq4x2UoypJ6Xy+g+qskvppF5xW4BLjnHI5BoS9ftkjRMIv6J7XswRcxFNg6GutXjNxg
km9EdVeMqTpDLyausxhR5q0uRzTHeH4tR1WESYmmkG7NnUAA1j2+B6rSFo25MFCJm81X64TJeID9
cDVfgceo6OhKQHnmFzhGWppGZFemlh3ITxdNzwubQRIp1OYp4AshqDorHIqA7pM5AiWqRyF9h01b
mLM4Zn+XE4/TaQFx/04hmk0L48E0yLAONWc7taBa/bsuEvc0l8xMW2Gd1uicOdRqjSL0NvUDHJhL
6JnOAuISw5eoldBKNWzq0UiwqlQmo/xfvr5Gnx1pWQFctRI9abvQJ+POgb1bwIACXtTZCx/Qj4Uf
adBF/UzrlfpE6Wve28IeWGb8eqAOVVUCvmWwY4av81VGSuURWG3AbHz7FtBxokxKcFXpBfZuy1N9
nXmxch7FREH0qAPQY36gBH2lQGO/PphjLX6KK3jaDuY162yFEBFQiM3fSX9H7j/OUT3OkFh7vpyZ
BlI4IEzSHTt8zaen6AKvmTVr2zG9FqAoXWVf1qpfj7bmUpFnv7wKymRJ70iVibXn9uuPcntPgO/h
rMy8V5wGe1K672tJy3jttHM8lUU/Sg7xdswFKxhO4Vqh72lrDndgASZcHYFYHx6+nD9FXZrmJOA/
A3vTmGl49hTJwrZR4cWfOKR3mZp8VkCkEDnZisaHxCEh6mL5/f5OCyskuHDvH/bGUj0EwoWQ+SgX
h1hUdCFbz7DCF1iImMM/CN4qrlwQhAeUBqhkSD2lMincq3Na4kjc3y1/QW3iC0B/elWkHMzmS3BM
z+PuvccdExmeQ6xV/LUgEvuIqxy6AfY99srRtkKxFh1mpCANMTDi+2pTgK5Kv5owTrSd01J9shDG
i+Ptqd9+LfXNMvIroxgY5/10rWDYYm8VhPeYjWyexHAbdrl4MmwgA5JIVDy50AZHhf88qnobDPkO
NZDSIbLBmQJQehKHRpaVjyC1PTIxtLmdvqBNyVETk4kUr51okpRBlWsZhOxVss6Hk+SIBdX87nW1
6YdLE8VYIU3KYglxQHoEsNUwXos2SwJsYqibWqoin/JbYn1D2ZHjYdpQdIDAYThdbF9NzSOEgE5u
Wb/gFIpWt5MXAa+klrcCPjetLRv7XcbCLSCYZSAVSapjOqyWMvF4RzSOjs0+UTfolcmQsy2GG5Hd
K/TZfwbCiKv7z8T5E/P+P/187tYAM9p1ofo249cc1MSaHoNbfUjD/O/+ENAd+vQzEwbf3CWGFZGk
VDyHTRTC9ugng292jfe/ErcUfXSkyOOvt/isgePFg/YwAkETYtVD9OINPx393ChkIDFkCmtBHddh
9+uoku8FFsQ/fzHp8SbeDNF6Hcnr2aLnOdtQbvlpLO7jsod0pAaSXx1/8p2BA+L9HJ9GrE7oQVFC
wgLnZlIbHUxTOUt/HyuLhwkvbyIP5CzFJ1lnZ2pyUwDSHFdzVX29JGlo5lWQ9P1UMAJMuULb2pOr
anx6ZmHDrriD39MAZxDeiivxkp6gXNv/S3d/53IYRYxB7DgswFF0RZAPumXA9pVnqzLjQHZYSUCv
Sm8EcsbJIdw2iudFAdS745etX+6k+OtprGFDKBJPaNn2Af5GS3Ut4Z179R3OfGoCZT0v0VbzDCxP
B8YIN+zC9/GDTYovAJRU4Ci5iJ12Gw5z9zEsgePvRwxJR9KCFF1ehSmLBULR92EuCusWpGcvfMy1
lPOt+EAufOUZuWHZtwWQrF0gwb44VvawW7Q2ivLpS2DQwOqeBwKEM5Qo6eUZneMZgvhY7oLU+loe
8G/PdBWoNUM9fiZaX7+RMsSzdY9VFcsbjJUPZ6eWzskkB+QTFZ1UWak/tyX/6xZXqMYVasFTtjJ/
ivb3rtoNUD8d+laTBfUvnh9jevZ8DvvUXOVrB0g6VypzjN0f15Eh2OW+qtUqEnn+AVFr2aDi6ivU
IFlLneB7B380sdJy89xlMrr6omsvDQbsqSetLLg36CE9eQW9MIVT/X0jLIls80KHMNXlDcW6ZAZU
LQS4nAgDFCCaQBZ8ISRNuiLKVXg4fe8HztVC1qVrEN+NpUw7ndjFKaJ4RcnGji+XeqDDRoTXaLGp
hv8IGhSnyBB70v4WO+fKGLURiY3Ttt4ZzozaXXvbNFCyslm8ae0o+vDXQAyC3arn1u9V3lQkSjhs
55EGwdPpkCby9lKKIBcNUsjF9cpT2+KRIXgkFKHjj6ZIhEBgpeiaPPvCKFc76YHwNt2+H3WT9kWK
sth1O615B+PDq18R6IzPqaGWHk5T79Zud//vSxTcsJb3nd91IXdvrMncQXhFH3anh4WQz77i3skK
K+00NqHUvrjCe8pNfpOJi32CPYaAI/RSIRT0eOwsecmOU+B3LAsaZL/Nrs+NAfqiH8Z0CKi7eufh
4Oqoeo/2kvSYIMrqnUogPdSixXV0Zo4T7sXn0cnnqkNWK9tsTRUxXc3zE2M/3EFeoUOpp1Ihm4iX
QWYv8FG/85pwiGljY3s57TQUtsACjBS19f+KxY7i9JwsHSzwPXTOuQQKPtVrdPCDdqmABg/ajayP
Pop5LpQ0+bBNSjmgS4k2v3oevH1tEiXA0CQU0aFPOnhUfhfk5mEpmI+B6qL0xx6+mGAjlnI7i1d1
cmxWqFURx2DhZ1wblq5YDU3+Gkg3PD/xDFhLgY2XFx18SSzbHqqFOworLRgevkGfk3owOgt0dCVv
gnP3y6RcmAi2IXIvRfw3Ns8l7ouH3CdB/cHGuBpiLoXLW222417xCQ2QdMBrEAWbKwOJCUr3+Rm7
V1sBxrF7IlpykIlPcyEbreW/vzICqaoG7OqsyrEkV+p4wDqFhK3LT78dOuERoNPK/oSscTvXydHo
raMgfbz3WULCImQEacJGTXqmHJzoU3UuGeie8sdjeLAflsATX0i80W66Qjl3Zk1R0CktAS95EDao
wzT6eT9DHcIGz8rPp0vUAYU49F9QtBvJf1xKHMGVx07plDO1q78VnKcxtvFnTtVjAKK24TILzFBJ
R4ko0kshoITUY3hLCBCDSSEDQmns/MITs9Uf03PgMbVmLRhWM9Zl0DW9kwwV0V0xJXD68/myt0VI
ZbuFxyGgTdC2M4t6UIScUeBypX2I8Ewz380OAkJS65JvIHYgxYf/QcZiWcV1f8VSja1oumaih2HH
17LUuh7IDJIUHWZmzGdU1aXtqTi3hEcZW+Cp4epeWtuID3a/JWe9JHuMafMrVTsL48AzRGWCcDAB
rUSk3dIBE+/Xxjq86CcFlvdSwKJDD3RKkAwkS9sxvbMLfQfo8alDRFWzijEThZPUmgVAAGS+83AQ
M1ZbontyY+p5tl7RO1Q6QBEuatQb6dm1gyT3FerrawyNqDnx8ut7q+uaZyF2C86XN2dVmEpkl4Jk
RUUWSX9qoZ19+aeZwLynwdV3zTVZhs6GBAwK+Tyzliv0UyzI0RDpuYjXeSL8ZALrUbWbB+CKvZud
ac2Mjp/CvxF5OdMFNe2Rij/CKl5S6bZmJT7fTEhZl0VcouthSI56adyuh947OK49z20lmyDCHBkD
+GWfW4IM8YXiWhGCsufSHmPkeAFxCDnbuTdGaVCrbxU9FUxFuy3io6QYWjp/ZkRlya3gsEfodItH
+3mILMSqyhsZ8vf8Br93hY/LtErhbO0AC4cRbRr1RJgFEYIQfyBUTLtQdeRmwy6ljqLPDPElOGDb
e4kNwgSsjGyMWDVHBCbrosyKOdfRnIpHg+Azm3Tve1AP+x3YfSh9RFxIWQ0fXcKbRFDYcOjyXZ3q
SGJG21uWNctVjtVmgSRfuiDKyUQOYwvygVbnNn699solFq8sUl74uGj5pn7PGkDGYI26B/kL2em1
YZjy+rLkIZbJXteo17Cl4IPKHDy5C0UpjQQjWX1OuivNKNlDGIh9jiYiybEAt7UJc7FbZguQKtb5
hb3yn+MOdx+Q2nGDvHebZq3ahVu50Iaoc8GotaVNgYep4x4gEgYFxf1JRyoifW7MsdidzVQeoIp9
5yX3choqcSLBs6JcKhj52yN/KRdOgyhvBAZMv3nXadfTyet/E8plVe/bI+bDU/pY9dM3gawMpWD+
Iftu2seSIOrzi2iOioR+g4WGstAF0EYm5oA2GrP1IusL4adVQO/+YQH6dNwA3nRMSDeL4GPHb3Jg
kdhXTCmcuvB/RisvMKE1l9PZTlt0c0vqI30Z1q/jnsOQJ6UCrh0Ue6QOXWW8xtArkXYsGQcAzEb0
9XMo1IiPJMX2CQAumS+ArDLKY9g+dvLhFkWW7Hg9FLtq2iguaf6tRPHYXn3BacFykVOhWTRndw6E
/85ok1T4kDJwRMDMZRtahKrt02ZTVpgM+obZI86EovDWjh/KLT5LbaCAfsmhflH29/3mKn31r641
AAjKILsx+aIJ8mCr97G7dcCv1+yk5T+ZJLsanP3oe0xHNH1E8bnl9jiRe9VMnMB+3nVD6l5w6w5g
twvBSRzwWydDJPSuGM1rypcEB8RZbg+rQwqxrevOb4snTv497h7XbQzAxfLmgdXlZyphx0oLBh3P
6pOZPWbipkbIzui9UTGcx8ZDkzd1/g1EfhRnoS0LkbZOFr7l4KybvYaXTkKiJhuMHjube3tzfVp/
h5/1MoATpSYJDwb0ekaE1FVLN00DxLnb4jEf5jySyQYExJnUDXSJeH8xmhfjJiEq+aBe8kjkhlfC
U6V285fRkqGWbkhakEsS9krQp3anJmNyIeSu/Nz+UfbGai9AhuABGQM2azXE7zbymCBlcy9eTP0e
pNabP93/X/v6f0J+RffJJQfj58haP0xFmy9fMrFw9YLY7XTD6krVwFO32M3toIw7spmG2yTfWqpD
QleuVm7tkCAWYSYPLARhZgNAGytOW0t2pB2fou/dwkUQEDTBl142KZo50bm17txsEGQPeUNL3nXQ
ybodsjBhAwwbMtYyYThMTptYmtKIH+hxXgxWFX2PCWCbvLyGLXTYyMaHJFyKHcypqE37t7RL9Tlp
v0eN04yhqjHy3w4pkhADiOo0CvRKymfEacic1N7lvK15zBe2AfK2vx1uQtFVh5oFXqzXZsqN4cB7
+sBGqyS+h0xZAtN/5cldVn1RbUDXqc//7BFS7GxGtL4zyClBmnMHZBo4Wd3TQME54cG+R6q+bKZ3
twIhfkdYNW7Kxcb2V6ocgXY7u31+uuXQzBN7GAqcP9ImtNn8LBMcTlp+hqv00JtHzurM6X8/txQ2
CrtIHMXVI1twmx9fA5opuLrAUKVGeyZofCY7V3DW07dIxT8Wzs8bkdngMmQzb7nQqjFRKhOtj9HX
hoYmMPn1GjCWGak9sz4XSSVKl1THgEA2Z3DZH0R+25phQkV6p40gZ7oEvbqSPRlBI0I7Wy//wTq2
skR1j2k5XZktubuAF8mNvgdxuDoIDiBewrpe3Wdm2uAjUuQsOlCKHkO5klaDvQCU63HOQ6rBA5u4
CfLA5Zi2IDrZPLZgE00gFDP+hApZKJhqGQxJXM2NtPMb5P3l7UzDKFwiAfnF+XXaZCVkBqfuAQgc
/HUG1tiOENfoD1RTrYWKyMoh71sn0H6okOnC5XfZ67Mzg7wVq12z5yckkODhDBi7/T1tZLmPg0w6
1VFTyI8GDYu+VBAX/n7yww09fP1Ntv30Qds/fR/orOYS909ivoP8yBya9ESgrewrZiEl+k8bLDX/
7RILk7YpimN+auDVhn0zOgcHAusX9zebunxjpq/afYuyJyEi1Zvrsd4wOkzOcLVy9bIFzvDa4xcm
UcEFyB5DHz59MXCTOw1XDWkHub6Pj6ergivFEUE4veoY2ihSnSzTvB4RlvXqZJy7zAZqMHCN7B+v
Pi7kU0QSSKPvgm9LDfQKEX2f7+nMimrmZRyJqEinOLEBk4u71AVwqjet7Tbop0hGbSwOE+bkHc7N
CIAc+iOBhFAMUgTAXhc3PSpi28DNntqYxK1XguPXYRVZynAbDuRK9leKimuKqD1M+J/JBjppglMU
id/TnQyOHO4LwZbO5BXPgVIc4h87EEm51KvN94kqfr/NGViUXpu2sFwJ0m7CP1kCr5mgXX0JqTCr
zofsZ9zFWx7bCIpxrgXNnlujHsOBErGTtaTlq7DoLeZgJKWVOyBO8swJ0oYgf0usM9uUhQoNs180
Dk1CrNomPVALU3WWUZscKrOSf7L2WqoNHBf9Itb/1hD7yrl522qa22mphzRQZ//0+xgyacFcCaFR
ZlZknaq8XJmdG8UqYCv85h3IpbDFkQWwq0Puorxijo5cUGC4JipwD+aOWEFlaeENbrxgtDIkaLmg
Z+gXXtOgvbQcK3g1eJGapNPy01hVBKmcI/d3lCQa1Z2zIPgChL8fYnDxSZJU8cHd54jwVGoRYBW9
xhAkEtOFUespSLGUOMuf6J0zvO+agDRyMYCIHEd2rhsrRUCGGnx+FMr9tpEyAhFt45T+yqDNcf6f
IqqNJZzWyTOBlDT3Wh1gy8IZKO01Uliq03NI9bqW8rf5Q38nAuD+mlaEWPqzrgsOAdct+0tK6lyZ
8drT8SwaDDV6+BsYjFmnCliHR766LDLUHN/8uihemkGd3/7ycX1ww0YJzITguUjczT+6fRNDI80W
7P3sltVRvv8tqlVZGGa0Vp+qkegxG7hT8r5umRMvxAR1QPaBpNWFQ0HmrDFyZ60yOJj02ESOOrQS
/BjLaOeNXx0xWZq8/NzYCKcNQje/zF50s1ByoEQ2xLeawhCm7Ewm7YV1Q7r6SwWIoLsUGvjHSWBJ
kLFLrY49FbCFzcNzARo78LzCaGnwNVdQOFz/MqofX4JiG9+JBcrtb6+Y9jEw5f42SMb477QgIk1W
wQKLPgR5zEB/GwSB4lNCAwYzW9SJMEALMlZ6icQzaygqtNR4XoeKk86ISYrpqAF1vRJS9ePvnBdX
mYvJnVNEpIHV6GCimvOJd29MeQMjDoRYTEEs/aZ96x/aIHa0IH0KrkiMIESJD+LRvBtcxU3YCdom
P3I47Bg8Qr7Vj/EjZTSZM6Edwsse92nBywRkp/T9kXNzn8e2Jcp1RE6iiTn/7+Ih+HTNmBvWHzKe
E1WKqA23F6dCII+LqX06qXlGhBrFHswwLxb4AXR+aiO/UvOVECi/AHXBQlAMkPKuTCTDan8uVwnA
YvmWkJ4kOtyuV2/MzMY2+AmiR0D3aRskOcSxNARdfU1zqzGRyz1uTs3gt9S7l+ffTCsdwuAoP6RF
jc8jX3fFi3iK/YZ+pocHm0XKuoWO+KZIpFk+08NaPuEd2KKUWHmnYEwJ+l4cees7JiJVCJSNbF2I
G7mF1GYaQ/xS+icKtlJhlJGwUun053qFoyk63XeN8tU51qr/LvQuxOq7QPxPoCTgOV8ZbTB3Dh1z
L8RiLWGPvE+2AUp/W8EH+5O0ijC61gUHbrtAslrhnU/rDLQ/M4D/zJBOMGw0E0wvMMDiYFMp0Isj
8erAzbWbjWdKR10m+aLRp17oZ4QQQFiSDiwdfxpQ5TMrndCtWUaieyA6niIWSgZUZ/MWUgW4CZ1g
JPNQyEdPmgVJLWdJakhn8gJSYeXLPKIOYmE6DDvySGD/qtXWedWIAPqkFwu8N+G+a+Y84onuRWjB
8RdWfs3Jq4dUaLuKUkzlrnWOrFQk14tb5tcrVQUHFyC4pm1KiQd75ruVhGQEqleJjbeWMGwneDET
VuKvGgyX/VeJJ6PwB8VGLSpgw1IRWb3ceUuzWWUS6etOy2jdZuqN7BqzTJvMHFpupPLT4GvOAeYS
AASR/AbuyIAijNtQvunId4t2m8st5td7WuktfnSvyfTxlYjg/f+5YUnvqrtYbCcobSMHGyQDgPya
5x0uiOd5Fcunboe1Z1srHCpdZek+ayU1NpQ1yrLnpOWIBztJaxJxkUQHRNubhweSc7W5/RZ/y+ke
nG9JcUaXwf8y882yiNURb70aKk2hy/gbVbphTHpiHOC10vrmR1U/aYQftqz/8FIinlmhoPHmfZdF
L4ymnO7R9e1EVl2XfNu5B7vCYUk7y58/VR0UcXla7Yii//l6zNd4T/4kyc470NGdZspVqQ01bLE5
KY2b9U5FCpW3r3quhYiBdnhQLClRMYOrNzO75CYYzgvtMdZ8j/g9+xkAx+7W7AM3w0Cr3xJcgrE5
N6C0yNlwz2dnriG7pO88j7CktWWCTEb65yLOBKJb/OCARP4nMv1EzRylF+DscFYzLZGSV+Niu0cI
d4NWY1Fs7Ruqn4/lbHouIxcqZcUqJjjkYfWXiDcVU72MMNorA0hbdaBlsUc55a0oddF5KPTB6Grr
dQGEUwB2bNV7Utxn3Y9vtE+jAQyqP0EjB8KIV4XWNWOjLaLLxcKfoThraoXd/olAvuMJCeEfFib2
q4bc/ImxWLGaQ3/u/4jvjU00/rQu8wGFBR7fZNfXqGmWWfEc4I/JF+ysWmmcXVIT6R0mRKX4n/ne
E32/9tpOzYtJfc/7ciYvoHPsl2U/FevvNNpUFNalGlPJkemXdvZX7g1iX9ukvpxg+o67sAtg6kuT
yyxEjH1HNDTCxBAHZGfNLiXmCdt22KRvbTmVPb8FhS+ecjNKvh+Csvqi3rV7R8LHH+7Yi7+XmNrm
earlMYl5M5l708n51k/xNJRgV+R2/6x7voa7R7XphzoqzU6szvxw5H/agmhF4SR71xcYK6u4tvpr
K7o22vWpJSsPLGu0C2A5PlHwVF2v3kQhqmnTVeN1vvCcJL/+Vbvs/brH+2eO0P3nS6XJRSPwoLoX
Plvq5CM9UkCbGVITDYwbDdtmQeF6clsDtpbam2k48QwJx/CJ65dpnjypxcX/jN1GrFORQxKJKs5d
GN/K2mvWiledCs3tJLvvSt4LaBpxVSOwPOkQqs0ASN8wOVWhPxs8z7RFzaZZiGo0TUrR+cvFekKP
TUwUdC6iPldQATcBiAaADC3KTCepv0R0bzePa4cXiZLimcpB/kPa2WKIhMf/qAD7O++CGWfbuOs7
Ctc4P7shZijrNu0qAMj1y+z8FovhXszr1LBfQe9x+4j2pN4MUHrpg17xKBdwe04IW3KRF1qi2bGm
sTzGMK9d24A3jPqTX26nwLtwiL5SXb8/40xDhlmaKwSG1o0VEUgxHZlj4YhbxOcpl/oK9fs3Zhpl
U+lvtC0TkmmQhDkSUcAnO8Aw1af9L7SxfQlwopztiyoYjZ/3v1O53kSgXCsCFP7mIB7exsEwIulD
exq/JjpLLvGt1hIOIVuJ9nyj2oeYdo4hAEfIa5VTQW9WJvgPwAOeUaRotGTifpxuzhh5dyHxj2/R
cwNPEEQcVImMXAcv3ZiuK+m+wNV/qQfZV+OlOyQQXcMHfB/VlnLTM+sfx0r3aq2Ze126mdz9HrNm
nPmodpxxQb15q9nk0HkIXB5di7cGtCczCBBAZos4DJm33bqb39yQFmQTuLY6pNtRMHmUzmU4Xj0s
9N6GPnso0YvUpYOvKiWVitaKXiPX7noLvYUdqeNkxR9R5SosFnb8Jla1e9anvBxWSia8qHAad4Jw
lSMkXNxmVgTiLnRO2PESAVDbPFchik5GrsN2P9j15OB7qYEaIRi0H1nN+X2OpRYYLpJL6Q7N8QkB
EFCIZpKZYMDio8Qw27njJHnZyHclcowgnaR/x2QIkHTSkJv/LZWyp5S79w04MhjbEvNoMR/TbOsU
vq4+j9f8DQJn4IUrtOJUzrfrxqd9Jw9jiDSFJnlb2+g6XVxuQ4B1+YwntJqAC9nl5YJ+Y8Z4p/Ph
Jeo+QuYsK+WrlT7L196JqePuEyuglbgLDyOTr1oNYTlb1yu7bIyaTei4ox/Lc34mQDfDmaX7IXGd
wp9NxqQjFg0fa/64oLgnLeU38nYF2uaL5NIFeeszL1d4g3O+eYsRLw38pByEYt9D/FrpjkhIxoAN
TaKPylq+ibjeTq2nh5Uw1eFx56E3dW3pgfB36dPXuJXzQ6Nbg9q99UQ3UQs+pCL5vYOaruknqovl
JkRRfoGTDwvZhLNdGq2voBjjvBSq8VjkRvaWVL6c3d7jJWyJHb/Kd9mEDlRyAd8U4AteI6qJfpGf
tyW5IQ6qWl+zucbDxAG60GjpyAX0r0Mg2rp5BdD2KQT5FeVUC5Y7OTvMQAbTK/IpmhW3ab4P1VI9
ePk/q9hSWHf5/F7yGD0nidFLHAeMN/Q8BzisUkoa4Y/DkNiN0Muv8ChpivhwGM6dnsA+2HDI5q1q
78yGe+ItEAt1pNOASBUbfTEZqkS/hnaaUCBsGILPgSjGv5OpQhaLy+1BQh1ThlsY0KURFjSKJMGv
q87OuP7wrFvKxoWgoZWrIBF9n6H1sI4MHqTSd+hm5z0lDB8qh/0IjaDlFQ7luz/sADq8tI73o9AR
ksK7OnIOFWDVMvqgjfGBVS/v5xfyPJyCA3Y/yvVnPpFNS0iakVYdaYL6OtvQkAAacyVK1dBUVrp2
MHrpKKgIN10aYIgwWmE88UAbjR1VzGPhIYVkOvupaMT/ee1lDnRlE2Yp+eNS6g+ANyPH/VZDls3v
J22isqTSYk8RJwOrFxRLOUYHGKabrMo2b7cwqJ5Ghtu3FJgiiy4AR9Xdk2t71ivg6ZWiwjL2wMM/
77Y0dRHW2MgV8/91VuiHurB0lWec+CXzULik5hYoz1z38GqkaWT/7BLPbwROldtBfUp/RoeM8zaX
N5qu2mpHKab/AxloVVtInFDmTGWcoZdoAgHRhrp8p363XhcTE0SvuTMaq0CD4GhwQ46cif3i4uCv
+HX7oFKKVg5KjsL5DC2D7fJcgEgeY4DpH2yaH7ujZA1OgBLJ80w37QnrP+hSmp+/DTKNafD0ACjL
S6lgFVesZcSrabiBQmX9z9LT/DwzU0oAsphZPUrntq1dZDMtYKLg4uj7PPBsDsYgcn8p41DrHkW3
DbYIePTrSxhl4CH33ztRkWr7wx18KyotAtKmRbMYEqgtwv9UDfhmGTTaZYWkPJ0ZxUBL4Q/5udzE
fFcvxv9FDMqmbMi2ladpJRqIfzsVZqD9dRsrGilka31PCJZd8Q+YpmoBp2SIZE30tJaZA9dHT/aD
qWUX2m58yIdStPNa4zTEg0evjJjAgoJhJddETuM+6hj+GlWdbigQa/61XWjt0JXsk22hdylt5gie
OiT+XxpCElDtm3BaSf5AZrxzPZ77tdtvmVZ0fhz2mObRfmSQpkpf6tGWgqH9NqSVanBteSocuvzN
uKLXJ7WhKkuV1mWyZddBbmDV77342fRzIWcCRGvqxlnH/7A8rGi2/860UiM0EJ9HP+Ef9cGLu1ws
8fY3Ie8mAWPDLPn6hl1BKcLrwqPkpfqKqTBUQf6bGlVUPdAtXNUEcwe1HiwWcgz3rvs2WF7+K1WO
Y5SkfMo4a23sHoK3hWPpY0oLOCmSQ6dblSd/jiItFyIQUZl7J8nBxp93XLZoDpcfaiOD3+rzaDdA
W8SJZxUdJfEYRIYsUE1qUoipzNut/GaYUKlG/6kOcQYXT0iqQz5qbE1gxRfamrWPN4lMyz6ml2QN
9QtncTauY1/i9e2VPUBzb1ia5H41aY6QThiw/P5JkASRfarbFcDK/sg5rspkzXSmIlu+EN6gVbuA
YzJ6Cq1VtpV+RnA16Zol0QXFG/89N6v4vY/gHing/0a7zTFBeM13CWxIxNPTLiI4W8CXdEor66Fn
p4Phz39sQ62Q2+UZj1/n5wkzA5n8KeHsUV6QoNuRpyJt2IBqtO3BBKPt+wW33X+NadZaMVnSUAUL
Uxqx1dus0p/Zcwq2WkQOSLy+6OjZ1D5YSzdWoKdQn+8vPAkwbCeNHdUIMupyj2FnQtS3ccpYH17X
KAJjQITpw2UomKxshnJ5Dh0fp4o43Xy74bAMLSUj3uwD6yF3Q31Psetqkls+54VOk4IIJ6CvmteX
lp/1vPeatRkOs1IVVNbLK783qcqyxH3kdOOFMoADtxm05V41DTuhM8MNzezTa0OPJ8hdyZINxP8K
qcW1bSEsHRa71YX9bsjUZ1VAlamJ3cstQ7rvDH2AnyN19iw2A1DHAXh1hEuZhc+87bDKX4hKgv9z
f98XM9qBxUMT5xTNrz6cXuJtou9CYRc76+Q42E+s/GyaIyuZ+1Wn99XrRkmo9uCPe6OIZaUtQmLp
xnyopAMpXAq+cQbjQSODOSgiplWD8HqfUtVsnVAbZ2lu8k3qoI5lDsJTdSCmQIFYQIePJBC5aFjG
pYgKsyF+XxrCJUQri/2nUHTsLJx62zZo9FTWcC5EL+7QJpPXng+vSCLNHVUI651/hRgccnwkRRUq
vXTVg+JDGzvbRdwOjRGYBf9gOVETM8ofn7doAVtvfbCbRHkwiUqzHRxeTJYnvNpWFBD/nakiQ9JB
7zkQUIn/SAVINErSPhKOcow82buJekdxgw/0/F8KKrB6tMmyerB/Guz9Hf7oB7eGlVUAudSHUpFT
DCsU+P+dMB0aLoTWSnWBecnHT09Tu3OhEAls7UXOE6Cp2vvNpl4+VhuzxYOO4mB2mXw79HnYPDLs
U4geNaamWtPmavILJdPrQQPvkcnsWqkOUCyjYlw3usuWrwSGX5tWSauNUZN+7pdaB5BuW4eoT0Di
TtFt1TSm++qWy6TwXQtFJ8Sp5M2kBNGqRPSuzxtVMBNU9nEOun+4DKEhpzlhaLOkfWrlIss7/yzy
tB+d5uuNfAbQN47ALfoq6czCmDrhUCCuEuCvVV+KejQ0q/d/ZMps1UGrttBKhXLVG2GY+HAVhhlG
hkDd4yqrklwHx791+O8RvTfD4UqoFsn76Ym6ZP+BeXZkhPlF+WOYhwh+1PNRrXaIP/oeYI/2Diep
Ogxr7gut/hmsKHO0JhRWaDiAiaAxCPNkbUrFCgbXpT7qKD8q+NXOHMlxbmbtQ0Wb3BMfPecKLZzE
4dhGleL+4OvpJOuLAtqEGt8Bpqc2pBKwfJSy6vyvQCDGMEIVxKNHnmazwD8VlVhxbCEmutXNQDK1
2du7OG16ZKhROVlVM/rwlO3//jR4/LIhpgXZi+kYScE9Nsno4+YFPRyOf+PWRguvs89X2F3l5gx5
F3favH0G9UhTUm0egiaYl6/3jglW6vyud2BER+75vEStOtnZAhQ4BeGQc2GlhuqFXSiBfn4IQys2
KCjrCW80qw8rHgmFUmkZoImPUnRau3xM3OShhx1+J7BsYD4obWjBZ7Ab++UYFk1auMsf/1Y2BomC
T5QOE0uFU5xVupFYzR02X0fqFPge+j1RXG398Fg8p58OIfqisSM92AyE59NNW/sCKTLf1Ia85xI3
9nfM5TUo+ZL3OXK31BzFmxalEec2JP9JeBJa0IJrrXlf6QbS61bJX9Sj4iLmK5Bm6Q/D5am6VTNu
/HJsxKg9KFYuMSXGfiAI0O2Zu+KSn/4z7xdiFRNacuEFRL3JJdR8ciNnr/8tRfCy+4bmb6cfHtF4
c/mkMApJWboZWbjwBqXmnPzAzQUsFihzXiVfRP5ba7Mks8R+VBEqUK49UjwBIdowxgE/OYglQJvb
IonsqocvwoeOmp4nBrpzbsh3LjJhKCNMxIqwBWjti3I9KTt1BpQ0T94i5b9R1wWJTtE/W5tWXqIO
/OxiU7bS/4T4ATQ/lQRJGnT+h659SBCCMNvp8sowl20HedOaBTOl+ODiTC2KBXA4clq2CzgF1MNx
12D/0PO4n7B2/y1B8VtunFHiVtaWU5x4aJpacK2YzAubj55k3K7d4EFgBb7m54ujZhbqrz0W89rp
7NvkgtD3V358j7+cdYN2IvIK9onU+FAGot1spfV2MgM3gbyU1fsyTvLU4ANqVw0SAvyiTanG3cBr
FnypGBfJw5gt25iHkWY5VraDmQJk5XdxM3VEGRA27d8Oix+Em9tjaizk9GDJx6gkhDru4QX9qxnj
jnkWcXyis4U6K44+qHmqCvDpDNqMbXdqZVFxDqaND3eHNv6X4GGRck21rIedGXOZ6IE7HeTMOKDl
W9h63ohyorYd3iQvbx5ItTDj+pJI9dgWqjuwH/t16Ozu8VJUZxFxbmwmghG6inWelfea6E3d4OAr
8VQ1MO9ACSF8K91Nlc+OWr32F9JL9c1YSZeXymaN1kjqzCHYTxSP4Fvqv1iN5tk69TbcJF3dPUEN
xj8iqStTJLEevbDyy6E3Fwp992d3SjmQH3DK+elDYbC43kFYZQY9ipYPj1bSiMdWLFAZ0IQVer1e
Wqstv/xKzH3rS3/OuKBZNVZspEZGqNUWRoTCSh5jCK3hIexRjb0fRc+PHdQJSsxXCRmow8/h8/bu
JhO3cOouuBu3819X15PPGY8LzwF0zKK7UP8mBMszdTMe0uNWbqozklWy6YcJ6gevNePS3ryq+UUs
QCORTTdr3fcMWvqJCD2DqKihRxHkgue1MBxI64Jym8tB+lzsqOTY3ZLMgXkunOkpipxVMK4KNlqC
dwOgyOII9tTbcayWAKMx+b/26GBf0D+GNjdtNImRf7QjmI/VXhfNTFzkRxbJ4Cgf7JMwHd7EpZf7
TtaFRleFFUkKFQkurcVG66SMhaqu6HCIp+c/oy0t7cXFJxf7Hd+qcof1yobByy+oeA8uuZyJo9VL
K+ykLcjJNkRB3/Aez0wY5ISu1Dj8s2FYZjHS872haIGPsOSXydEmg7FjpXNG5Vys/ekF5EQshhaW
kqhMvOfo9sQgR3EydWfDZaBDP0HBEssXRv/eeIb9L3C2MeK5wuXVQMHBMZ8Lnior/wvJvToyxdeN
4JMhBARKHl7UzDiqOQ40U4XuPczU/VposJTIcdFTXy/9BBOGMNf6CWu26T7UH8Af+0uT/7ZRaX7g
jSZJImlJrRzZUGCC4nEXhbToQiyEGurNFDqA9nmmxasAnsHO4ZDaqnGPEr+9VMJgZw4TbZ427Inc
JnEW6VDoQLMCjJwyS8gPQ7g6G8mELrEyQziwpz5xJw8kghDVXDk9eKIiR76qXSvBWTf7VqFLiptd
393s/WnyxKwM3dP1AwGy9TGG4QFnBwioak6NC1DgADM5ei6//3lly6evebnvWHllu2symT0F13/F
ZypMl6l5oigJoMJwSUeo5Xt9Kj35UQao3fyzx4VOdKfxybJSmIdgsdTGd/tAswWNELtYLkN6U2+l
lgkYORWjz0zovBU3njcSCgW/PvFij+6UpkTAGl2qZugpeRivpVp5aMdfJ18aDqjt4QN+NyQ4QqVZ
mAWmIpdlW2k7VfOOY7zixoG2WeSnoml0tO83yziLVZp8QLeovDuB2FdtpUj+3SynY9PZ8658VoBL
O3DLM8jgFHd2du/BBZkiPLOO1lf9uB++uxJk+jdk6wGhELoAA+3M+aJ7qS5I42O+oxNTWE22XI0w
vM4f6tx0+CF76Q0mIGzFf78l90AqQFTj8ZpEVox7gVS04Eo4VJr1NOakRNRWOsSgEXsFuto2Ro9y
ErD2mY80GVnDjOFezFdYOyQlf6QE4DQ/KJhByWhd9BqCbq4NprInDB9j5+5GZzB9h6lJ0+ygdhrh
pZbRM0tp9EBwXElcm5YfHow9Cz3T/onp3n1AGzw4wMWZ6TRhCNDL2bSQuev/snk/pgPbPl3MiLjv
YvorK66rtV9L5swjwseIFFuIiM94S6H3IgApLK1sdo3JeWiQtTYGD/Vfzrb8as6KfEelxxXxJEsU
ciAe4UhZYui75tAf4kH62ChnRxgJJOvufeV630IVOS1tzkDs7GUTW4kEKbbROqSZX6lqY+FKgIAZ
7Ds7EYzGeET3JtikOdNRbgW/s96b2Z5KF0eZgRujeGaerQC+LaAeF0oOpd7lY9l0UKhLTbUNA0+z
1l62dON4oD4x0H04cVehvItg3Dgrs8EaL5QXm8og+JDBogOiEyOHy0Vu+1W/VT61utpQ87GDdvrm
VkvgRhpWI5l3ABvxDRMb1usxa05wQPE8F7ovC+VFi3LJ8OxBN0E5XWr8RYsSI9sQ+fFpSVZfXPRx
4Uv9Axl0WQGoBhzJ+a9LAHQqMVX2j+ShfcWKsBu/URrzHkFagEdV/CdqyG7YsXx0qg1PqQ93DVVH
1lkdvaVn57QpNif1uekDB8/mo7NbLy9S1XfQXZME+n4CwyB+LB+2uox0qND0zMc/RhxGOJqlu6fK
9tmt3ufBSFt6fnP/vWG+RHnznkUI0Td5XuvrZYox7ek1b5qjIg2EyviyxlaMdta1wkc1XTUXbd51
KMIRnkenhKE6q6EuG7HtPO7Z7KxPioErO2zQXd3RL3hCR2WdXfEb5nwJRN4LIYHTrkAAgG8w7MYc
CbhTiOkEfxRwQvbQrpixgvtG0DsI5TDK2fd28mIH4um3TaoOCLogufJ6vck89aRO/kKy8dM83ZAG
JVagpyxDZ7FPmWyvq5kSUJJcW6fMuT3lBp1E6w7Kx/haajMC+O3Wmm9diPgyPkwX9Qi499Uyzu7N
Qf3qe9IEXf77wFG8epxk1hWbwSZ+Dm1edaH88e/OeV3505cV3NhVuqa6CpJS53nlRKMzlUyGOalL
rWvRqfSpZlaqWNtcoa01OZM9l9immrswtOwT/v0nHhZFTY3OSlKHp7w0C+b5qiKFeg+xmN7TPOxI
Jooi/wJVRwtj404HBNqtMm4jncvwlkhdhHeDQdgPaoWkw+j7IRaYegz3xQELk3BAwArZrk3xHxZ8
Lscn/qjOzG1AlBb6bBZsunEJN/zRqspS4iKVnXOCj3HSXmdpSzjbzMa+w2qzIZRfTBjcOXTWmkIZ
nYd51YICYMnglOqFGU+iag4WlsfIhDkBM6/tW6pRCsHQuPYx+43vBmZhri2/zdtRaHEs5BRY5VTm
s13rRkTC6HTmhikX7hRQsXMPHNH67KGzwBzkitsmkiyLgI7X9pA8rrDKyleKwwX3uR6hwh2iHAcE
94nWU149KNa7jCZ/sV3Z1GRk9Vf44qx9JCTa2Mx/+/I/xvt/weJpAaxXCeKnpq6Ui72NO09W32he
Lxci0ehs1nLdn5hFhulcZnZK+SERdvjWJIWKs/GQHX6RTUzo/XZPfXDvb5BtJ+U8d8Cu8W912n1S
pXjI/ZP++cay/zZf0HCnfg81cmjlKVXxa8HuFC48xuucsbbzNaLreiLU0gdM/sMxF3zx7hDhrD0z
RMtaDm/Bg0qbvbmgRZmmHIx19gTvLKEAYJm2i/fAhhMROyGN+8wUmhuwWMYCsAOUwkgAwh736krz
9HweE1PeB4RPn9pDFv9ZqqBWwImUH2g5kAlpd75kZbBqEppa9H050xk1tJVv9RaMc9vsFsbBZLUc
vCc36Qmk/KCWx9AN6yaEr+V3FQWZle0pyQtaXTL38lbRnxFFwgT4C7Xm1RWt2j0wPIqeTrR9OIjZ
l6I5rVkps4RuuuxcuJfKMCpnjfqi+L9f9niE0vEPK7PCruxrwWD1mcdauRX+J16e5f8KfISz1W7q
6swJEvrGgQik2NA7IP2ts+62S5aXKAlHs8uPyUHWHmrtY7uQLYltJoE/wQ2fj3ouNloB5Kc8flsJ
1xm8pvJ6PBuGad4ygr60P9t16nDckWcIReOh3oCy3lzRKuOiJqrgi6ht8WfQ0mdQPaPY2X1jaUlk
eDEmi+Y8KfxPK0CGg3TBitCqyIU6IlHjDdy96bJn28az2Sahg8Gjf4vFhW8bgNtF0g4bNg44ZVpW
ZQg2vIvlP6XHlI8sz+a8ORQnDBmGX7pM/5kjOBwMSTHDrvKqDSrvZZn+zQ0xjm23OyuZJGWKls8O
9fMf4PtHo50EbE2WwbwfHAw7zAUbf7PxHIAr02FALA0fmvAXlZdRwEQD1y6tA7qeoQPnJQ9ib40W
auz9T2Jc2qK/GBBfvOF2VGWk5v6lOGTIS168Ot62c0VaJzdatsqNkWJ6nlBYiNmGDPpH4sQckRAu
gp3mDNY+7y5hvJ6kl2YrfneLfSlwCmcwxrigwAV3jT5jVJHm6b9LLt5EQk0tcj/C/MiqQ8e7yoKL
axnUkIfhSyzr3tzlD0VoLFGGfiHAM3ytioDHUATC+YForGf9fLIFIc93PlESsfnQ16fDEMB87OMo
FWXg9/+hG2HhJ6EWVIcMUTNoPeEXkS4iVlHLsNsd+JOVmLedZYFbo0W2nRgWUj07NjAHJKA7qKdK
aXkj9nGIHIeM6cdV0kYxPQWWRRIXkyinWWEHqOLqRtpTPPhHscpjMqE1inEu1R2LMhD0M65VLipZ
zSAwvv5+7pRZQivjLBT8WTXQYGuSyxnlxlpZybNOJFvSypS0PrgerImqXjrju6BkC7Iru5SD/Ait
FqwVmkn1GcdgMJj9ZM+3cNbvo2XkEHtnWZc8OR+vnpoWOjWeZh/d5jRMk3g4msTwTIf4n7ophWko
5vkwf0Zvbfgq7SLMLaBjbrBh1I0i36lu+CwxKdrNFC7r+CeH+qg7BizYRJvuTYjdx3lpgcWCjIsU
rUOvNiT3+BCVR3Tylq+/4GzUM5kLiVYxV4qg3/QCsUF567vAWqHh3H2xsrJplWJwthJuunjC6vNV
uez3i2IxfhGkXiEJuhxDZf07U+qPieo4pJ0afbUK4ii0cQki9savvjt/9w6ulcEmsiu1+P254FDk
b4f1p3c5pqvky1mMnh6h/Kg1E0TVrJ0qX4RdWmLjhRmgzgfXuWZzZJ1I0Ndz6bFLy/9uflk2y91Y
kfA4DsMQbH42bcxyZBb4D03I+GfY4jsDEILnusUTk2kRc/HVXGsCruL5aK7ITOBqGsANauURytaD
xGEwEKY1W7vhpxTlgjKu62oSb9EuGG6VViROMsquMNy4a3mTP9JnsOowIjYYUJ/vlbuqJ8WZQK1U
f9CrtCWM2xuzAr4JFJQxslT+vXVbBCtmL9CuvGO2TkdCdJ1i9rr0mOUCGPoU0h2AnnLY001MAxQC
hgPHVyHsCj54LteNXTHluVrk3K47d8v81vSno3CO11xjFW4aL8sQMd6UEtmMq02iJL/48P1FUJCP
6LS2EGQS11DGOSKTg7bgww+zXTCU8hXGHzjqP8B7MY0at1bVrKp9xm/lA/1FZEL8F4Rnu89NpAtw
5bOvslDG7ATVhMlC02UlcO8pTmzacR01d2lf5Vu346FkbEyuw6ljr8TYABQlB97nG7ViOaueMlaq
3zzghFyoU2WTJ3Kb88OOnL/zrNEj84fRYaszHT/fAZp8tawRRhFo/Za7WKobXiRQDh3gpju2OoFe
wwCvh5a/kOSctl0nEGUFyLdvAyBqjwpfEBPcGeA25bURJS8ud0zuLeBEDnvvm86oujYHSZ3suSMi
ijz1+qwc5C82qJHSX1zcPWQjyqOJJNqANnaQqyWxy8YWz71qvE6v8i88SpCcXg5/dpjzPFY2LEfi
C2M38vbtRZAyRwwCeuGjodtX58s1bT2IAUEmBeKK2POCzndqdPt94kSYF85KK20ZvU/FSpift3DP
bZRgwhz5jSFdRM18rXkWtSW6/+UHLCwTnDNEn91F07mLPYUgL7Zv5lxx1rI5ComEvJ8ERDGtO9sO
RGnsv1AvOV+LkbwKRHiKwnVfsylebb6RToGFOR1AZgmHiGS2k/g3898LFfZnJNFK9M/qVH+claXD
wmf9uPJUqdK0SRMCzaqxQcabTsUhN+jnlLBQ1BBWvsta62qkMIugpiDIWLMD1eDdZUINjYjg5I2j
/OZaEgxu5Oi4NoFTIzuXXQvKnGEB+pAr25UX/XTrDmhS7M5Qb26n9baUckvtjOykqXZrPxhP37CL
tIhyn9Uo1RZQO1a0vwRY5qTfbiU+LfoqjuKWjdNZwUJ/XOYIoqt+00/v5B+ub+/OMg89ch5/I+0t
LV4pTv/mcdhewdkSwsiLaxSkQR1srUdcD6e+TE5EySDCnWLE775EhJmCS+J3KQYdCr9A/n4V6b4J
rwFwSZIKT1DSaQJ/CfgGWS3h/m9lYh9EktiMNUmkmH1KO7Mhpt/hFHXYBlV0EuxekoHrBzgVjJd0
kCMRkwE36OVwKG2Qe1+DBBnLHl3zVkD/65A/zWgefPqCT5Cqoxw2oZZgFxftKJUFa3Z3TuuJjNG3
2ZYU8qmEtiGlD7qoibJFkrBMw8Mcw+fSYgKbvqQBmG+xufUVJwGi7nWSqH4QWRmxVwZ00rbdB5O7
yjBFYeA7nYCioC7aRLLqCDs6xRLwgk8jDixPjenI4/VPgoUvuW+28db9ytXhgFftnAdr2a6lleOo
EV5CksvEID6P2606WB2fnlIBSIu0nVgfFWUfzFAtv00yoA7v1/G2kMIigVmKfksIbV56uLaEQHDk
0roYT6L5GVn9mAwGjqXOjbK8Z9CoFOwSyd4k2cRZ6OIgbswtK+M+r1JMaTycsA7JgtAxGMby7XdH
Rsi5Hx5n5XYgJ3dhcllprVT673/wuTRE1seMj4LxpTfQpOfyD4ky4fXc+7FabdP07dSfn/MAu2om
JFq3F6YZO0L/F/I4Y9TbgYfAXTqM3sXYq5Kdym0TfYtFyJOpINlRJVGhpUkRgcnm77cgj47e9tmN
Emr2xmePNgxzymdQr/nzfssSvbZglT2G4YqEeST8pwXQA8v2nJjQlqK2y/noz8IPRi49FjhqgZbR
bgIVU9TBTlvSzaxb/YRikKTHC7hSrGPXsKk/0CAIRps+tAe329AX/NorbPweaULxZ6mIHevgytHK
M3/is7VRG7lRHx7uTcD6U15jTLp25Q7wGXvhMEqWNM0Suer5MI3ljpjCDMctxx3gX7YxMC5r9QN+
w4jG0sEtaZPPm3T1NDwjgxK/Y8U6LRGiop+0ASIXSzcy+o+QXYVcpPs2MfHeFW6NIM8TjYck6HUX
u+IgfIfWGg+WhXKYXQXijpApkYUWqS5KKGI8Ll/Cbpd4qW46gQyk61O71Zxf8fiDEXw2ECgZH0VV
JcOVh8FsQheaFa4m64O2hYYjqjJuFQERkf9L3VXKWpuTNzwH6+xOU7+0Cbqx4gYAStnB34pllfAT
tWO5D0fi4WFKeFligJB1msFlu+peJFdWOIPQwKBvSo3AiLLh11x0PaMflcuMXTj9x41/hdU6Bdz+
CmvCfezZn29Er6TduNK3xA5QLS3yeg4RFT+mBZaQoOk8fw1hZHVflOLfQUsQzyh5etwGsoeJtvKK
LSW3lk/utAg1jXrXOliL08IAI3S2FyNHesfrH1tHVLvRDik95PL/vse/bXKQm3oMY6s9w6kHbESC
abXK4TH9GTqSSfnww1h2BTxTYeY1+uAGlO/ogZwUPSHGSMmySzP/A2caP3TD+XKFysv4cDwqnr9n
djONLQZNjDjUnQm5GDblBEmwZMmaUC5l3a6Kiw8lz2FU9ns7nZqWJWC+0gAfZhKofp7axfmUG3xL
D8385C3uMC8YE2GwPwFLzaNePvSHLWEEllTLYLGGRLECQm5Um+jAjhMwCM/2TuM7gFZNA8hesCyK
fWmtkqzCSfP4sy8qak/SKbmdPj+qxpgT9nrz6AzHNTO68WGtHevymPQchaiVAtQBIXu7AP8XZN38
DaT8gKvGcgPCJE/MQsNV+0Bs5zfVRZ2mklemiUvSPb0ZW1v3NBn9SBtD+bY2Hiqabub2hPBkSz3b
5k4AJxPKGfYarOgG2YznM0a5Y9HZcHVpYmfniCN7foHfU91jvoAaTCbxZexcGmDyneqJYgAhuAQQ
vtEfF9C1erShew3O0KrTAJJZPlqsuY1xft3oTslavlunAVwFmA7Ho1WT4CE1n9atWvn5aqinD1TS
7FLA2QuIzEWjZItyElUVr06ge7ZK4EthsWZVNfpeB35YRD7zthNbchGvKL26LWZgjT6l4ybpVlHB
/ZzKucjaCCaTsDk7XG1DOZHRYgjLUB6PWnfW7S5y1xzZK7x6Ppa8GuyNgDWLXKe6PGO3OrBvsgXy
4na+WCtm33Q82ZUmiW95OcI6kKNFuiXFUCY7MA60L2CNEah5FWqk7E9IU+wKTkgfaw4VLg5vC2Z3
eAhBXW7w5b2ZMNclsPQcie0/o+YSUPTvKvL6h1CR8j0fC3k3P+EdcWFTIldz6cxaia2sahJm2Sq8
Lo2RFvXBan8GFhj9wG4ojuBOGgckNM2W7MBx/f9Xj/HaLDd21oGv0oI3+k/EzDzvjAydZNP9PKec
Y4k2Zei5T1FTW/ze9FfS7uKEeFmQAnCabX9zBEXxDCB2qYB95fbUX5xb94L7M409HeKNnXbraz8/
Jh1dgXHL8Np5KhKKzPL41S940n9POp2IygltmHt3RhVsdtntnI/reodXPOXnygNkauiNgEfiA7O9
jMJbP0hR0rhnoBliwIhOd2LxQtPgQehEaDYAoDtVGAJ+PT7VqCHeB0iWn8yRgwzLMCRGRP6PecHq
ZDDfoD1P6zbkk64BkRRelWOMUci4sUgmyfUwsmptJCk6fuf1aptPkiYa7y9edXFUmT2jq7RFbrj6
UzKcgKL6F1zH3pyvL9wVLRubRp1O2PEvDKR8a02Vv3hDXqa5+Gh0erUaRAmKcS5eGzFESFaX+54c
7noxOgWdjtMj7c2W1ULkXYPywskafG9BUo5u/+v9g89GVQ3f6Zj3mcyvC8ZHrIZNmksg2cEC8l37
42EGzLo618RpxDV3+9+zDVAm1X8QjUhW9VJlccTG/wSWdL9gNOrHOEIXB9ibqzYTEO4Z8aMyKwQD
KVsSQd2faxmdmdx3dWMAV0nK1MAHbI42cLsloL+el8P7iTGjFZM4jlQPGdvcUaAGnLTpL1l/u5j2
JWXM1LvBOcnYrrUv13bMCTia6q8X5zVd2BT1RP4JvWmC6vDQomo0W4KueFOBGXL0qcggLfUBffup
hZbothgVpweES8jrx0DGIkTITAQsxMOu7jmvxOgcQ3Ad6DCFlne24T8OFHW8R0HwrO3MR9saHeEe
yt5qJhkGbVov3bjc+CnYBuJIMMWqZjx4zJVBYpQmbee0u7VYxNsSiKPk//FHaHfkX8kKV8NAx12R
E0gW5uRcyNITMAIwHl92KjrKsfRV7wjDgI/QeMcNWkOnZ84LGE9cmy6+i6ydxM0bFhBwRH9eh2ym
Xzj4JjS0nruCsi7zJYgwr/huQIk/bePa8inmqQnERK9fEoQYhfFbJCKVf1aDCQ00nyvIeUmKaTNa
eZXg4EeR6XSpWdrHO4EdYAuUxIe/m/VDTwOs6YM0D22MqLsEgSsMxBsZM46aFrRIskejs6zlqZwA
iwwA75488ItSSB1lJSkOl5Wm+7b9EW6qY5koRX1ObOYXJhdcxXuIpNkkRCr9i/t5pX/rm7VGdl9I
cgxeAmiwiHvzgkYdWS4qm0s+zv9ndkoRQBhaLyeDR4RJBYJwjsODGT/9/E7ght5fZvVhfqFJOUgC
LyjjGoW2SvgQHEXMtaV7jn0tpbYOXtwBEozC31gAc6G/rXn9rO0zbDP27ohYZ0/pucGbDq/AUA/0
XJR0YMIhundbPCRWAnU7o8QoZ75psPF3mZyerRRb+5BuhK4bQzWXOwwkFnyMapZqsL/kZmrQB8rW
40xphQbpbj6vuhPbJAjJproiPwXVFvIfzLAFGrTeFmp6w2BzupX0YTgI0RCVn7t4t9XrfKWey9l4
IN1V120GwSDYo2C/Zw4Dh/2q1W8WTMNm7szXX/sL0Bnwr1tc6jY6BgIS7oQh6b15dM8SIXFXQn40
vUcbzvHLqEfmTBbGmA266p6pNlzSo/4Xr3NKAxYZK/kLKD4RDfo62V2IcloW52fg+y+MQxWN2d5O
QbcSb+85zyI6E7K8UXN2ZqkgnGDyp9KQQNC9FdTfLd/vqp4JuESc7h6PV29hFtbevAMrI0Syp/2n
uYBzp20imK0crTANf4l4ZUGVS3QwTBUS87YrOwe0cyx3MPFHIgG2lrJLddb1OMBDeCGZCQjg9evT
fYtBW4SqQ1z5ckBpbKpZ5xhXf0gEzDbWuzsmPTZYt6hwc7qiwumHLrg6+sp9xMVInMZjmvNpYWFN
Z5k5Dhyi7XZTTMgWDyeRFYxzcTmBpeOQWDKPT+V1tsAmnYtmP0wKepMfjygtlRIemiEyVdYe0e5v
LFvJlJW/5vxHSLIuJ9wW6CYQPkpARECPQDz4EYDo3NQmQEfpLJhlvgAZRQ+aCrEg7qdiLxV7i37N
rDeCAm9cKBkLB8eQbBdDSJLoNzJyrkAhUhkqBTky6FkPIeenlWUCJ3rYr4pKwYBa2hgXnwVXdxV2
/lJpG6c1X8jbWffGRkKjFo6GFHcmN5ivJf6Oc6/PB53k+l3Y1hfH5/g9hU+hWXl053ybhSkX4+Jy
2jrrp5loLtGfnUY49auuPwM8gU726IMN/AjIodWq5KpStsCTEJbzIQjAAvAw0xB6C9ZiQvRI11Ph
ApYhlZZAMUW3S6E2uK3KZ2TS1lD/nxthpyIvH7505e8SyzFXnx/2OpQxxfHIic4351ZeYX4tJKKb
9rWrKCp+mwQbaL9tRs2KXDspqBfPE6ftKQMAUfQpTn8ckO8Ha5LL4dzq/CzfcmE3uU+ps35vsmcR
jTAc4OOuj4lwmfK0nhaZNA+gGb2QbSz4uRYHSDfvb4V/LPPZaHGp2SzamOsfDaXq6iahse88oyG2
nmSVbM+EHP6IzRNnUD3CH9mqAqXW+Vmktj0HWCI1xZ8TztuON6gMH/yyqsX13oCEiB+SQKC2kVbU
46gRNi3EJK2V0Bd9cEpIB2SOrIrOX21BnRJ6MW5EHXHntQD0IMEg9kscgQKkWeUPBQ6GSY3ww4y4
VKgpJx/eJjI94SIvI6Gk/Kr1X42x+zIV7A9q9GRFmWt2tRLVLNxRZHLAA90IMr1nO/xTkpJ6TnWf
o6DtttPcefdiZeq8f2HY0mjM7EzM2aAJL2MINmPAT/PGMp8uOcr7RDzPYcYCxY3Y3zLI4BQXoHQ/
Ao4QrF9AiDYpSbybrHlvnUUM77ManxZPNQyI05zaOL3w8bJCRI5OWpUvxAT4wCVC/BReHTcXQf3l
7zuGKUqLvpsnJM8zGMeBQupHiqb4DnZYF0NNPTxPKnXfppyvJM9+RnLnC78EZyJcbPQvtEYMTgYM
Emc89+WwMuwtqwdXCF7YxrQzAiHr2CbdSPVeQqm3TAuvoftnKmpx/dWEd/0ysX9tFDmRqtSo+2mQ
7OQdivoijptJuXQ2RhtRBijB/C/FUS13jsL7yGKSonnVPdPCZzGX8Xh5fzWf6gkY5wSU+RA89lTH
URWwn/BicqOHyPDB3Z1ryEJVE5a9h+3YzQbXvLZrft/M0zERrbtRb+pb0nwm49e1hoGlmZBzUz+/
4Zv2xqSA+UmxUz8B5YC3CinEsrGJ3KDvs8s11Y4hSgtqjI7EiFf0YiducPKi3KoAvZ8DdmlbRL4L
ghFLJFz9yhNgMxH248Gzr/H57cr868czqAjHnGZFIEsVSbQ24s6whou3/1p8NaN1N2u1QCSdpTWZ
I1rA2Kh0Zcw5CvqjwCLjBKPDaVubWYupN7WKc1SkmdYttqpJMy3z5+86LIFJIBOOV35wYAJ5HWvE
Dko8EvXpzHBdeijTy0KMuoleF3SDYvBQ8XjgMwTbd+vwoSRPvWJLrUCXxxMiek7gfk32hMlewsiW
5qC9MZsGUxYBSKa9R+qx3NXCh/0D+rMn5pht38huYACqXeAsxJY3MS9B+qX01ZZPxcY0LpAsTolK
2yxrJi7Eq+8RSoNNSIZpKU0n1+QHA3lgxW9XzyRr7W/zMUrbkr/gQzIcmP8vAvB9wbFE6+5fPN/R
9M0QUw4/jcvWdAHKqVmAK/YE8YCVLSt4ayv99tb10PTT9TZYDTRXKcOoXxvAX5a+8FLegxKsO2h4
To3zF7db1XQ9qT3KYY1n1a9gLhEjZzPt7XkWdBQ6elfuM8AT+elh//w/f9bDQCk0lgWwGITdm+Wy
+U9/UGN2/u9jGPSqPoGMkVZAke4a/hS1AjfG03o1cCQ9nw+YXuGC0n87F85Mz0Xwmpa9D9wfUBZu
RPBr7WQT8Wd0U+XfBQ0eYQj2vrDKAwPhSjWk27QadwYKrZ1BkgjdoVZEb8rQ9Gh8AUukqHz9WHht
9NJBzwsIfajyeM62jStETumopl/IVNNEw2jKIhwsbJsmTTULc8kiAZUriq5qCivrUAo76HHx6E+g
gR+ecFmY4h14yBMtNEY4h55mMSnTe37zETVDDlLuDPttoFVsIuDXJ/ll2uMnKvsKncIt8C0ynzvm
862yHybHDT5UcPV8dFQ/vHbfA8shWy5Eyu6q4IPzoix9vdgon8kYwuf1CwTk3TwzL02ibGIuOo/M
uvahqG3YmGvOKND+xhm6JC/MWjweMCC4mwXGq/8y5lq31bZY7iPRxQXFAm1tZ+4ooIcbcGhHb1HL
iME+wSXN96ItASIgmEEe90JX+2ckP9yvHutSz8y1ZpgdA0rcr37JDCr/JTHNZRslsarc1KegkZrW
e54jHwJnOjVbCAd0aV9Z5BcdaHVdk5aULd2Nd8/t6Atgwxdwf+uTwxlpjwTcXmz0Kn/JSd0XbNDB
2hM5P6mC3WHcEytlYAuel0JR/ahGIyDX7lBuw4yQ91ncsyIZtZ9gVeynsih02dvi/xT3d9hZLQ/B
HfYKUfG3ZkSJlqFodsabhCHjjyc7kZhua5pMe2lLwXb6wba9y77sRMLgAg7IrPxsQKCrg3qEHdXX
k/rNEpVcH8LDyRyERnDYWU+foAUfEMMbmbPuaHYo+AJ2AweVIO6Ei1PVbvisZHdCLG18yj/0Rj1u
dtU87bYFwFAclPSAr+HQlp+vR7YNeIuJwfklqfwL3RGHj48DFU75NcTLRQsNzWT1V7X1UjkguQu6
Jl6SsU+FUmP9Xtcrb0LlhpC+oBQNx36gXF71yP2uncTQlAQ97947ON5iFBJDOemG+wKyTTIVlDdc
BgYQ8QSMNJzcm9b2qjcratWuyzGEBl3GjOlscuNpRI019FDEXA6Xza2DEacQlheGIfpjGN+WvHwZ
wbQchCiS9CDfEqVw9D0krvM+wHmrTAx9xgwOPyUDlozuhfJ5ZvjhTMY9kmDF7tiF7/DLEgsDUCTy
fscirJrgOdec8wYewbhTii8pklJo5diM8alT1mc2DxH3Yk9loSEMjowRq8xGAl96jUwFRdezHpD6
Zfs/GXrB1spuYtEbBsUeZ/qR+7KAysTwQooExQ00n2QHO3+GJTAFKLOAZ2luqKpJvg48Xb3Zt8Hj
de1nAFDBbkuY6pRVQiueDhNknMKWiSXd5clSEURNdRK6BILTUfXdWB63PDPjEKHEV1Nxxyk1xSFC
xR9749dffwyzN2bOLYX/YNg5jKxxCzRYW3/8HgbaLmAoMuXex4V8nwoSzN8YQ6s09gWRIF4jp2Fe
6+ojoC0EXnFeNktS7amxL/QsHEBn+RXRN9oDaJQRpKSG1tIGgo4eCzTkAeJgiTGM7c14igA8zZrO
y693zuvW9J8DNoTm4OZa5NvWfmcVrhu5cA4ZJONz4NLA/cokSpvLxOBY/4dwgVwjiFsQ+3vDVYYo
sTLY5Q1Mo0bSU3u9dAkvt5bOOQOOum3bs/7e5/0m3ld0CurMMTwn/iAKCkajBx9Mj+hcPnhAwy0E
720asxPS7fJ+Wy0uvEki6v318/JtT9/n3+hhE4iZPKUzrk104zCum7Zth5IZLYydH4M5VWyE0vzn
SvyhQVRlU7B7lulgidk26uCVIDolqD0J+uh8YYq2fpiRaCX/izh3KthlRVPtoeiHIxG0tu4V8EOl
KzPPvqWxJFwLUoL68CbBdHyy9r2jKq3WQPndJh7BvX+rieVfTS2XUcrmXe3lAAtbrAfOazSl+gY1
8Ekksm32cd4zsdA7LY+9K7/6WfCTgH3CfJLFY6SnQDXVQdNDxopFMq30BrkNqgD/cEcRphQs9BEc
jp5P0N+U9ke9GaOkfDLhBBOGWZQxPWhxU+nTJd3NYmYXsqkEzp1RVXTL3Msam6s99bex3bhUxpjk
30lBXdQb9mcAwp0ghFfLKsMmiThyBDPwvZM94WyQigX82UbCUwpfAuEq/j6KIzCuMc/TKe0aHKWe
i5aXiqJ6ckY2fCL8J2ceLNFo06ryjdpTqJCFddEQDksR6HXbWGLLzRS52b8FdaeFKS36vSLBKr8u
DhOcPIg3JG5uNFYPUemMEGWQLgpaMG6wMv9yIfhCMmCXy+c5t1DzTyBaHOZB6CtbL4xYF10XPboL
VMkM1XunQ06HxD+bHZbT4e/Czq1d+s39Aei3nCr3Akp0JSU9jP/6VyaD3g9vH+90FAlcJFsMfmk0
ezx89zzPxWL5T9uNFYQYJ8XhiFLBaPiNNrXR+rz5Li8TN9sYJ3sEX+MJTAL1hrKEYOw5lygp1vDx
l8DqIhpc/rAinUNjR+gNp20Z52kgFPEMXC94VyAa5uM0oNUAJeD5rLPoPi0AhCZgR7MlL5FinNOY
4kaerMlB548YXb+Q1DzKSURZmTBlajE7gYdcxVw2ff2JnjY/uEW1bJAnhe/yUMzTXFDtztYF2IoC
c8ynfaPmiWIm5GSpbLDYFcNVRfMCo1U/rvcB+b18CwF0TPCgeOLdkpuWbEtvhTXq8gnqXROkQy3R
9Ebqt3o10B5Nbvfqbt3l3nai5VnS33dA9FAwvT6o0DnKaBQ3gfWBp3Clm+Cuxt7HR2CyL1lBLmKe
WMosPH7aauum9vCOMmZ7n+PrBMKFT338QY+w99wL2H4JQBf/fV1NgRGKd3GObhrnom8GSHFuuIn3
M/SdQSZqAqLcu41c1ba5KfUqjqVszS/itzoSeuueAe7GC7b7PtcY1R0gPJFtvQymGTd0o6hjUr4E
XhCyVeVpvZGzo5ICk4RKfiiHjfJGkYJF2G2LyNGmIb2prCqTpnXU5lC/u1l4KZg4mX2mLi7b7k+Y
L8F43ELAoBet5H+Y8FKN223MoDcf/Rn8U3jJSYeQTF2aUNRSvWb6jDS7JtVLfElAA04TnBeT5kLj
gzIbaqNSbnqxuUnGI/ByXXwX0UPfanNPVhIFKwnWPkyaMmLoeSb3VC8Manbpqw2gDLGIPhr9r4G9
/8phwISbLCqaZTUW/rlnevJHR40XQ8Lr6rKbubMLjnw5FVEh9bT64exYl/5eQwenKNtXA8lpkUNR
Ye/W8zfymEJmfG+KYNQpjLGRos8JhJhYWd9P9AjmvbMo8bdxpHziB55zCF5S8z5a1UiwPB3tK15Q
txys4m4opk9Y4AWIbm5FjYEe28OXLAhrSPZ4z6OFMAjoq+LLoh7w+kplpibA00kK6EQwS7OOXMjt
yRbw7oNU+N5rqy3w7QVFwLSjrTHI8tzPS761yS83nOXmrAsEnNhQkH/evan/a2YqJ0kgNgXdF27E
6m/JHi/7wE27hFqddomxP1NGrMKb1taBgAlLxUkNvZ4Yu1Ch783E3YMuomXGE0dYj4QEzANcmxlw
1lm4VM1b6G+TCZAfbX5jatsv7ffqMn8quiPQrO49y4HYN4LmYgHSXx1jiOJJesozI3uk4cUYd6jO
/VxLLaTlAWNRTfAO6dbC1/fU7zynFWdnBibOpzrzLshJHXlakohbcgqpKo5PlVqmWy9ya7RNf47A
vPgFy3L2StO1yU8tg7EdxCwJIOiw+bi3z2e4JOmWnPMelVrT6AMCbctwfg+YOksbC5iJhfBsX2N4
UJgcd3ERwSU6t9tNmFRoZpLbN75lnweaHkMvIzjXwjHkZHIoEz4M9JBFypn7S792/yrMykZ7h0de
xFbm5tbU9dij12z5ElSPgjl/gbgmXwPZjjgiE7i+As3F9zqe3S28gjqnnSPus1e8YolG/QqozpV0
A9Mbxdk0JHUcLK9wIp4lY7YjpecHKzhcDxV33Gvg4ZZNLsxYTECj88Mcx0lgZ45vk/dtAWxteW7z
0jWOzzTRHDROHEXs+zJGnw+7bKzLwxrOnO0YMymHefGShtbDbemwOEL/8saWo18o2KaR8qK/9pMf
Anum1aoZdsd31JtSCJaG3F7vQEXb/h7pCzLhmpXuS0e/AV+TJv4eZinQPOQPbQ5WHjvTsMNJG+8o
O0Agdw6aVczy9gfbhD3DUmsxnXJVDjZCh9XTm8EtYWw9NWgbGmZLONYoSzS93qpkizciexFIotO9
1L9YeNLGJPGalvDBFUA/bH0fBoG5tz3mR95vQXlcIOa4VRPXc8ZZ8DxV1P4OpBhxeJcZWUzRrtuU
xfwZuOjBKz+5JnAVysw3sbsZXm/0hifzM5EWAijdL1DeRkVopwWohMz3pWDtH8bUE7YceyuIMVV/
FQYj340rVwOw6jwIB4fKqZbRa4TsyHZYWrnv6c7icvMaIbVpSN+VUucEIuMaF68GoafuqSdxBn4X
EfOHyNdfQHdXe/i599nxMHoVCyE2m4madFrKmyOvHtwMrXeJSWTnwER1wcQHckMdg3Km5azEAJpZ
516eJdlodqTFYuu9mk7eiL0ymiJtFOxDw1dU8J/lfxPnhJXVUfi6hv5ILLpg/CnjWyWQwOHpfhBo
LOUP/219AqTUNc4Su7sMQT4R5Nc4pFX3AP+l2lzHYL7stNDgbPQIqNyqaqF6mEDQrerkT7N8CB4T
3A5xwyBX8nc2cdujr4hoKGZIiVTraawd3ROoIWxH0d8anUdDCVQTrlGa/N6BPmnFnjocisqj2F+q
aG/5H9dUNkdWatIj/zWLCpMillDCXo5QHtrQ9thX5B1TbBoJpErH1XjO0xBvwH/UowmPkTS/sHWx
syfkunLaRhmsrtSpRmioez+Yi8A2ujkIoJw9P8AsXZWprcESpIP8sSviFgP9WVYMYfVPk9gSzXjU
KZx4INx5pEwGfFRjrDYU7RwiY+MLStPz0UnTwyrv21okO/S8ucxHzzqiwlcEoi2GQqaz+hWpn5f2
pzBfXvvB2DN3qucJxK1aGVsNsRh1c/9lejLjLrZlSzddfnubpIJThQ5oBDLdvd/PDhS89TA+y1bc
BdWvcm5xUEhL454K8AwhWapO0tBhW4xVZwgXl5eb5U5gNKiEfD8Iz/mB9NKZuDJL0VAt7kd/5kWf
wAsvMSKPlMykmqLFphiUQ7WoLdTePzTObFGiwIYb+aWNjvcLeu8dZMpUP0l4ugcggNMfDwUz6bwV
MB8U6ZHGxXPAFuyPeijoZe7gDzGFuRDMvb8oyfYgtJM4U5Kovf+xvM20f75p8quEeAOmjWJTo3xd
4M39YHn6ilaZ2gX9bngjZzY987X7h1MtLKkQaaaMOv5RDhmco4xNmkN8Sol5uCP7WIYhL+mdjuYx
2JMNUvjGtAvDk9G/AM+hYCBkIZljPqkbO94QubA7QFJyhqkiQE97S1tYRhGQyIqDFLJxwguM6M2x
r0slbS34fCDIO6a420369MKLF2zl4gxSp2MBqGNm3L+Z1AGu/2qkMVG65qn9K2fOWlfW3qJywSMh
0qhLTAZmIkt9B8y29JlkBQ/lud384gCNNRz2VslkhIrtuSZmuLVHCkmR/y+yj2aqhYR8SD8g1ltX
wTDnf8K+YtFixDmRk1E5HyggXOMpXuEC7ZBzePxtftg8N7u7Mijbd3pSI4rMHBp43eGoqKNbfOfz
6Eqjzllc8o6U90799FaXLFsW9zM9yXJ1y1DP693OtGi/6aWWlCPXKPUOoDBuvVMeXltskMgy0lKD
1gIq2JKUUsjR+nqQU1O0GqLtg80EGrno9x6Cg//gjnCy9c+M1u9RMukZ5PSGuT6B0zGoG6jTIsTu
6ruoECMETzxlqIAhOhZ7QyvKH6cAkepJiut1SyDBAeWx+2TvryAK21Bs589nNtUAfrM4G1xwy7BX
0Dh97U4FkZ47S+3oLopU8ylaShXFSMPvyo95BQHCKepcA8WOCGBYTBOnBpdgDpYCvE6pHOktf6s8
E2almhZQoW2222Bk/b5rW6tzagJeyQBNPjLjE7vieKLCjXCSOulUCCT2YcSx5jDJpCxMrnxhwaFL
f7akoPdk7Gh1npALaTo2e7tFXB9jjII0udsfIh6JuTK3P5HoPc+BCf3U3eaBk+Y9L6GHTdLkHmhB
5VpnDG7bT489twlz1RRGeZHUxl5v61nuDmGatg0+qSKQpJlwTVY0PjcxQXlRXW8yqlu1WIiQ3sEI
HhpoBXBCBY6RDRHyCMDKM4+2khh2d0FJXeu45WlMC199HOw3xuLllXoE2LFw61hLHZxNv/jwXVTd
HlqKVENdHl6jbiwUYLz2ASifKM6ysAfHMKboHIyYYfw7xHjWD5V5J0XvzXUUHkcuc/JrChvoR9Rr
sUNKq18Z+gty+FB4LmS5QVZRP0X7RgZGm3HuNSfAraQYJ1F7g5mNGfAKYEn6XF9creaEYO+jcS5B
0shPv9CwUPzoCU9VdpXPBWmMAoReh7WCcCdDENVIqD3MF6JLMWkV1ZjOVLJ0JX7iVPDfsYbWFJ1W
K/+eczD7jFLzZ/eKyG5bt1z+I/cyg3F1Pp/TW7i0XKuAcGkvamOelLjcQPLmtDpT/V8svY88eWtE
wqEbdHDC09K5M+URHKrJ+1ns728YpZswjvi1ad4KkeVh16DkxOgI7tI6iXUys55jCyxvXlRErFXa
lXgFiKFueAHHsYfHAjRe/eNYjd+fP9CxDFUgiQopKEs5X02R928h8TyK+OI0MDzfZHDn15mTnHm+
ZiNjI24eqwfR19Y7+UbGM8stz87aSwYHOgiRVEffJYxxZS6iHjDWiyLL0SdXXTGSn8RQdAw9vQG6
d61DHcusfWBYNsAx1bjX1RRb/JT04HNpRGDLGVmDBNvTPlEqKWABz9HM/czPds8Q93IIX+99v16M
l06qw8UvdzmftrlcUAmHSeQd4GvkzV7IIQTlXac/EPfMAb6CBUfmmV0Y2AuXkoe+dFuWozcPOOB3
Q0s5cxcn1TTSEHkaMIxSnUIEaypfqQaIdvY++ldPq74Uzn7IDUoZqtZHpM6YeypNlohFbWJNn5ox
hB/N7O2TofaplVCSwn/fTrnAY+zq0AQbJepU95Pcupg/O+dgSrwP+vBHEg3ZtuOMOxgfFPszq7Dc
ppobjNhHWLbUf+4tODF5HQtxPfwWTRCU2klh9QBYwoS8IRzgfwlNMH3xkoQVxxqo+jR8P+wCTAOz
sZDTKcf5Q69a9/K19QUJ7m8fq4mWpJRgu2k045xJ3RJygt9ZXR45KL1QHHNaf4PBdY6cxUQEt+CJ
a6XvkpAP8GHrPiZ4h9EoqXPIxbE5YkCB6H7fBTKOvnpYze32qbtP6x6tFaAWppGRs3N33FGNfB7b
8gDzC4byhSCs/cEFUiuKdwBq+/otBvrbS8cOzslQXyiXbcWVfoyvfM5ceWpPOCHb/1r/4MXMj1Fc
1NzCIeviAnlsUIRyv6butYPE4T/7yXCKBnn0i26SCHmMIoK0tD9EaRKw4bf3N8Wh70yKbJcnSVmG
UFXJcXtuI5i6gqrDQ8r4tw+lGnBrI+ujcKzP7/dkY3hJd4iplX/7SjLXMHEG2a+boTq4dRSUzFef
eEwntn4p1apoLbqI48g20T9/2PyN68L/rOAYS0mcwNP9g6wGvBvOxO49xmUpmYndMxtU+OBU0bic
kJ9JN6bEphBS6BntLv9hATbzWTpxlV2Q7kSWNr6awvXHsRznZrwEVFb1avxiNOGQUWNdAbxBGLz/
SFXPyah9HGoJg4X+Io8P9Wm+d2opEBlZnT91ovNsj/2DfT8k+81Y1oJc2enuWEZy1S7sGkMxGG9S
cKF+Jh9e568UVDJKlYdvy5RD+wUmzv9Ne9NGQUuekTC6m77ukhBAimQSs2g0KJh0geX8NvApOa0y
5z+5kdXfwltNuC9BwuXAIGQPZ3rluyJs7M/c1leWxecV/NiEvtdiBRiH9dGoPkL14mUNU6mGXhwM
7b/r/qUOyr8BMLl5pobj3hkCfEcHJxM/+/hpBNnw346ftm1hBRmXOlPvbkD94ORSfIQTHStaEk1q
CbZScrP6rYM9fBUdS9rWrACZCdjwzgk7irERpesMOT8tfDDoqCvpfyKZ2t7omnpQP6W6R34xpWmb
bL1WVVzA+O4ybNG74QZLmZoHcbmxf3JcJeaYA8Es1RNA95Y+PGCvkpsMv6Kn0Zrgg8SpZH4eaKMu
b9Rk5bSjl8D0fkQHY7aUvJXuTT1uXKsnbLFn9utWHbO3wmMTVokk/S/k2PbWRxYfzE4TQot400CZ
ttqVW/m9Fl7GB9tJyaKy3PTU6FMoR+BohUQvy+YCrOVzIWKIkamBjtPoYWoKW7f9tYOnANvDGdeo
L5HQYXwyJjK31wk59B/5fmFObmUepFNwUhjkjZ+wy0DGTdbdeZ7WhqohopURprmIwRUP8JSZxqBC
XWUgsNHv5PnnT8RZ43Ak+NKQowBCtnJbFigoxuqMq8lt4f4d7ePrM3WS5YIYN1oN54qoiqStc13N
TWAGF7Tn+X3Q1kQsb2q3febqEH9vwzT46HORx/HbhxEo61yH4A2UvlxnW7QuXdsbJxkdNxNlK6zl
DcymvpYeFARKLFYX8V8kx9a4DliHNTeMDk0/HSFkO6Y47oIZdB9GJmeTYOdBmgMyCdkkkXsryAPG
sLyv3SaLtIfNkxDo7+thmpALVQkiYE/en9vlOTLS2CxoWcAQbbXCYVgdBy7tD9/lc08Qy1P0UeVk
bKEqeHtFaLmtdrFJjGWqgtWDXTzCzLKxLplfkVTHWg87pnW7m/yt3m7FD3yxgMRFJbbw4aDIEWCg
wnXoBuTaMtucMaPUTyLa+K0IkoHc+JljilNjKJnRnyZd8eMGH3yt/pANAnScFTGGD7hZCpV+zFDW
k8XCY/35NnYcBSLTHdRF5UUkLHD73xDoWSsJObdPBmtTes0bQVsmi+avfosIKM8RIhN3wa7kA1Vi
I2MinYHHSTiPAQwDxxFLDuagNeU2Vnl9UmVxp++dGuVLGkbgnT5S8SQHuK3hPgjeDYytGhAsKIe8
hMR1pA5IjfYkHEeAOd0WmUAOQPme031bF7NqdUFDR4hMeMB5g8apu0eO9s5b5dqJJh+Kb7uN51F9
qZZOwy4O86u+e0T1n7sNAENZnvo41Ok6g3IvsOU9o/7xd8mmEPVUhog7qDlwOsaPa8ltQOCFSqbp
Hc5Koz4nFVVwOd1ogUXE+MK2J0R7dqSt4DzdhMIUv2GPG7DqBwJ4HwfqfMnUSBbTfPdjxsD29IO+
4Qh4NZ5ia0bJo89hv3o9FG4q7uJXxSAISU948WxAdAnZfsp4MzGzjofZXvkv5qKEZhO29mqswAJm
S3FfPK64B4NV7JJDulzXLZmUI8JEDPfRGelxIt2a/O7pYXOHrPJePG8JIBe08do7WWEqtZL+sGDv
PEWN1V1PyRhcPepuKA642IBA+CJ7BKdqRXnWJusm1wWcmDwhRYFrVjQTZ5d5b/QvMOqDEaaEl/Rv
Lnrw57I/vf02xEvLGwi+cRJlcWxzMsio35+4Xku6XNVli1qhpZa30ChWiZpRXsPLzQqOO4JZDhrZ
hXSGYZjAMLgf5sIMD3rbnZMzzyP1FJuB9eMffU1N2xYhmJ+Evdq7dhRVQSJTNmBNd6qENb7clj7a
KRRATH9CYv0Kh1Az4enXdidbgo9vt6tvevR7CStGrLHjWZ9biORd3L1xIBwOdv9z2ntfqLNPDk3t
xdwRDQgYTwGv0awSbzDodlcTuG/9s+AmWxzMcWLp11brMRSkY/mCuOZNtHrKXPu9OTPaeaOJ8sra
L61hh3ba0RDA9EHcYo3YqaZfymuqCfsxt0hDe6wyZhpuRZx2Uk1WoYz1go1dez6uzfdhYJYjb+ki
CSSXXuYvwqx9PxK5G1IOMZm4po+JjwhrHUwDnx6OA7PqkdZXrEmzB2c4mn1Bw12wvcyMyc6dUAn5
XGwhu9XfURDqh71XS/pEwaw47/6KDr3t3PqriUgDhHUu2DdPY/9GqUddIH91+/kZc80tVYs6+v9p
HSqbG3Xl5vfOZBu4bdH1zBYBkE2dMx9Ny3Ly/0RxpZmr9pNO6dh+fX1R4HZVuF22qiK0CTPFBBoQ
HKMYWHOQ76HuvML50pju0x+RHA58P8KpMlW59EBIujXyKtv/ejIGcZlP04Yq0+qLmxrN8Ru8BCjm
KhBXhDyjBQYOdlZWsxxrcsBJyOG+1gga6te9d5PRU6IjJT7wJo1wyeBC4Ls272JYvpG/G6XKhHMN
1JwjhT1FwXHNzq7/N5a50xlQVPToxJ6qAQ7KeSyh7wjaGSutU0ZbkEpNLSMrP8JQV2OvbDZ8WuB5
KpnFVHEgNLsc1hOR+O8cFz1COlnrGKLVom0D82Opjpeggd/FrVo/HK/WQjWTQzRHvuzdMiF3M51Q
ZjbO/aPOlsPwDVbXmzIWlwOFPSKiVqpipwo8NhCD4mkdUlEWR09ermnvaUNn+JGnPD7YBIXsA9VX
/mNHbQLbjwey9j7eJqjNHJoVrXYfJoiX6vh8HBhbeQ0kQKDVgkSS6pQVg7CfbbRZwUULP7fL2pnQ
YBwNx26UedpTLu22Tgze8hu2U0DdqZIo3mW7bEKxG1lO0/cLq/cXJkvklzDZg7Xgr4SSjcrHYEef
ANyj68RvdUwA5l0JrVyjxcFUL5u7L/qd1zAVK/G6qxGRLNTGNz1jSWBYmUI++lAAUQa5Og9aOP6i
XTmEQTnH6Ju6pIjYJjaADz+faJKfVnjxEp2S/2dH9YLluR2MK1FRL3KzKhBtb3lY3drmQi0fnJn/
Z44ocTJAf9WhoGDNM43te726ndsSpxT2Wm0x0eDealo9TvJAaaYQA9SlZ2CarjXn76vNRRneOkDq
AxH7kd4FJhGhg1yYzW+0f60xyAK562IPn0+zbXeU7urkPvrSv9AP+LoD7hzA/J5pps/7mHjppsfj
d0s0AIdhlyOMYwEmvu7OR9XFzCb57C8pnspzSAltscZgC/FzFWSWuxpa2iftGqyDFMl8rr3bKBMN
GkleaBwgc/6JwqmTf72N0/My4nRQKV6Vr1d5NdXOgKa1nT64iayscOddXbq+bfCYaF+1HrZyuaeH
pT0Fb2pjmiMXODG9JY2NnufCR625unIs7VZUd6N2hyHHaVnz5sa3JcaE8vaWhpee0Q2dkyirEPIr
2G0KgaKnsWNmfyRUO013EOaTmfMSNBvdRGurrruuJ4J+OYnCjV8vyeB5ouneQOweRax40u3GGbSF
CxZNDYsH0Ym3u1bvAImjXOjQ7tBjV9PltlZaEAU3lSS6UCpEizwBqjjn6krERQ5HPetl/zTUl2Xz
+w3EqGteiTRrMcTMbuwbaMu/UDAqJvYV2v/K3ZhbG/qweH3vDQbVn9cmyP5mD5zxe+eAUglu2tpM
ZSL/BitTnY3MqK1Wr/rmrbbag7/FvnZS4NEskhKpsW7KE6jEms4l2PvBmU/H+gh9Bd7yMtKMbweO
w+qHjMuVC0kWPEMaUAgCm9lYLxTFMyJzNtdfosu90K4bM22ft85IgrNyEJeRVRien/H+PND0FSOk
Y4m1Bkr3nKO7w0IUa+ErB+kArHzQW6EIdkEHDClcSetAvUkj2hYqFlAKREOaNnDbr0aWjUFVDbd5
jMQKQso3ML15qEepZ6xxpFcWLPUZbMIrxKnjbKOkR3JUAYGFpcAsiycI0D9/i7Qq5+ketlVicTpY
SOG+75k2lts2peTc7Sb4G1k/ZEttAeOoNbenJc8vJfpoYmtlBkSn5hxE9cIGOwADS1H2CFB1tMSd
EwM8AnKEKSVY0/MY82TCauqpe59rtr4p0GEF91D0G6Ak5ELQHg6lxOZ4kwQuD6VKWqhxhNyCFOqZ
Jadt9+Ur+UcpNokEtww7NUvguoCl7QV6Tfb6sVsaNgOxe5yTR4Z13dlWp4cCi6GINHySZXBttdY2
YiTnERRJzl5y6h+pWp13DJNaqZQROcxJx8ieMnsEt0OveV6e0yqytlqJ71QNNOK7C/Vgp2fhDval
I6+t0eLy0nyIu13qCBHWxSj4KUO0m1PsCXFhpElOe6jzOkpX9ToMsuS3r5y459Xn0KZvv9ZQmbLv
CvvKb1Qle1CXxIqbrDLN0gmD0P8kfNsFGfln+3AyKpSGsLIugNOT/Nv6uzOxWBa//S5kZy3Kxygh
0vWfz+waGfwqicD6kX61Ltb+dzqkjwMuE3/hWaVSkPKkqAX3t3QXUSnHObSmPtAtuQd+Y7WX8Fis
sWq2UqLQ0el53MgcjZHGj1HJlZn8Ss/EhwHo5ivT8ytgkLX8ZcvizbBJxowc1vpF13WHIBTJt6Gc
K8Gk7HlJbnN8mFbxB6dwB9pckG9kHBSheLFNpZkmiUtZJhJJBnfZjjNXaf9BpVykrL5hSAC41mWf
ooSf+IhA8bIO6sf/xdaMcHEjxb+Yp7bfwMo81FvOiNGWlkqNU6Qa9oTfh9kI8rZ8GFLtmaAYgqqr
2yE7z8aK9Q6y1TWq7yescYDaK5Z5OfK7Epa4cofPdGvPRawvgHzIKAik8d4ueHQC5iGdaeIxmLxb
0mcrn7Jc9GceQdqGeV1KmI35vdJwRFyOcgRolp4Opp0lTBHGbY6gvh2w48bEFLjfUDdoiJYwLfMY
fk2tePkru7zU//n0eNN/KutwKW8zZMNz3wJEzu5BiUGEZGTZZbI+TEq5l5jFwemSJCbHvX85Y5oA
VcP1tlnic2sTYrWk++2+HkXj2Mg/WzMH9I1k8WRrOLtBOelK2z5+txLqcSnSlyBvr/EbPvuHdIlT
E99IzEzrSy6DjDyjT4zPEjoLa2GFciXEbNUL5NivmOnQPx20DjNH05m9EtynvbEAzEc6PvqGxvlA
9lcItWrLGIHslrHev/SixDPCE3WBD1xTyXYFS9VksUur3tiFA+e4pvTVQVkOeNCQ0tzoRwpZHx/c
7XfSovuT7FV68vUyWq23+eepdTZW61hJoEso1dECDgLaDoJuzGlY87jLeYdHtw5Qf2uDCCqOY0hp
whdTnfFvTFppESgOVrBfQ0CkXM/eLaLMhoqUpFSUZAz7eFkFYvnBOzLAvLvEg1qYatQYR7JcJWFa
UzriRNxE2DC7ocE7tVG0LxlfUhCmOG/t7eTSE3HM/lwXk7RknFTfXIUCYFMSQGSINB3bFOk0pj3P
oFkLsH1kZ6j2F0FINw1NE8BtHu9b+iq9UqD/N9xxnaGJXRvNxu/vdxWbGcY9Y2N6qqkIjZylBoHf
1HkWih/PysKtO1hI7buNYVihi/e8DMTFTc+UrYP+wGi2XD6qk1xfNkE2sSdG5TJ3avQsQCguPZbv
vpp2IR8Thjz+Bd1aZtHerP3lKqOtWuqlb6cu+bZHgYBS2Mehh2ZbYb0mP2dGhF55UegADxlcI3DJ
jHMjO4/f4HEN92gcVCs2+6Lgmv2neGpYC+JyI5DAUSutwB8oM2DtxBjus8spSoF+cUab4VjeZ4JM
YwOYDbjeFA7KDTmcFJMMLiGOaJcT9rpaQAH4CfP4H9pFHb718glnTSl5kb5cP4H8quHWFBIV4NFc
p9BdIxEquZItUxGREnqwaWMxtqnHaOSUbCP3VurUIOKL4hTwzUYAKrPhfYRN3tzxC5aeHt7zXRgP
Giyi1dwB3uQG16b+HPJHg8PvmEQsKtCnmA/Pm9X858fWjJlzKrmUbgrxQaV8LEVZZh6CyMLhNa4j
CflVZ62s/ZY7gZB0/usADoa8TjQlUirj71dnNegxFKyAQaKIOrfzbDYYK+2O1lA/aTn/UYpz25MJ
X0jXvK8qXqhKUb1QYQEnwsYO5GfykhBPOS/OiQF/lPkCwjTfJDq4CMWQrRLikY1zhvU5/gEyz6Wo
s+4OKRo+D4QZtUaPBgYhSMFFveXR0nugezkQMf+2EQ1XGY4gFjVLMwWVcEHwctXIisMPFXlWOLVB
Zdey6SJbDBkZVZvrKXIW14QexejLMbDConFISE1JzQidL71KP6g/MPtzOf+Ym9+L8DpljNJAuEcr
VGucVyqACP0cjvbPvaSqcsUVq+D2BYD7/DkVoYksgFukwbzcK2hhK8mnB1bJRR34L1kjD2giJz9f
Yk4uDvbuj4VGQj2fG7g+PhvgLJ7Ct8mH8qB5GvVlBGrxtzqGISNZXumZ5sq33UUdGt/xnwhiX7nt
Y0gKx9p/HbAI9ann1AkhT9i8G0t+zKiLwxsZjsCOblJbEo8IpLcQDHxJze8VewcbY7c0v4r7gN8B
RavLS0T2EdtZaIYFyHVRSSHYRLoMKt8OfDcKWqU4eWUc7pH4gem6zokMVWm4aLxaYPiYAoeNPicI
+A5KKiukRCdQSGTYPgeIdPBG/u90zkEjflu5Svr6+LatxVxNiGc0q41P3ptYDQYGTY/DGCcGisEK
Q8y4YYNHHDt5rRAolLNjYBKM6imuKYOe3JCOFm77ehzA3prNQy3gdMYY1Dx/1HBWgetQyLKOLVBY
TONwF745JQKwYuBGY707gBYIiEITHRajO6byyhzYcgM8hvpB/1z7ShdNBeGJNUfT3Z33D+xqG9Qr
NoxiJJIrUSwTnDYH6DMqfgM0mOUe2n6WPXLHmbWE+EOp1KR1bi+attb7/AxgAhW6bn4b8GfHd1AM
vaSwz4AVdQqPaZNhiBMHCVWbSKT2DIBD2QxbvbcMiznxG3qsyTa8f+zIKKmp5Au2Tu4ecQGJ4/3h
/MmJxqgFQ60dUSpk8nvTx5oIiaPxBl2ZzpIS9TdVrepFdUdexwLTVyaKxzmYzO04wV97ENhL+lph
Maxn9W1F8IXwYO5MDKY4HtRYP9IFky2zRZDOyBf4KaJ9rCgLVKvWKUgCy9/+gccHuVzIUKrQNy78
K6OSpzlKdy7T0JD0t1RmmbGzXOum8xNJnrTcKeEn3P/tGsewyMC6IBU7ydUmwqjhlwolxaej9Q3A
XNmvmd+NiMcCYxy8oUdlEKPivGzBBpcGSbjYFqCOEX1XnSGQMk0ikLGIDfSNkp79Kw8N6nUJGPXR
Het8OpTkSQoHTV6YpEmFdfcZjKPmfTXjUsMj4CDsBvDhk+kAZ1zBbsOEKxkt+H/Sy8OlutAgvYC7
olBKPB/IRhdQ/NNR72RnIlxpVNj+FOxfvBG0qZttQDi8Sxo4fCgPG0LP8Nmaluej/WlVPOL+L3SG
rsECHruyHDskCLC+QpQqgge5oaXmpQyVSWnnLsRoVZSrf4jCPtCSdNLyd9vZ0m5Ms78cp4HVfK2+
0kl+ay/KwVaFWt3yVumf/ErYhcBhttgutmh3mRX79ra0J8+Yd97TLPsVIXGe3qpDDY9HM5ZaeVb1
bRWvqGBY5iB53xYP/IvCSgluZ3al9TT0YYzSBVN5jL3c+IfO6Ax5VvpUlKHMxHfLe7lIGLmJhnMr
ly10t2VESRNh/cTSS768ozp4svrHmnYFytRXzttRhQ1BgUdJ2FhlTHptgPhcyW4IvDAsLVxOlpeF
0E7Iuw7FQq7eEcwY80QkTqbMPP1qQi4yslh2cqJLHkpQaN0SWjXJJP1lKleIiBAm1gLB2HUOgl2T
2U4Zm2YLJlKFiU0zbcsU6xaQwL9NrZuYLHlzhI5vusDXd4uLDP0MKOnj0K8mW8xMTeJ4jwG38nCi
Dub7h7b+h7orYKD7jzbmlIcGgFk9smU03DL+hWbrljzR0AWPO+xqpvKdn7ZK4N+gaJSorD9Nsg0P
xNkXTa45zLshuz3PsUaHmK74TRoSbMdPeaT4PQ5hxpHj4Q2/bc0Wn+c84jvqfluTB92gOPrb5zDa
8sVmz/TcZOUskzaTytOauRNU2Br2K+bVp3+m9uYTWgYdRLhxgXL+eJW1JyQOseUlWolxBaRDNQkK
PloCBWd0tBE0BE5Xdcm5iyvu0deU/5IyfLJJ1EsobGhkHphU6AHtpUGWuXpKr2T4LC7w9PEEQLYe
HxrM/LDFz8adXj6Ycm76sjoK4hSMmUmh4yP7RJQN91qNy3W9b9F9kOaL8ogUQUm7IuhQ4Vv+46Yr
NDUUQ2nTa1aaQW6lEL8J/zx2smmutI3XPoMxxuqlcqI9X1erx+Zl6flqNw7UaivbxEnR3oKU0Upj
IkqNFngnnnaYQNxpg9CNGu/0lEXmcPiGoRapq03N3KfNKZ8HDJe1Cpg3/CkCxUA/GLcxPbS4rB1H
tiYroCLgNnoKdgzWWGl2ZtaGLlBmksO7htyBzY4geEj/cOm/VYEWHxwlKfFXDGjb18vJy7JH5NQ2
Mqm5WEt8/NxWSEGqOT3kGiTo1FzSQLVS3KiqKlynvKPWhlWKGJQyEUwkl4369XcdZoH0fswvnKKL
rJG0Zn5/wtSLPoTysyW/DRmwKHfs6Oolz9eWsbJeK+aFGAasuEaZdvD0enzs3IDQxnkziEJJQqZZ
dgVlU+aGJuvEWNa6KBja8j6KoUwWQ/iMUCDukPFt/H3Sz5aH8B/AfgsAZRmQQcU37JCgxOnTG8JW
y6db+1NlYGb/UkC1rP284c3wU9mTZ2FI85ErxZA20q8JvGSFzEOokO3bWB8OZ/hDyt8B2IXXvF2S
U1OWC4i+uEv9JEBBcRJZB2EJaOzGfKLcBSnA/V0B6sO+6YuRKisEJ37eG2Qh0YtR0LYyhGgz0j96
N5zC/LjI40Mg4JesjXI3DDGL7Nw1HEt7E28qeXfsLzrpBFWAg69ET0HNo1QEq7KqJIk54cDMxSjc
Z4Hpyh8N39iulA1oZt4xk55slNgKH7lu8CDPKFCEOdPrrZE5cO3iQKgkOeismqYH6fDSHZkUGqT1
bkpwYK/RNTlvfJhJzFfyWCFyyjJDzUgs2n02rS6proFQ8gGa82ftvao9Y7M/Yi23zfRHjjtnIaOg
IdB9qke0PWqsVAWHVWZQq4RtU4Ml5ZIjz7P9ot0PEvH3ynX9Bmw0UE/TgMESa+nm2zrSykN/mXH1
zAUfkK7/ans/xMGEU8dqcI6e5asIlRJGOQGDCT9Wn8YK3CMPsSNoyu892ieHUYxoplMJxOChFKqG
qnfIDrg2y+IlNc/mqyRIgxd3dSvEKXNrwYYEU3Ad64nU7sn+7xRN4JFDXC9LsPv7BN9wJcCHtPw+
hgiCu8i8gVmWiVkPfgl8uVGaEONkCjLobo9NRuak2iTEsYTf82d9M3yNy+C41G3LcsRFj6i7sL++
Rf8ccS3ZX9aTe0fbxcJ5kS6IPU8XEn6TaY6iujUbCIzBQH/3zNwtoNbV8AFID2ZfSpNoOACixw1d
5DD/2NTqRoa82bHi04bLy2m1nfB6j9/wo9rSWMdvXZ9ehljkCL49uCKRKMRj+9Eopc/A7IRuc10v
hIGi++sZ4KaG9zJop9MLcgg9iilDI2EXgVmSlOR1WfAoTPwX50iJbKPbuUEClC0jpVhIE0LC28X7
MDxgB/0GC14x4Lu4RW0RqN1QIpOvl3/iN8r6NWVgDySBoR/edae+uuolVvSZ27h7L65esH9Skwwl
jCcTiUXWkuRJASVtDvylGJb6XOx33D2TFAzo2N67/LeUP4Kpl0PdpS96fGMNfsZoE6BUCVDtan/X
4n4Hhy3B6jzte7AJpLuMy3hnYc3sQ49qkKSyRy4arnxeLxxUyeX8VDwQzJEgaYfs3WPeL9HrNawc
tu+l1wzFwF/+PVev6Y4dkxpJXZlm6DO6UWDnsrwxpjb+uGJTmQEstWkDHQQl5gXsk+H6j4B46Vf8
JRhmUKzy6GZLQcLd/wDhpRgt9E4cfyQDuHDb9625LjKC/lqEI7T8my0T/iioX8bC/ikypRAIiKU/
yDPq3ApxDB8sdkwkzHsZsyP/6FJCd5S2OKpKHwKBd2uCascISawoQpmXxKJiGiwnq9A4hlMe8AMu
/2GeUmFh0V4OhOKz76ScgvlOLJcUToEEnvHCtmgwpr/W8WCF1UMET3R328upXPI5N9iLFeVfioek
Vagmk+f9/teM2m6+B3m1/OAMIS5DDJbN8H1YWmRO4yr0RQkSLuaZZ6RmvohLavpenj4I4VEWEMLT
vhrmQLOf+Zck04oTXcwjXyzFq6sa2Y9AMjHDm+LDRAdxboTzvqXOR037zjAmmC9GE/1/MpKyOmsP
BriHTBOqj/DPvE8UJ1wiYb9AR8IwdJA8ktZZBoVQGHg1BSqtwZkmIL82/Kp7NnZpEnIRiATUekqu
O/Fo9IFzowRbozaQDgqfHD58jJ/XDwqY55rdwhChIZaotExNl0+R7+sDV1j7Irj4KWdeBNPS7wTp
gZQsdPcW06bd1LTMmksZn+Qq+C2BpFzHgPHPxDpIv6Pjfgzcg2MndI5Gt7EjXtY2DA2jLJLqtiF9
y7KmXvQewX5SyTp7l3TZdDLj3T4pu9K5ZaRlrtV1n6jHzql8UuE8a1cCUio1nXJ1dh157xIsDm7K
4jCQTuU0Y+4pIjyR7jW6Stjr/iqF8aWMjpJDttdLbfj2TvxHvfO2+Y1uzih8sYYhwiIQsZ3b/4+z
Km0rBO74sUs6LcR7sAanwhYnRK+qc2UDy3Aeg5VPGeSyU8+Xd9g34O9I6Loabp/Edhz18ZWffOI9
CvTdLU6I2CHvBkPuffjEdYSpfeVrgEyjlJrNTV8ciads+fhHXq1WM0Kn9qrjexO91UucJBhOrlpZ
uENbBMXrEuOmy2xMuUJBAEZ+FyH3P2DoESFxufh4EnAXgNYzl15tje7gzlRJmZGMLNX3KFcFd25A
c2aXqJZWYLQC6ugZ4bozG3kZT18eA4KsUqIqHFFJP5g7ddlDhqmYokG16AN1s8qQdzWX5cjVixnW
RbJQ1CXBO3cb2QsPu0K9VQy4m4f596kqyD9htty0F/kY6xcw39leWK4CMnnkydsOXGps10AhIXt+
I6OVSaMdp7Z99RYO1MjRfgOhqG+1+wVMf13RejB7S22HopQPjSgXNkqHWKDVVdhTNekyLfI6DwOP
sCKDupTCVQjMGpEXYk+G+yTgBKF74SJleE5T3ZPYVM5alVOYZBHJd0dxL1WsKVA+d1LDyZG5OTJn
3xyYWu4GbTxn5AknfdKxeQrwl4gLpWrR7U9W9i1/fRmHDVNjUCe4WgaKTr7PmzryGKbQaQii7dRT
UADwSvJtSRJmz1ie6AUO61s9qrCs4S0qz0B1KdQULhO5oX+n+Pjrg6vL05E3BbTc8OthYbKfbXps
ut6j6xugn52DdrtbdJ3TZMgTv0g43WMBHm8HYvCYyZw67f8tzpulUzLjLhBT4J0nOpB6eCFAztW2
tofj1R1nFqGUkpKBouOQ2GDp7oWdIz+3vF66rocV91FJF1iQA3gYE/1pvQ/MnqzhXq8itxJjenSd
5mgwaTvHs9FITVmtEHr0USePzGwDCBIMwM8t+REExO50FFFWEI0gWL6uBannvVoVBivD80JYUoKI
kRi011QkDfdTP2g2dyx0KyQwgGfijVR1qCEnnuX1EWMj6YfG/UnGefFdDZfXpNaOVkxfr5BrkHvq
1r48Cjd12L/xXuMWgg+5vb2U0tBYyEE7k1Q7Oxlvf1T7yDknNWXqGf3XCE5OJ2yZIpieqh2eaUFl
OaOIFDP7IpZNaLRZnEc4pjdYSGPWYztB+UWbM2ZLNBDCO0VsR8H8Vv0pS94DrjwzOo3aFwyiA9pb
oLr7WKF+cE/Nm1CuvyOK8SboOgyjb1oAtMQFOqVsCr6+AoJTSmJ4i35mRblAvRXN+yPq49vyCqBQ
V7CdJSKsKsm5wc8X6Cvc0HJ9n0LfpjQQbA2lTIAD+8SBG/Abv/KlmSA3Z8omZTPklnQbqFpYM37Q
7djMLQf6osuUcex/LowV+KolGGhZDvux/DCAuT8RlQo/RCwiHImJllG1xnh4pt47fCUWagf26gTT
9/bT52yMRTS0h7vw7Sde9zUMS9TVH3fQxUvCEwFVChBYigGMAI4Qekxy5NDGXVXbVxLGRMH8wcIB
7nnYDPDYUZgjhmRP8DBNmJTV2MqMnS6NIg728yYC6B8k20vTuVa2F5YCXooC6bUkZybCHyhrs9ya
VYja/IE5JTRcTff0juaZd6tlvND92w8K3Hd4kEGsWdWcGkQGCD4ZlZQOj3sBrMjT+h2yFt5k6D/Y
SlFFDabVHtLU91n3/IXE5hzdFY9Q+vZFZGoe19lY5Bim0YMGnGmhaEZ5jAYGk7Kd7DnfHWxj+Tzg
oZZa+S74v2CctpdxlgoK2PR3Fv2iXo/stzlgAPnCEce0CqHDo2YRm++OPeiNiP6o56r/EBA6ELHk
iE9Udwu7pFeZhMA4hIsygF3AN6PUu3Ud373hYFY875I3KKNhULdoqXzIozVeUWHNBJ1SBPcUuGuY
ueazCog0JhWzkkKef0O6S1DQTrbAS5IJZH+4BvfOjocyFojN0Tw6psTIlLPnJX1aTvZXOqOYpWdo
UyE2HIQELMMtBrlYWbV915aVgqTR3jUA6Fcr5aKyeUgIrzO8skQRa4/r2AOdcS3SDdhHbtigrNhd
+B/trKhNrivuQMY91x/+sfXSlH9ukHUcJKM8EX63k7VBTLPc9dcoJYhdozuboD2qItDew5gCMos+
dBFljrPCDjVbk5NSTBtjFsTLAq2VE5Sx4jc6afwMStW1NUoWzzMVHPnvoX3Ec7Z2oh5PwsTmlSDR
lvy0yYiiPKodtiIpItlSFT3R1sFX9kXZIgOp1/fJhUhXiQsKgS44Kb4TfrA5nlCgcrVAdBbbtN0g
7UXD4yqGkD0w1UFZsRU2NVm4r9e1PHoaLiRUFaLB0Lx5vZ9bpduWwPECWi0mls3n8/x8uHXRZFD6
gRTtHUuVgalRQ9cQvGn49HmUebrHtuplwHOM13pIVqH3IOcZW5AbymRkWS2+gANSu1BJubtFQ49E
iXvTamymqvZ8otxJ6nzifOiYNeIBlbmyZ1P/FVu9Ql6s3NnNocj3Oyu1gmyOZZmhZ2fevgM3NN19
xdpbrC3eoTexE6T7yfQ0bt1WwEmiot1mscgT6Dz7+EpXcGi4TvrNIRxenaW3oCF5AcRe8SpO2oAR
6qSeC+X2tHDgWMjPI+DTFNQ/FHQJ7wZMmqrDCbxXMaJpbHafjEwI8IEZL2kAoBwCgdHtn4jHj7Nx
xgAIrgS51+tTYQ1orU1qw4EzQ+ZpPBuapybe1ef721xtAHBK5C9h44kakFYfwKjvzjOMP13xh8aC
X1UkjB4V+GgRlJ+KqmZdsRkFJhhcb1/heepSEOuqgA/X+YUJysbXvJgHps1udcivpHOXZhhCUkc4
HKM9aSI/VUEuzfkATzzdM2I2wzZ8/ex+oPUXhYMLqemH8QvIzSORTYTeA7B1Uj7Yf8VzDiIYkX81
2l5VnJmKEtdrcss8xS5+Lo5KB0hFPE37mp4xwEbf8Wse1Xsg8iuEGYflEEWlDLZblBlKqRO3X//4
w8Ls4D0V7rbaGq9+h4FZonzeZxJw3j1q+YaXOyjY53Qaz0NnRbudPllQdlw4j3bX0TJ5UvwPn58O
Zo5MDq1oDJZTSTJN8dsallSpALP8JOv3/NpB99rY7MGi+sSYPK24PO5hIjESAuvVnSz6C/NYQwFr
XtPwbQ7ogy3cQrO8eKednGtW2JKg/4ZZKOj5PdYRmytblpyLN9y71KH85Gf6pDXSVeiZBLAL6w0/
QROcu0ieeswfZCMI4jlP/xOez6Gt22IxRk5WF5ntvPH15JSmLBwxkC7Tov/CAmXcrc660VeJJTlI
cPpnTgpVi7QQGx+84UloO52b7xgqXhKOJtTfDUzzPJ7ufTavk+nw4jCUKTeHLiTNBjssKCpRm5DP
Z69Jqnlmbnh22NJcvVVXjs4mnfyq6St/uxtxji/sY1Yaj/bMdMwnsG614FNLb12OLHTSHtqMYtsK
JeCM4rRKRQFroXvkWWOAapFBUtiVTIOquDdBObdF8XX8/3AjRvV/JfnCvTJNmscZMUNZcSrkjXPx
9GhDmVrmi2sx73LOxWvmc9bJFie2Ivb866QVV91tK2je8yG1VztdX03P1mfLR63hQT22zcPjy2nV
u0ivJk/la6cequ91LB1RBkwvXIT8WaEFRD0f70lybZNnaVu1i6GlEl+RejCDr32t2TaoEX4iXXR1
I0SX000l4OM5ppo2bqqt5UCMqSfclvP/N0UKXUR/Qr7EUaFnbmeXPdmFwRzAh6GpyY+BJKLcBMji
BgKxKZYw8kjR2xLZIAQMSvlb03dCbh4YJgh6AZFNFt2qHmqPbMiTu59EUwz08i5WNM498Lngj3kC
bsSxhqa8RNmS8AsCKQ5Wv+CWups6D1klJm43tGLKK67ki0EE4DXIyDgPwAdgs708EkZsNFfpBm9a
6iU/xnfJVK4pHvzM361g7QZrtCFTKfvv4z2WGKAIh8/X5gM0IGRE5m0p+4GaZkPX4pcNyBAbnMhg
VyeboDdh3pYCM5jInAElOut9Ldi0wYoKpu+h1ZMwYfwnPJDLVuN39f1OuMErF41lK4m2yMLtVbS2
VJBkFTzKrTXXBkpQ7A9DG7bAkZ+B0L9k87CHRolb+7554s6XQ1d9UrNBbLz2qgZVzIsWogOB7GsJ
4mPARjI94z2giPTEhJmjsX7iYJRe+SymKcPwLw53DO9zbS15SYAPbSuJThgP4MRYWBMFQZTppbYQ
LmjDuTPmlnt6+12bxBU65UcC/93pNyesWvIynwMYCt8NXZEgd/O+A9QqAiuh9BFAWlJnMMyzzJiv
3dWeAiDqQrh7b1aQSiPwrWGfKDHUEUSTiBOh7iJRDAs+ddSygJunEnxBxvml/JQZzev0G0qW6UjS
quv0A9JxcHt46MVyTc3FVPxdlBAr5XBWw3M1kCoc3LoP21TeRzAlTHa/wJeiomDr23cdRc9TVwQ8
8KuOP20FDKxGdLZUBWjrsjalFYKUCQ0//lINpoMfjVl8HWq7+1mo23npkO7E3rRk0bwRduZzj3Cd
ziPu+sHGSDEO2SE2t2woUkymhZroUO1ej532xE2EoWo2qGTnTlLnIlbk7ohzQPrJoEXxZYxwCG97
xwH/8MlC+g+nbpffIrf6NsCEyLe8iUDcsgyff9YbGIkUphzEox76bAb3cPJ21cTZBXK7S0r8kD3r
6ZoG2Bc1jCGk+ZkZUwFsl5UdP0uqGpqt0v+fNkTSD+t7jX2M2KbU74k/RWRJ0j2xdx5xPNvYzuJN
LCDfR+ZliAdruxtsQAxG4YUCVfWnH6xnm/dZy9Nmct7734Yn+j0OwPzwD69EosidrqrTraWHv0mz
K3N2eQ+1UFGIyOqOGJyiMB+KF0zPU4rsVRMhJUSZxNGg7vGedGSty7oWzrYbpAFmWdniUNiMSumX
NxbNpM0lAU5Tbogety35siIfs48JmamvAUkA488Y6UoYE66/xz4nm182YiT4Uj9HArArPWOUMe3c
Gf0XWhPH3t0LvqG2qEVA/aEnHX2woh5CA57wUwp3J8+r+ZONh57h5OtKbSqXnm0mllRGOBGFg/KF
UaPLW0SFEC+7Rjr1hSAtZinL2YqE3BUwOSDd89EjoKQYupBHVT7inWnxHhlPEzPXTgZ8vAalcjLD
blVJPfHTRlMyHh1rqfV9onUcaEjA4DJe11ULvtrhonBKrQUz0Aiw/2ieflHXDjeeqjOwCSF8ilja
8Xsjm1EAb4EWRmZVugs9U7TdIlDPksoyMzBiES5PgsjHJMZUUCvWQ9dbgfiIaJW25KaBJ8U35P3t
u+pwodJg96+w80cKjj0U8yFXVXUXDINNa4WzPKderu7StBi6koKaugVY1z/tciTzJyGCEZqJ+c/M
sOvSZBbCeTe2ZXRDZTAC9VPmsmaD3/I0wkCNnnNfOfySrpBfe2m4djVNo5XPT/nl71LQRZqmAd6b
BtwgPnqzGUJzGPsX9iS7g/LllDUA1FrjkVT5hmKknK3h8Ua/8tfbc6mxNvL9gr32Y7lCWdsS7w8c
+SBlAcwDYvqdXu5MftIppjDNr4FseV6N21evTAEilfkn+x7bX+LutPYsECP21me8Xn4Bvwlg0/1P
4G6GPMg54TjvxWYycvNB9HDdVuCIK1vxoRY1cTQcbkisqNRkap8VSznaZn6C2zq08vQdjR6PVwab
8glyhIO/Nl0bgTNJ/s5JEv8Qo3mb5lE+EmB9SlaLuQMS333T6NfhjrOLxLa8Byh4xXj5ZQ79DPuz
49pdyyNAgvvEbN5r3Ldattp15tJ1QVAe4z5OxvEc4K21uhyKQORCJewby01B4XbQqIYHKOFa88HA
EN0xdgiwh5xnFvrPtYkhUnaljQfpOJrAH3VCXGy86rdEoFW8OUfGVtVlhlFsSaAEv8LlxFzvl/Y6
8hMJFWnHItmJF00iJnPBmCqrpazcElc/SnY99Wj2GZCPv0hxxNuLw2kKtIr9nhWDE+/20s5Jyy/Q
H9CZg3Hm1FjaD1t0wTz2M+i+/l3ltr9zg3OkWsWlEieYZbmIgBkB5+Gj6r15VH0wQWY0/uD05erg
04VxKllxhHiRbb9u5KgQqrOlIYcB91vOhRTIBNndKp6MetxiJA+OsXm5Gz4v408x0/+FGFxlZA3T
uOixOJAOn9S1wqQUsnCzxDHzSyXH6QFIWlbPgPoSp//8IPdKNdMguBFocgu0zt9eFaVnwPR6AJ+q
C6AQ5o3TPCNw4RpItDFtI3S+HSnAovb7J0Tiwsl3WIe6yBI7UI7gnF9SYUw3KjXBaRAjIsQO65LG
CpUQKvUVkxRb7dJeX00yxWg+B6Uq5kijoSjXEpAqpupHZyeeIADbzoUPWkRVqgNSZ/3mPLODhRC6
5kpAcfGSEUjSPx6Zp9kE4nigOc4mAwCfbvZkhdyxHExAEHZiYCOuhMuqlzu+S5h5INGKJPNGMDFI
tfcAtEQW6YbhUF4b+/PGGU7jEWfTNh3OeGn5y1Lf3d8XEi13KaVloMcFOKX6oETP+Jc1ElLap3/b
dbhkZgEvbFigyWxkCjvuYP2UYAIslMWSw1UH9jJPhUp5JdinVZUAyKY/AnVEVvi7lPFq69N3CmNn
X+sUAZW9soGaqF2BCXu+5IBGVFq6pIr1SKS3jweH4DiqgL8Pwbd6Hvvgpy30cdqsTVXKjFsOywbd
1Lco9UpvY6+OYKvFw106M0ndiTcju/XEKeFlM1C+vylRVlR2f0cgDQApxQdo98I4AIjYw6NqOREK
/4GLfdrEAdb+bPdTvJuODn1ZqWq0wdJTHXIEbE5TlbBmM3a5XbXvdGku3bo8JppGle2/XDQJcCfL
afp/gGzXZqg8pNKPplObXT/ApIHxR5Byd6GKr5o75LP/ppQhvdud1Hwsjc5mdlODeEaqv8Kl7MgR
/ij8dBSinWWoaw43RS6dlCP+KCOvn1ix3/q75T5HYAaa7Tf9WfpKn8rWgsp/n4afXNnLj7hwO3vk
vmjoOhUYJvSewtR+487Mn2/ekksPON0mVxmOVq30oq4qJtpnslYEWAVKbxJ055+C7dmrFs1r++Rh
Hmh2ED4oomR5iBvesf35a7KGoY3VP/VvALxRu4XDJTmJuWUVBo4LvP+syP6VQYFTvHAJAWc4aIUt
95DY397JPUiiCW1sQuiCDYWEJKKM2lhWuE3eGdFufY1MdPFHSQGBoFx0ioiLctBiG3OxDroFbNEN
U6VtD06Hsl36u6FGXaygjEz3b0vRorhig/Qn1VdcvXGnHIT4CDUkkQiVIBlpYEFzdFgIiHYFIMMv
zsDhdTSu6sJkWiE2+C3pzjfK9lBg1C4od9pSmwNdF7egI10Zo/bYITHNXxmW/ox1x6MqjLrGeHHH
ZOb5tmCh/fRVC713CsuWaeyj00DVBQmnAKPMnOp46xQcGe++zGABtO2OLvr7Uen71XizdIprwjNl
fBkdZBQJs18qOQAQmrU4GrV1kFhAj2bLepfs9K8pBMHjjAWnN2hRk+V6SdMy5iFca+NbXRAstyvO
wxam3QcjHIwSoyqaPelAdzQ4RvGlvK8uerr6uOEF5ojfKxXIuv9cgrPnkFrc8pYDYm+9x/EkS0Xp
m1OwCJRnRBfl5Eoz4RfeNdesBQ2Buu2VhWbO55VDmMUo+oSt+XNfitmh3oUi5L4yD1qCY8p/BTQX
Qa/zvR2q1LSHvP2I5Cqch/Uu/cLyb0Wr/PFplya8hYfog/VcMGdsiD7u5LsR6CjY/weB7m+U1MyM
KeX2N5qszL+BgitHEmvIugpvUGbreX1AzuyuKQ2lzIj2E4n9/nhWfT3ENOfilfn69eF2hGa+PTGc
baioFOCqs3U4SoqYhfZ+W62vzVXunUyNH1UUJ9CYu6DT+yIEwOePHchlUOCNmeT8+zMLtjs0cDdG
zxBu45SWXLWLhphU0+nJ7DCoqS2oJYmDx1I8KSZBkqITl5etNjVM+H+MKGkYSM9QZcwRYMkvQNqx
JI1dsqVX2U5QtUWlN8piDtUpjnKlXfUQSPnqsQz/R8j4gvZiOeneOL6krz48GuOLltPuL/isHr9n
7c3Y0PZknPcie0cjDDdu8dF7mNfP9K0CghPhA0eZG8gwFSY/DUeqnQk1++AoIyXIZNLV2Rv/2kTp
Mpff/fDX64qBidQ09ZCBzxNfrvl4R/IhIR2C4vynQ0aY0bUjvq6Cj7RoaZ6SvNv5w9lKmntIuV8Z
bkHUmdzQ2yMxPML4WWfODR4GQZEtTwZTpxxiZO8vobTACXbbJu2RqSZyVb3gqdhEZinTlszUSSrP
bwIsLuomg70Z8MX37i0uHmPH6QZX6GVmsO5LNLK+fUfz2L8q4AkHlY5mSeveauBLqBT7RsFF6nKs
bwMgTwlJp2LT/EzWpQNVKBp4H+8Eh0FD3fdRq6rvwTefsfJOVDuaDb5TjwAVpi/YtahR78Ux511A
HABqdVtitS03Mz9AzSI6X0+fUTeXT2vx6UkMoNKtttIcaoc9DRijUhZrPYr+zVCZXQrgsqngutCa
/luH6gGK3DpB1eB0U57ybB+0PA0y77/4L6mHTHgzkWQR+20Fh/Zy8+Z5j9lanXRURv0zcTs1yQ0R
pBqI1OF4W30xfBV1ziHjSEjzErD6FM6G6A54oq97AUQ6zWXyssuTqQDQCR02ZLgWn1RUmi+muP1q
wc7C7j0l5XMaWzcLvwKnVrfBV9j2eXESDAhwjwBEZBCY4KB7I8w8w+zkN/9la1cyafJ7Nk0RZ+20
9hs2f8z131YFZeWdn/gNS/xhG7PwYF+nR7V74SEsea6m7zAcAtjPtQU61fmgYwwgnR1hAjv7jKIV
yHdrjwIUsnQZefXYKA0jL/IQkEBJkvABK220dv+PJ4pbOWdeKwnRVjBD/aXfBbYqLhdKqHD/L8jQ
Vb/N1W624kWhE+SNqcgwqSJGcIcFD194WZCY1aQHqBzeYAIO856nPnDwZQV7UNw8TJkm9ZMqlG8N
dk939ITgYc2suHj9yhxgEbW+f7Z5JLq+kJPAczFSOUlOLsAOKmXHJRYE4fvf/Crf2HHRg8LOHkAF
alKCtW4HRI+JHween+/TT1vLVhrk2gjdKJ6ZBwJEth4JUBaL8X2ewWacsxI+mzdaqohj4EthWy70
oOBu3iB4kyQzGyhCxcOUTGJvxsVlDKnE5jimREhXLDzm2H6AUMlhVHs/oiYDm9oTYWvIgmmvYip9
n7E8GE00rX9Z2+qCSQA+8pvca2UM/45FhAwXhkq68NQitWZeImZFXwbiX2dkgT4fo0IWyc1qqCLw
MpKLIKrgFp16Ejh/LZd+vjgFU9Dwu1pVkioLLAEfM2w4tLkj4i3ttZoG1KBpFse/JuCykS4Tcrcx
9d+9kXpJcoMVasa1L5gIVQCjr6WZHfDhF+q6YK057NpxZeytk9TZzhns3CT/qc2HzMMO8MwWZeE/
cOExtc4mgj0mksVst55WL8mwuQoRon7DWCyujK9drkH7X5tTMzDEMv5U1xDEjvJEknttD3BYT4j0
3p9E0CGsBnu/XSGzRgyqw+KlCvi3XvxTnkGiyz0n+eLFku5tsIAGvN0STMgTafpbpaL8W5+RFZzg
sMEhAZ4AW75x9KLTsRFwKBPP3H3PAZaKTOzYFUFSYC+K1fuNGnieTlr8MC0HGHHMktnz7QFr6/WN
uum2Nv27u2UEMGdD/nw8aBY09hA8LcwIYEiSzuxH1ReZ13sGit5kn/6jIY96XKdcEkFabqeyQlY1
tzxj5+ExhsSh5JbfOP35LJbFoDrE84jSQCda80KICcGQC/uYwgIhV8AUkhIzvnG19YegjIUHsV9v
6Ct/DZOdgn4ziR0AIR8vrlYLpAyLKep2iJfI2oMaHO+fIfzyo5mzhFJJ+TL61EbKP3Kp93cqN9a1
ELIqZ1DIG5GJQb9ONG7NXCWxuN/kQZims8/m6b3pH1cj1qILddt4Rhb+U1NFxRLeVKOhfao9/2PV
a5X7PkPHDYEBGMQu9DqpQub77UHFhDzzzxh8eKyf5jA8FPHSeDST4hg4Mbp4WaGCXeo3FqJxHlRq
PvLxeiyKmzit3V+UhtbqQYE03ptD2fMfdLBRrvqy5sakZFdl4WiAwqSdOtU4z9ds7VsyrnuCMeeA
8vXcIRnMVdHTeksl9EkYhqz5J1koNZ8w2PCOhuqHlns5PDo/VW2udgy+TKH0Y4ZU8pp5pfRlCqx6
fgTd9RKm6hUqcFUopdLTzoiS5yAc9M02Kdsyw8Mo1C+cr42SlUT89lAXcEuQ44+sJcaHUBd8CY+k
IX2OoWu4BatTKksc3sgzdIFt1ir6J55/ueLkuE8XIPZlbIkRR3joM5Mxac5Tfz+t6cD8Wz+D9vQC
N4jUHdg68Nb0AgbKDMGiJqdHwSfDm4MEJncB/thp6vmyJeGlInaYEu54JREYG3nMj0W947dhTwqQ
F3gtUocN/m7BJ40KFAKdSQ2MthERSl9O1Z4zj7LWc2K/vvNQOc/hMgUvXhMxkS6aIM5AkkMZpu1+
D1qWbc6AHxs1YiZU/Q0MhejMXQ/J+CVQLDiVCSBdSY5OEu4PqidChpnWrtJiC3NdxqX0WSGyLRG5
mD5jZwUPsBC/goMJJKr/zwsNzr39Yo26a0ccYzbZgWtA8lPC+T7zvCi25e4MvEFJGTvbnEpMoGe+
UoF7QIwTNbTLxbmNYlMsEU9H6oGRn/7z6ydWOp3Q4/TI+3h7cQrnzhvN1h2K3TUEcMDP76PFyCbY
WjvAROqJ3dphLEDQ7n7RCknLzqE5fe3LecM5Ka9Sg0Z4O6TRi+bxDQOf9Cckr50hD6XoVXbziy2b
QljArCd2XD3vxIlXk1++28kXqIWkp5s/zZEYbrgk6EUwmAOBgp6xVGAwVH9xxIkQIUoFfvd5epUs
CLSEPQHSsbLg5MnU00B8b2vqGgH/CaNtgYRiDiRPzcgCjTdeeZPXg8U18dg8My8vvoh269NughzI
XE3947dw7s4n/aDnz+Y8bFEczsEnCRVQozrqQ28681PvS9vR8C/d3sSrtQ/e+Um3osmrV94dnANI
eO7ZGDGLXMRW0KLBidlCLLmrxuKMPfXut00n3Lg54tjZzou6zI6i3DlYsIIPWOo+WPfkK1GjkQ5i
oPr6Chhnoe7ujoCE78LUWE+RvSHyyyRt6Rio9lSblP05Tpm9C64sihb8OTYgn7PYKpQpZ5id8S7I
XvFl1GKH9itQB41verq++aMMJ4Uut2+dGVQXxxN+GR45BoSiMsjayVeusdJisTaC93cqYx7dCTIW
/WJ7zhDtUKR7OPtHUachhP8oYhpUZcJA5XhpSeycrsCpO1mqgzsMytvHAVCzOXnIVByjAO5w2SpV
oW0yJK5pSfIB4NLrpjiI9d2j/dBAsb7its1OaThrxD3U2guUDAquROxZl6nfUreqmhpvnM0RrPsl
7mtg6Eh+Scsma6RGoZflgd0Ctx/xEzgCkxdat9TSECpHVCRpAO1QMOKzzp3l/em5dAP4u/a48nFX
NkcELVJyR2mAJNjly2I4xZ+OJg1Ehp4U/T+xZHGkVIxCb1ryJ13GIjydcXkOvSav2kT6MseTJNfB
5bnoL0364rTfW4MPNkGqAsrKQsvfA6DjBQSBDdEVnH/FdArItAL6w1goXLRAFiEid616/cjPohC0
6U5jt+4CAjSdUoj5tQJSjS9HPz5qSjklxc7Pz6PWE2WJED/nzBbmFwGO7A5k+8Ur1keyK8mULhZD
EdAuLZT0VABMapfhg2YlNfexsOGXG6cyl6xDWNoedJOaDHa3ZAvXB08WdJ64wpyNlR5fJt2SvCUX
h1W6kxjJCbGfIXift5PtYiTSjfrL3klvTiVvPerWYElH/LkiMVgOUBkj8JoB+qAdQydnmqLtAWrs
PPeR3GgnGpThq6u8yZ3OUCiJZjXiwwcl6zi5Lbb0pLKAym+rQ3R5entE8HI4eDNBphMa7y5KZJ3g
z7kzF3DpTmvvie13jPq2D2av4q8fb2Tcj6QNWV5+qu/Zn7kdyyvQCgKjMVrGu85wYPvp26cEW2V5
t+/m/W47FHo7cUQ61nqB4+UjFNVazaOuC02UxC3Prz0GPgfgk/YsrmyZtfBCxhSTssPNwIoa5alm
eFtTTrkuxrdTZHV+4smc0Mbaj2PxxNq3YpNHV0XpHgjEkfw0Pmsf1oFaaVKHqSnzL5k3MeQrEp5p
qazfx27bAgzJ5cUtOAcL/dexLdvmb0V2Zu34FmcOOzSBCdzjNunhuMqmVZCDo4JTSAr1UTbxRVSy
9qCKQJCbMt9oBwT54jNjRO6Y5k+qa8mYLFJGwLfVwCHY5yWVDs32SlZVpqVim0CB+8fBtMm0QZaU
/9r9GxCiiZjsZRjMoo/v2iTzfMTk1ryPECVQq4jVRr2vTOuRe0+OaGzGn/RgUAAcu1kPVfXa06qM
kUlDqeVmsvKu7wYTolz1hONuhH9mJd5Gkaw3peAbjUEHV00pN3H7ethBfMWJm6KyHqj/iAzbCDP+
YLBokH47z6EpY34cMliSZjK2MR2tWjqKJ8IAwCgFD9obXp/4N3bqy58/b3F0zcTET5lx91TWMU6K
Whe6sJWZZ0ZdcB8eU9CU5xO/Rtqtc3pxZ1u0+QEiGYI+27m3kdwLzdcVuFHWXjKQRV6tf39SMeN1
kRWfCtoEdi6fvh2h4l6Az6OMTtWpP4sp8O5ysiBdbPg6disUxj/A+ggFYTEMuXXAzg43xayufdKk
CA3Q6S6sSlturd2VclZw/1aImcI1UB8zAZrBMqqbsY7R2TjCwUkPIY0l7uhJBpQG4VlyVW8VIsfi
wU3S6blqRPTRI9o4lNGqC4oi+XfAVkybIQQA0qmIgA6lFQ32yotSp2HMnBNUWNrd8P3YQ01X88Q9
Cb6PYRFvnOgDDmkV1nyKEnEpNvRxxel1BBIyHP/wooRl73aMOGEpAgO5XehktGygMS640l9b+bDv
n3tWrkat3LNXHta2gUSfN5HOLhTAiBTB4rLC1m4mPyQrCaLh6E72OokzGsVnBVkcqraRiFaCajfo
3NWArCGAOXtj6nraih6RazNhPxrTPKZFh9v9UcfTxwDSSW6OTPMV6n4dMo7OdD6Xa/1Hp7DF5J2g
L+j8SuRbvUZc/FOAHaaitrDstjwPxbxi5uMQw9IjyQJI5Mm6Bi1ZVv7UF/D3kAoa9lzSYNY/C4lh
5swwEfNnUv0/722bOUlqhjoeMAauerK0//QGoTbulnufOBCKMggAexRWgF8CLrRuvRe7eysb4PA7
7EO+57IyxBOkEh7NrOIVGMr44ZCX7ebLbpF5OHKSG6d9x6Kyvp3firqJnwKb+95RFO7yHbWGvZUA
2UCXLvP5uycCb/e9MENMZlhHXgyWmzgxqaWDC70SZ6j6iY4wPNQeMkcG7OCQ1ek3EO12hksPAUHK
fXdo+sEYXhvZw1opsB8fFpxNhar2jCp1yUzwH0nR8G4ZtRBvZLTwnbAY3zJIgE52IRsqiv/qdKxh
1rQAnE/gZrePhN/2YhltzByjU1pUz6xdzHndU18NeJxc1u5SX0rp40be/5cT9QuUpngfOdhIGCwV
DIVIFdPe+dW7OiZCBlvPJGlAG8w+fmJ2FBwKeXYIIUHSzE2wJMuEvOm2MrPDXGTOwZF43RpNP9WM
b5Ks1/RflZkRQC1oOyD7tMj/9H9rhjLlxW+oSWwPXyrO+cB96ATM7I9swX2jIBuee2xLbAsdYsrV
c1fy8oSbNfk0kprvVLrbdrtRUPVMAiRsHmp7yam9aCTmfxPFOwYCxKUogmDKfOgSdN6twxZGhVBV
HrH64P07GT+ETdn1PyUYrilVCOi2NoVkQDLTTSj1p0p1UqytYmDFEwSA+L3UJ0B9ILbCxsPupkf3
w0XDrtPyw2q7hBmiUaZRb7FwgciYPwEHroxKNaTJXqTc19IOvSoLzjOYp1hLvJxusfhu9nkAEXda
4MIY/r5Mo1dnSJNG8WXO8qPS6Zf6OkEDAZtRySWCsdDdGQApwKHOKc4Xg3+mNwcI2uuu7z1IvtkQ
kbyfSasbEZ/129KUSh/GQSdqdx+9NARou5kZzeiM5qfOUuDa5r6JDo8PH6I2vRF7Ghugm/jFLoo4
DGl74zuCIq8quHw7Rkqz0xo8jVKdkGDNVQ2PWBR53arXzV228RCW5fa7jN1za3tOPA5naZf5lFxf
+Oi6qVEjsrIdT7TbLUTStNHAesd3JtXHlVUhz7kDamM6GsyKh7nYzn0LP0K5OSTIr9ctBEa+JKep
dPDF3npmYrJhBUHy7i7ZRpNZCNlLDrQD2kW5H0aFdDyAzoGmc2Gfg6v9IDkjx7ivK7Lp8dJe+tnh
jyv+MZ5jpp3pOcMEw3E7jhdkFqvbWkx7zg6qwGgLvNBjpukYJxaf4Ezy9cgpOG19fw7fxuKSHlEp
kAI3bL3GhC4kNVYGHeMwDBOfd1MopbYLMu87SlZZ4wVK9YcJ+5NLRZvIvtaSsApVoGxavgA54yS7
hrrtozXWQ4d3qwPmyhT1dVmD88PHlkuchIGuAdqyu5OhpLrVNu3FfDHcdJBqsdSOkKKgdnr0aVxa
U0uHordDfAR7YQvrs9+B4JJIgP+iWWVlgJ0cNbkkyAsQHtH/aaXsBoLKBxVe+VRXurtWX/gyIxbo
tKuAI2EdekvGmuxia74e7zToAmRpHjeqTn3klfB+j9y9ReHNWV0NXqigBS3rqQV5CgWZl+RrS3lq
zXVOs85jZBmqG/4rOPMZN+BgobUzNRPOUUUkC0OA6tGRMdafWMit+O72hol2ytOapxn4OrtzveON
LUjfa5+Fdinhjbm5WtcfGjBJQO1t/NmXWptLR8VfgrE00taR0O+5DuFC/g1bnix1lSOmaXctPTvQ
JOc1Gs5t4hKAG1zTNlTTiQR2S2UTs1+7P8zTUiKFXmNnUMrA7TpPUC2J+bqMTAMSHZBzPSsc2roF
ooQjU9VuNs68QvOTGja+vgIbbud5VncCW1a59zCwmHxmBnAiU76bwNNTQ48aUHMqhOj2N27ANI0L
0v+hbts+Ix2JB10sk2LbJ0C4wpFtZTeFTxb19PDoYlCvRiApbeNe1a6taa0l2f+CdLvqou4sGjjr
ryYxHR7EfSjURNcASTOWX821y5l6nalmTnd1I4BNkTuSxnIrtlZjn3LaQNnZXPg7ljt7a+De9AOl
9RGqaaax/lboTgfUhRVunvdfWinKhVUt3wQweY47p6LWZVmrkVW6WO7y3L6DUAV2Td2ki+5Umm+8
OSNlRCTx+wE9CIryyi5vjeR0DSuzYC9XndiB5N0xNr1kFOahupDgfJydASG6Cn3E7Xq846zWHzUi
XdWJ2vW9+031Vb6jdYxY27andPBsE8nzaqug3S37XyK+N64AKG+xcQ7hjSga62K+6gXBEDjrw5cO
MDV83B03sFmQGLKY8uxGQ8vbHa0179FSyRRf6CuOfgMp9l6z6Zlo80BdlBjz45Kdn8BWTHSpT5NU
WVPSbf3UHydnLo5C9mZN7srtVwDwTH1xexP52TD1IBxSXevihoQl9V4rZ7r2ti9QPxUmrtuiIq1T
VemmSJXGXp211Q0nVqZ2fXOm16esALZ4RKPjKyhAH8ioPNwD+69C6RHd70NPrvdoDVKh2Y2RkihS
x7nlRdw/QQ9a5rlwjTKCwIfzDC3T+e8+YOVbAQxBtU3HtIaQsm9Q4ftsTM+C12I8BCZW5EBVUS+9
2xNTQsKjMxd7YxmKAmT9+WXJQIyuR9fCHspR0CkUfrhJrcYaVoSroQKT6H8vA34aBF6uBMx5A54O
2VQjPwuDivCFjcVEpd0USP//8zOucBkzlcOpOqVa6/ab2jEwUpwvJ2lzLPFfE6lCkVUFM+FPFyVs
IFPI/lcqey8fQQbS+MK1tkj+gL8WEX4h7nYVotaYZcnxaw1dYI59td/XahRLv/4netrvl/F3RelI
T0Avmj98H/aRyIbrWVRbH7CFq7435CksGFx8HiLQyPJuP27NtsspJuQXKYMj0cBNrTLpi15KEFzi
1VASTvevlQlfnhdYrUjfx3Y64TIX7m2vHkiKEy8hl8sBW3SS2fTTbqF8pq/tFMeAMXtUEu6djxQ9
8t+ada5hi/E3cQbf3hssBSxbQcHfcw+tSw2cfT2NlqI5CBEb2fWVvfYbplVx9sjxe+suugzT+FXb
QWFswtBsfSbYP7NO7K25scgwYgZHVoYm1iJOOntO08mUqGCMRb3f55+XsifaZIG0WTVXJ8SxB4bI
SKTu6L3lZZ2YiKDX3VF7sWKLdAEUFs6Q5Da6cyYUNJVlh91FpP1Rjm0H3k3xuUHGTJGUT+RPhTtX
Y53Z7aZ2pk11PrBZdR4sGbThY8pblt7tN7ItdgD7tKpxG1m/ZvbLwec5Nlgd4PwB45PH2hblxTLW
ZQV6J35MrA7nubavNI9mhtgDDTQbobTLn6Mbw4nijTqrEQyz4CVCl3DzdpxKRZYg5RElPu4Wqp/c
+9eDIRE+jflghzfMd/63BYzWdm1ox93hmCASBxzS/uOLaEqc+xZXjxHimIajf9iyaRFbkm1MOhKT
fFQPz17ezyNr5gcKafAWTFR9DCljw6DC6TLh4bpBBzM3EFg6zuAEMnAm1/DTNxRydT+l+KzN1eYM
sY/Q/u8LH87/kugdKbSdBkLnXkcnMeYmi9pfH1ou9p32CseiK4WORgPJ2coUrG4TV30uF/WnekrG
qz/gDqRdIMzv6Pup61dFZn65KYHXxL/hz+2D03Z7H5qOUlFk2g4LpGcPXD+cjUc7Jz+PXrJzhYY3
73U8pom+DA58t6iNewSPTJPHqPTwpREFo/qmztV8HoewM3Note6BiPeWvQwFKTJlAJGJfTxkR+VS
enscIUZNLZOhqUfwTGps71yJCsYEiqkkmrq96V8joOfG7QwkGKwcVLGLqNmKI5QWKzy2xkSPEVxi
V4Qbw+xp8Zd6ycTSgMPqrPzzkFf8OkoC8YOvfFLoAhfuwQkcLFGjiYdRWbWD6k9i/fb9PTezIfoH
d9oJqAaBev1i4TWL4q0dsIi0PtvTArHswV5og0A9sVqNJS09OHCPCDwU9GT7MqxKrCPe8OKwQM8g
IZiqE3McAf6fL/bBac+85gHFc+qY8VhWHPRodb2hwFFIpevPoZXNVp+FsFGkzMr/RWevDE5VOebF
pTrYCydBqO4ZLywVSptVwivyr5xn/dbUgkJPwa4UA451ABjgez2tFLYMt6KGMSQzN0kBOtcrirK8
UmdcRdhedUiOnwPV/XaLdITFYwgchMdJS5bqDErG2mQN7iidhNve7HuRCGSIVSkoZ7EAk+KeVYIh
wVPdbDz/qcXfEwe0lBqPtp5rQvXSyckK+6heFy5fcwPnh49ou7gvOLmcEz3Jhzi7Y3lERDUTxNuh
kElpdvAySXcp/PE65zECtxPGPxBjM7acdtNhOtvit+/+zYOdAiR62rF93zlh8phY4xPcDbc3f5Xr
YLxe71X4Oo8MRAVZRnU6EI/pCLmXueAUXpURZ2fQxx28s0RTNHYCUxPlsEcbfdb0QXZ/J3PXHeME
VC26mw3yWIrPJgYRsYTgkyM84br4CVpFx6pNfUbhr5LjTzKSjUpxrEyeb75OSn8wQcUfBl7itjWz
ABNTji4NRIJCx+ggb0YNm515dhMhM3leMUTPrcTpyiWu07PWqHE93iRT+RzV/Y/sK0G2mRoWMKij
ITqQUA6giCNA+twQhKsfa8pfS8hCODPZ0UTDyc6X3uQNTL4qhUZ82+cn6O0AG5Z0gKoop5JME3Kc
NFLoSCYGTI9AO/FYcAUAQUMkaS2dVLVKQbH2eHey766tOdfyTy/mSdWZW4qh+Y90s1MCpmjGMiNj
n5HAut85ft9eb8ESQ2t1cxA+SdLMAp+zJ+iDjDdqiJXhUl2YHXmP6K1tBhurRG1ReqijGbG1uxzm
SLCcKJgBzQBmEsxZ02V0YPEpglIn4BFPQFLiZQdQnIxG+182IXaUDBLbkQwWhnXS/JEBwTLOF1Bd
dr+pnHNVJJj7RRtEmlCKoMzPSoxnvw3AxRgYaHDdLyw6JffWJv//XKRn+ZAspKkNbIe9J9lD2Cev
ulwbeRjP4Tt4iBAaZ+uFgS6YlfC7omnGeoRZPJhgzW60PZALZNqAbhyc0xUlQfpVGKn86lOAMrT/
Zrxgd5Ns1GxWqKp4lkiFRB5mqEWF/NAiFFc4I9BifZzWCNbrqJPL4btrLNGOrNRz3b8//V+ZbRg1
ax7V+wOBjDUPpJs/bwIPbYiRM2obcXALEWozVx9muET9hVtofIXIGOH9urYhB2649SmuPQlYqgQC
rGELWg4Zqc9jdH4/ZSZ8KigOr3hyfV8tNRRySd5MBxbL1507nmwXfwiSraRnE/66H+OVqYPe+jo+
hJgnpfAgu+8qMKOqcjhj26pzOTTJIng+G4IGqkKCmtipSxA31zuzAYHOfcLv49aTXP3Ayn3y2t9l
R6xFrwhsX2TWvZJsUcRuVxsewBGPFS5agUphAd9YtLG9TkXyR/PFMd1d6btIymH27Y8DqqEN+dX9
L5zcRRCRoyEVPRRrnDRPgM8/V7mPDJRXHyyUEmtwnUNQwo8Fpewh7Y+GkqxA+TPD3Ww5HC5FM/5f
OypuNuo6KMDMdidVzbRYhJ9CabtnTKrDfWJZWvQUfvgINb4EGcnXuK9WUSTgNDKDmDrb2pb0+hw/
CxmomkEpZovkzKUFGhunPqbc0kdDd5Q65mn1Qk+aKxR+RaaBYjgTeXU1BbCERm2OMWScjUFnJ48H
LVxz9c1q3bVkpgy6jtCXxkBSLuAKlylxnE2FwbkU3RYcEwRVdruEUzqAOVJNFuku56bIAd7sVhRZ
/1T1g0Jda7onwrI3vuOSrCIZHGso/pvP3X9U92weNY0t8Rda0sythSYTgAASycxCjFGJQychDGbX
X6AXkCqMo2Ku1OlzYC23qv/bcR0DhEme8x2GIDdo0aUonjxad5y6JcuPph15ksQhTIuNzKJB/Iab
vLPjovLnBV2J2+mPVuSDZM/vwHwjHg/IlaqRF+Er/b2AR6caPg+RNvp7vLdC9qg1L+Nxfbp6RzMs
PQVBN9J02WZPxkEVYIwK3YRyUxzf2v6P6CI11j1mNBFoivESvBicwoRT+Zgy3RIDezG7LQjKZBt5
O8HURc45joVqJ6RJWLEkaPZaFkm8OuIQQKsE5UeqGshgRDeNPXh5NuSZr+ijaY183v6xC5MYzAo3
59r+IzY3TcWkVFGfi1mSlJ4F5Raqmmuh6/X2Z4XzVEKcJ1ELMbx19UgciJz1LNaO6mpJYkfDs64N
R93DEJAvxQ02CZt61qUaod0qHWzzOyFDVfkx+rStCBgJtjNEWhWtz6slio6gu4t5zAQszgNw1qAJ
oiEW05l0XRBTZn5itStigrcIaYmZ0uhcn8+18oGUYdoap2F0TTS1KUgU8UG7ys1fQs6scC99Cdco
wISdIqIpauyvSNQ2wFmhLdNIfqKsDswCcbk86FAw2ClF8biTLGjWhy7LF1SX5Jlf8EdiASby7I5a
R7GRggy6Nh4cDHvc/BPSL2pKfFTdMq/99Ipy4GnC0hUxLWKTNcYSJvF62QMRKEgcMH9huhPHlq6U
Snpsmyr6WBRNxxfVLfxVxvGnnnsBs+xG1wgr5ejLmkQ318KSXlhTEDZ6AiBQ4Ad7zYSZ0vDIpDX8
3QWP6II9Qk3EC3L79Tnz/pX/5AA4ZPZ54OPuwr9TniWDCb+/42sGtgcT/iApGHLmlZmOGG/sLeom
r49yw0dZmeWvkvdpAytsig0XLMI7dmWQr4hddv4zYEGU+N+0j2QLXK3B09E2ZTds4Z8N6tnrPGGq
7rgfRZNkRDkFTb8vpdky+Bw4ucRlCYv1V6XMr+IZDcW05VAtr1ZrpJpzgb4V0ShWVaTk+0e7LflL
5GHDqovopF+MFjO1yA3sF2hFvIq/cMEO/Xw7kAjMq1FJADe4UY9JCOfsWpl5zLl5og38OETAGrea
vydna5pEpNFCCEV3IvaZ9fp+fSEpwOM9aK4Do5lTmnAgIvdk2eSZpH1O7usmY3lnCyYd4jL/n3yt
Ua1tIhCWyxBGj4hIDOh2RnIw4AGhqj0JFKiRH+6llLDsDsFhv5j45Nmbhk8nnv3eFUZB/oxEz3YD
3EW0sFfhCN6Mu8tetje38nn19a7o1cEHwUkDiMNY2LK538fiV6SWzDNz2Lywot0BAlxl42L7spb5
6yKxx1uUbYtPOmtrc0bh/ZP2sqYA2A1Nnt0PGfnkqALBGLqh7F7aagdb4/doGpT2u/9jtoxRTkQb
0LeXhOpakaE4JfdyYvMbIIJB5sotDoUWxOzlTfCr12rPJjaPrREfd5UZ7Z3rayh+KUaKlvm0Ms3K
vOrIgf8ktpYbvpJJVVvYzFVGLdfnQW/5Pwu/49Cqa1mXr0gJbYqBfHqWD0fI6vcWFqJJ4jK+iVvR
Ur7eA1gOEAuC1c0cOfQMyFzeSBioUdjfiBwXw0qWr0CyaJ8UwzmdeOjIYabnBXZoBziIM6L6ljSz
/IFr7ifk6iSIaPLbiqodvIbRsSdT0t2mL0U+wX6k51ogCOb/CMN5yXhcbZUuGIe3K15trmo3oF3O
JSeZKDmiLF17VJUX8E0LMg1kNPFdsqtxqFNSrENOvbAEatuIhqXnvgu9K2eKJ94k7P9WOgAtj1cv
TKWx8VMV8JY8qZF9+LfD37kdKxd5dl/OL7cHNbKtYQbp4/jtsGuQf6dWcxkwfjxJVt3cpop2dRCh
aid8vyviibBMmtgk4yzkIth+gG/Y5sNv9V4aCogJor9ncgAwJevBA+3Sc/iBJwSwugSoNczSnqQy
Q2w79v0qq/5fJPyaqCE253kVZ8IEUWMcjFXH6g52njkMI0bGioaCkKU+qMNbV2z0sbZ+XbFo1+Do
M67nxWOBQT53q4lBdNEecuToCy6jSSOIHR0uH2LYp6qNkbedsVz1JtavwKDdYkCLVN90FDBJrUPj
MjsMhS/J1bN4EwRoIBdgNYbwzJdYDO8QKal/rC/n0Uim0XhWRnkHhXIAtj95HZwxkGRbAyAun+SV
42O5fArA1bKpBq9Tzo0Y4sauGVFkmL9rDWTVbPewCkKjon3i0HzD13StooP0Jo6geBp5fG1eo0F4
o+id5ZulnzYwxyvoSnmhlIYniD6gf4Csd2EYMV7OsI13uSakYbzfifAjQ8/GJaqZaaTCty0M01TV
d/mOYoZRMkiHcDqmzHtjYNNS4V0eScBjDgIQwBI6Kw5UeSeSewkS4iuVXuhy1y580vpdZ/H40+zT
ODJruFOyXxSDzcjHDfBKAPn837JeGVefJ/3/XBPngdAeg5rZhmZsrJF1P1tvfqIDxqOO3gnNP7qg
I05HVwq/Bz+Oi2RDdClPVVNSpqYwaYhQ8qLi34+jy6ikk7l/uXrf3Nl66D3O5Ls2se7k8RcGIhZR
u7ycGKHquIMtzasI+Rs3J5Y5GjXNTuQhnX4yUwYucTO1I4dUM3d7slnoAD4G/gWXptafg6H7zZ0i
7qyUMx8nur5nTssTviC5l4UbnPiZjtzTqjNXCb9NuSv7COiJtgt2a19YgTaMeQJs9oF1pLIDEEEm
DK+GjWXRv9tsnd3EpasuIPWgXE2536LQGkBDKb+r+S/AubkovLlTiWf9Ub2cQ/+WdcV/V6VgEAJn
sFl5XiO7rHAFHbfkQ2nwCcP8QxyLJB8ty3k8HIHtoc2wNy1uMjuykOTN4i+cvT1GZQxDGLTh6d+9
0BDHjz0qowwC7t4OOTHaxhaROWRBJ2QVsst2PkZPmdqiryXqCKVbROomXgbBZr6Kb5uaEE9G+be4
33mN/Syd/r/zhsZJL1MVEmCZExZxhU1GfYOQPZY3jxP5RA/eqystKn7VJaJ1R35gouEy79PRjOBY
XpRosTa0XJTUnlRjYlr4mdg4hgrgfNppO92ZgM9RMTmh5YizpoxvbZjZ/gW0+SWR199tRv2Fqcwn
wC2eteLjq+TbMbH25J3qgZz3TlNUb7H9pwqPOtfgglqVIdesXr64wGwhATlgMbvPdeCnHH5GhM9s
9Jmyuxaa6g89kELbqxC+NFbTPIBb2qfXpZO9KRZwKVDntoz96GUmU9f+LY89UN97IROmxfuSLMUP
XBT/scSlhU18xsm7pK6IBaE28KsLg7hN5OK++sGYibW1vLvYBmzF4nBce+lMxmUAthm13v19Wn0j
ruAJsrykPAlvyfkEeUn3bPiDd3kZ50R5ZBIW4V5/UQDvo+OelYTpSh+qB6tq2210XrC8xPNTKZ77
4F4i5/n+UxKYxmQLS4IhPIOhnEQ9BNfB8Rg0CYOvuqlcY3dlYJJeWC0lGYdUxktdUd12WucRsCQW
FcYC+dfszCmuwTgXeVWppig7xUNjB7DweViy24jkwpqDpoMnzBIUoZ+P1z6gcn6FP1mClKm7KqGC
/MPlprRsyDpzz95+LRk7zHDy1tV8UfOo/umFJLIl01HncuhFJsalOwtl2ijgc1oennkDRrksBsB7
66V/QoetLFgmzk6D2n6k07LBdusm0vAakPv2Fyuh6bp0Jew/CudX2ElLoMpQlz/GovD8jA5Nygop
nuay59WxYQcAd9bIYy/F0TPlEAnAgHtuw/BlNCarzpbWFHbjA2K2aiKIHgSaEyznNS5Gais7lr9n
lZBxGd4l9BFCkyPOwiXXMxb47W12yjnKYiofsXnmuHowZ6L8mbVve9eJngeuScujdSuPouN8w1Hm
KzFa4pcniWF4eVWUTeQ9e49Y051MSrRIQScxjkF8PHNlFbroozG81WaofPYJB7X6fxAeHWqj3RRI
Opn3iN+bSwAVXMeyWSVARI5vzaQHDK81trQgYAKyh3QjiRoCd72gHYHURnsLDlN+6AiwfTBu2f11
KCSKcxxQoeNP8AMRPGDfVzTqvlN9GNa0vo6A5Er+4bwoPDRcrW43z/FGphv2M5N/w81qLs5xiBSE
BY3Fbn7w50DviZUUTwZZxuRXvtRNJzVYY7sniYdWoVQey6MT4/B2wFTZmd1OFH2kgXfi4f1gp7um
cd7H81vomPPiieXc8wdAEKLxlP03f/ONyvH6gqEx5jNn3c8egzJpWtoBLKIaslWEytyvfSQipE7b
cmPLbHKIpWeYr51BhW/Ya310xNR9Wwf9vglO2VG0yXzA3QR8KtqKbR07TxORdTABpovkquScwcge
1ZlHULyg0uAjldddw9pU2EjTijPr1JTkQTq9GJhwuqTZLgZox4cvXoeE0NGuRw8ypjccZbZJ5ub+
OyKykStY9Pw5ETufL75/C6UAlC/8KGhRgBRaAZp89anDgRSY0wNB5TTcfwYtzi4CDlCL0AvUh1jJ
9cVSGvm5wtl8KLeeA2nU7AK2T/5rL6mJi8hzfpHbP6ORzqVGfpKYK3fyaQSJcdGYX6bKuAhGMVow
cijLZP5NxwgR8XWuZgvhuJj8oee6M6G5A8E/W2Pj++WraB6F6eCmAmhq7gI7e3W7CLAEjc1i0N5T
JjvuoC6cES8gJlLoplTr0l5sGbErehE7hU2FRahXA3hJPKkUbMlj2FLbfFl6AwK4BtAYu71of85f
rbP2WbkdwpAnGZ0tJoPaSSrYjU0sk4iqjWZKoIRa283ea5P7EBH9/ZGjgGtXxmyDTj14XCY3bDkj
5b+90geXpZHiQr8C+nPQ+tmYiT7wAbSOKorh79wQxDDYVEFwH5CjwG+iDnplWLsHnqjAu7UpHQR7
JOgJH8DOfDH7p1YaH5+0hJ+v8SG/T/t0NZwmdwII0YlcO49Cj/cQqRR1no1RAvt+v6sTa76nctco
Lp6sqiKIK1lzIJXgcJR6ZLbNFxppkE5ws/AB/2lb/iNDnM12FA0s9LAYD1aKQJWExufFsEHo5D0o
rVdgr43dTAqV3qJd1ciICHVCJctmSaC1PZsYFLU+hfS6raVBP7bqxiCcWuHwrtJqX4E5y9eDef+o
E2pkqfu5obkFpqBRk+FRcwMecCGHgIHljuWYOnIvAI1fW8/+JEX+v5JNx6ykm0j3t8VqZljd+BwD
D72B15An5s/LF8asQaIKev6McRS/a1NDcy37RWYMDyv8DhZxn9dFm5WERY/XDHIdOPIZaDHdDEAz
7KrECfyMfJC1dA+kCz8TiahXkt55zYR+QBa5W7by7LFytSOtk7TPqJ5REuDhCKkSkIlSiwRuv1B6
5kgU9g0IN10SEoMrmiyf7sb7jQmK1V7JNzkHKY01EJngcdUv8cDVTjOL41AuKmJCP5s4/iPZpxmQ
F4PFGBnatjikdV7C6B/HyxdhukdBJLEeNHDqEiuU/8Kh/WM+U+9T7SGh5Sqy4uSVY0DTYlCMyNqJ
g5m5TX29DTNuu9kMhrXad4a1fvg8bWDXQEY44kVXZqe01zkv5WLkRx9lIVTTYKozKEZlSO/ifzzy
5/VkyV9bzC5BMYr86ZLUNJsQ81NK+Q7OumqewXV946ecttAdY52aonKcmI+aVX34Wgl8ptnpepyL
5na57WXGnsfQsJX/DSjd8BScPungMhUmuCIw50fxdMzVenCP/uzqP5bM8oLlgW3Sr45m29z5+Yf9
0gGqfYcfIS1KiAdU83WWM3LSJjSjBeH5nKIGwJmUK6ManntubuFSv2TFxNkSge6nS6gLn6X26+PR
7/u5fFdAiNpr+cQ58L8lZt/L9+wffTRsJda183PzsjCytBdTyOB8lPmB/Ipyzkt00/7i38nNcrpQ
FR4h0zRtoopnwgaAQIU8HfqB9Hele4JM/NqgOB4gXB6AaYVyWdKtIDm662p7aUs3aHSQhQKdmkZx
cJilk/QyQ2IjvFsKR5w+9WPeFsQnK73Ojw41nxCk55/E0YhwuuRgJIPXLQYn+SSMARHb8TJyayKb
DfS34WQ3sfm0+0p8EQZ7XOg0T2B+kSMsVWn2w24rCfIW22841+OaDfgUH12/oaNzt3QLLmZ1RW4J
cm0swQdWawaHSp2pyJnWMecy99JsiPAM1aiGtBemCQEYYm898XBneNgV44ZOV1obvmI9wYz06xFS
9L7cTeIrBmQiqhbjZBSD2cLW/Y11rm7s1B1X/5moMBHV1vx3iWwsLbUuXbu9sPZolwCCRm91N5k2
OsM9pMqDIj7vSTOmqOe0VZJlvRXkNpJa4/uOxYdsrdBraVuFL7Oc2SIRXm3+N5Y5SXHHYaHFdF2l
whrL8nDM0wfQjGs0+X4/DKYmqnoIdSUouj7/+WbKKO2RsglgIW2Td4Oy6ShLnpCaU2mzGl69VdFJ
utdleokeYh0C4Mwbx/xT2BWQ/ZfH/escvDiwypF57Vd396J9GinRO5QLzJyDczp/KI5Zjm2iDMI/
94W/trJOImVv25bmBxY5gOXszdg0bkbzeaWqg8IX290Y8M1wrnwCvrxUXw8bwI+qIP3KvnpIPBSr
CMYoWdK9gQC85CJsUWFfQBIwKYHFkfEIuzUSpmoltneiDz1pPdpMvp7125lWRzr92Z4hVEyUN3hE
GfoHQmNJHAgkoUYEkwfCi5VSgpldQjD6YPBNll6xumxSAB1SwdagKauOYrhZY4QW2AqtbWf2WuUd
7MOK57vdeLTbHJWHGkN8fKR7FyTTX8771+bDvS+a8Xh4YfysRofzVpJJR60iu31+WfwHPvqxy6rq
DilJ+BMhv8MW2OWCKWexvEHx1lJ4+phEJ0J6olreuDmZ45VvOD4QW18kKXsPbg+ZPQ3/8LF26U/8
OsD46qMJ1Fq+b8jfe4xfHQvG1eXpQccjOxFzB68yqMWaiQvsYIKxWRPbHzHt5F8uyBPYWMtV3VfO
AivPatxmkjQ/Zi8lQRH48ZFBMUs0RbrOaFqUM6yALXtDVshGn7PRZrkmb4MJy3g0jyqoxQj1aGJ1
paG+jT4f+BqhUfpNUyftmm0EJr82mpzyzgWkw9BrH8aa2bfexJzzjbw2WMAtRnV+mWoVo0t9ndIW
JX7Y5rpapmMS/Eg237pa/lmALb9Vo+7C0KrsCUb0XuFVd+j8ZBwXPR3Z/VP+V37uA9aJHv6rGLTS
2hjKkKsnhDNiJ/KdgqVZDggvd/mW8TDgLLITO7iTm2bnZm2uAGjzW+pZJwzIqhyVViqdM2YkrGjY
XnVsuvDRi4Ism1X6e+MM6RsclV87a+vn8hc0D/ArNfxg+nFOqIfUkEjLeDdRIOxxzaUcDhC9Jr8q
OXL6WMgKV1DRw4ueiZe9NzoPQLAKV/5yG7bxVB8JodCyHtCS6VBLTdTpX2PpbwpBRR0oqqGIVSgG
yF9+U7/tCzXqdA/QZDwHoQztcoDLeLa/HYI8gf499ZJzeD8s8fu7JfddqHQvbtK00wOLvjhZQDCL
3QAQL0lUtHFPu8wh9gFYAbv7+Jj9WPRaF8vkxgvdX9upHfGxtsmW8CwOFjdGA5Ppr54JOkDMl1tw
Eif5F3WDrup2KzFJ3G3jJFXrfuoLTEEQnfZxTvW5P6pYIhYc3IngOLRWLqM7rxISjhJgEqy3sqeB
HPvS5phpGVygm4jwAH0ctzuydPnYZ4AJKHaeznftpznDNo4rtfqmqUaIo8HUnnDuRb1vnz3v18/V
K3NRcCrm9NRG6eTGv1B14M8NrUxrhVxTYVwjO5e88JGRrSJtosm8ufbY6+xUb0q7lmFTCCd3Fehk
AoaKottYuINBNK74x9VMAPdvsHYE8BRd62dDeLVANPCha9JOnIJCxcOmFzGS2iMKpYA1NbVuvwsN
FhXFbxs26QCEWXU3AffJTUALO1puhJSo+zuI52yIcHC85FDTo3xGbvSTOM9w4/yrxmohRiUdD9jd
l9sSII8HNp71KfobKWANY5ggqYxUl32QPSujJobmLxkGWkpbak0VUmdzbZF57kaB5WT9fQTiLrLf
D6T5ypWnmPynv+GlmsAqT8XvOqY+vEHAJVC55+rh26ev3RW7gwd9oShKmvqUfLiHZVylAX8NM3dY
XS+YJ7dWa9Rhho3xxh7M9EzgP5nkE42cTtAPtvMxUzxvY36GI6sWT6BjOF5YyywUAxJqG/GuBOLK
34OCSM9RgExenN/yk2qFfcS6gho41DJZwG/vOvHeWR6ktYv/YD/KXenJ31818Xrxc1V4oIOuyMm/
Mbach81YCgoxGpvP/X4KPETKyzN0Uu0fAiDLcuMhe+RTzonZ9w8/ulbuL3e2pb6sQF2x9SV1szuI
eeQwrpBT4LuY+ubFUNaBOy8nrBxJPSMgeAR7gVvn7jM8pA8BH35lDhSYftheEIL4k5iVOUL8JrZr
KEzaWYqTM4Dt+czSPnXq8BYHBeBwG9ZKZEHvUCo/fodrtNyAUZlsdNDeRV3vljCPvb6SBAkP3XEx
P9qHnrS5zFw+nzwoK+9T2d8aNkcG6zYiMxwJENW62U+HaQML58FisC99fEZWt4rvlt8+THTYQwhY
aYEzMnAOBYaWr8jzPHYmqlKN0NYNTYiGffS9tpZ0RQf6aFjSWaQp/RFv/f66oyHEctFeYf0w5c5G
xMZAVscmNPd6bWgwm2z3RELcVro5MtIRr9RSVGtIH+JLZEjW7Ascbbo0d12vRRkqhTeinZjGg+mK
Huwbh/vPXrMpN0VrGpH/Cb7HkJFHdOWcPHNbANQ90KcsXrFdoSzGtPfji9bS+NDMFm9uwrNQhfTs
bErRFQnXtPhuIf0R+4CUJu/AI9zClYCmRZGDaC3uGMjsQpw3YNO/DnS4c8AOPBvRvgEd4xyt/gTO
JyA7S3eBU2V9x5tAOZd3T/zDdZfVM6pqZQpmSQJ0XTZZ/PPPHcKdsEyEqdf9qB0fCEyRy0Y06sNa
plp8xKYvj1JGt+HZ4wfvLqlEmgaMYv80nr/RjuzfwMbo/WgBM0X3412akEVuJViDMLAK8z263Uk2
lrFFraR72fR80HhDxj7ntXHZbl/3MXYpdvqK2cEXMA+lUJM/v4ENEBrgMjp116k33JBj8+1pD640
wulXFZ1rbiBTJ/chNgEyLBaIIc1NjVujjroKpwzKT1VJEg8GmZazs5tsu5Mqka5bV6TS5dXT2+Tc
VKcawdO9dtOQU2R32zNBxRR+9EECbpa1Qke7STvdNQZJ0DSkve91PgwpTfG6NVPcRO3t4E95Ibiz
zs/bSLJWiVAQH96yTxZphg5XtzeREc1FHsbGFcRSJ+uzDz3BZWd8ZfTDPQpbrztX002saJhloBP8
GaoKgGCRb/w2aV2ao6/oIHwCmriJsKtUS3bTDBVFpfn5b7MZex1rEGaMidYfh1p0HQ/GN/TZ6pfl
lL7fg8Qr6aEFPjRiK1zA74MgXoQkKxyfb7g4Y+tZsZb4xxtyWQi7PnyvA1WNPxJsyk2cSBZwjlIY
EpAALed/AUkTwyNR1m8UT8MUrbjKZP0HDHJUV2KugM+cSmYwv9Fj4/Ns3GNYgUT+jLMwqRGwi2HX
xXo7ZTvYbWIyULhwaDryBGYqtRZtRD8p29aSqnwswyHWizKE9oelD0FMHVfUj7thel6MbygeJnHW
vP0/SsHBMkPLhb/SIx73erLKRV4CcLW9ZCNnZxWe1rTz3/Zx5WimgXMAB3sL4HDBoM7sBaTurNk5
rquH3qmGUtjuGbeZcAsv7P7XAtGGm+9PUKCf2+h1M2Ldg4eOO5rT9kbXbHaLorJ4PHu8nrJxGgr1
3WFJUUDK4VQzsdePigHtyfseUjJXqGVH8wtZg6hbHvSueozf3QN5BDeGUITf+puTQQpumMWqISMy
OMA7YEIAahImrS4zjPKZ2UWA/nX7sfRSxUegyz1sjL0FZGFBjqDNC7/hWtPGNZVAGVhJU32yvzRR
TSA4mXDe5JAJwr4KMDfbhvokPFH+JqUCk8O+buMrqwqlZa6nzUYjuVWkQNJlFyYyYuI/ekNDMIum
ZF2Skc3JHH2rHS+wtau3KXE8LkxXN2uJS+lolGADGTlswXjKifE5THGJVqFUvexZ2WENxv02lsOw
XXcreb5QRsN3P2foVC1hynVhzFn6pSAT3bBKEQuzTJ1fdIFMLPnwB0b6INrOdhFzlJ5AzJVI+PoU
CT8Ow5pOAfWf/uvpMg5cz32qko+h+IABGlqnRwGFSToXmrg6agfR+FUckl8A36KXwqx0XLaK5lkU
sSgpLSw/3sjMSnmg3MlhFWnPKqeFVNokC6r1oZn6a/PH1nxTMhd0PcbGvuxrs0LnznWuwdr+b2mW
UQn0/pYWPdZ1DrWpV2WWtqxT+yOObRIs+m2UdyLmpHNwFV1G93OAwf57PNH922f3+l2gqHGtotzc
4un9Hg6qiIliFsQt6gPuDK++knIRb6KRjsyXdT8mxP3mMrcLBJZlBd/jDHpPGJGNB6TDzmAzKfTu
WPIwkfjWuepJ3CoxfWPqx8OHDjgug12YEWSXLEllzvKannZNWtHHSUzR3LDQ7ejyZPTioxdbEhs6
0x+6huWdYmmSua1llKtkKWwJyjORn3vKwJXCaw/6C8r3rNg5teeCcs2Xqvk1aNd/XVlkRK3MgdBi
WFB78GY1nEsXsBmg0Ng0NEGb+kNVmwxbbMWDGRac8wh94NXuyzEJQE4iMFbyFxTzoUtI9CxI74UF
bIVs+OHzX27yxViAeMZJEUi6sLX/HIFOVFyyU0I2ZYtGNSGYDcvc9PXmLQ/cHn0FqecNfG/e/Feo
lIRU018sSxCEPzyQj37U5VwSzCdT/VkfRLIW42pwRb7Nmn51IpLK+QcWMnWbwVX29rq6+gJN+u3J
c+L+zmwj10WnsgGzY1j7kiZCoSWgWD3LIUl2sH3UmYcpCQi+TKLMMUDt+vQOucsiLCvT1U7CzBPo
yljY33dWNaLKUuFWkbUPLAquFKVkVGGGCsBmSswhS6ZTTwOEpTacj4xfGGT23qoTpr8j35Rjx0L4
lQxoPSZeV2th2XkrauYKBUkCKyoiDl9aEZgidZPmP+TVNn2I7vlbChgkJ4EA33iyLNtFky1bKt5B
bic63xFw90eXUPj5CnFwdsrgVKQVmSCL6OsiK8xy9+Pp0ti+eboJ2fHhk0mGYSU+FoMlyhybPeWV
niDVTbZCpmLaLBGzQSHpoNJrND74/cFrv3Bk0/GO5ljyw9kJC+rueG3Vy9ToG4i/LuX2RI9yHAX4
PMnEwi2u0tfPDzPUj/iRoV+M/LoccYmtAJ9gxG1fsWe98lsp21ufgHoRIWfVyw9k1KWXHIeub85x
gKcJ1986BYBKdt4sQjI1LZOz8MUUW0zBCf6PK/94BCfVzF1CR06b75itYUXL1rXuyk8T2uZeTxfn
Hqby4Y93o28Hh7vAwfhhDDMoPfAChDkng//+O4EkWemClZd4/snm27lCeV5u9tVRHrXM+OkVK37t
0JH2ASU53VBBu1x3vcVmUZS1HEopD14DaqKLrt3U+5AUsRUbwFHWeT//IYg1J2kyaT24cinN4E6+
t2PgRYDUQpXqCYXzG2kOcLwXJCimnQCGUY5KvF6RauAW3KuDrR9svL92tan8Ttd7s8ejxJQIAzGS
LiqWqPxxjPSFZN0wUv/QW6MzkM5kIYmFZeuNRTvSsrs8c3KqJoM680XNPkOWT8HOKO2M678RceQw
/PglA3VXY7ejLIVMAx/jGNlhDNmSgNGAW6ipmxKeK16mOU1i3QYJOS5vA0LCa0czFP5jIchLXtUv
lljbpBYB9OjMQ5zUvcci/VSV2MPxzrV8PqpB8TjMxrM8q9ZJdwp1Uz9KbR1G+6XSVXqJZBY43X/Y
hZhW7kNDfGldtN6BM0XbVe5EQmOdYHcU2nnIU+vCS8I5IwGqXfcQWAKjI9r6rzIB9NXniNuFsLgo
9O5C5jSEpw5PHpiMnKhfrj+GiA3VaFJqnCee+So/Q7il0f75glgC85PojdFFzahRFmCjnINA/l3X
TOCa+uqHVF/N0Eu6S/jbqprnnXLrashRStUHGlKP2g8GXWEh2Gc3aq7Y+1nBbeL6Roowz5guCnOL
b36B1h7jhYkpHy9tRe1CLpH4+UDtgK7JqGI3uiZ61CcZVQidtdHk+9/N2noputz2vP7/Z5//6ZlP
K49HQrIt/JcIKU/yWYasOBHIitDyAQ6EcOcR4XHJObBvbeMgI1kqLYT+Z9ix0NTQv+XDXc1D1i8g
2IroecEa6AVJJ48i8Kk21huYxS6eXHHqhTU3d5TPY6uhNTVp0vaBXmBB7nr8Ow1ja1gBKcAywKHr
e4ZkDeC/HIvhoLmLqMFUL50MXiGD848j5HOIIFT6XQD++cxbzt88pvg3SLw3K+NAMGDVe25L6EF6
WgEu6beoExyLnLXLr++DK8vAzIfWQdAOefP//7HuHIu4QU9zFQ383NRVHQ3JHMv3pVWAe9Jh8UOv
ZT8VCRLd69bWq4dkEhaONAyHHAhC177jNAxIUJnNR05wOGSKjsEBm8iZai47TCPhCKLI97utzjea
i8ASeRFiWvQAPbcUDXBpZ5hzP7OSXYBpd8fFnWBHDIocuf8rrOsXg0G8EHEnLid/QVO2kaDuBP/k
KkgTVsy+VMS9FxkY9wisyNPYF3oaRRsGAcPtIjixNHXSr+AIKDC+uQP/VrvHqHvm5ypFomQIqNlz
OSDb6b1DbEgjx7PrWUli9ubYRA5FaXCfpF9Zh8d8Einll+2sf0xKMMSPfScAIgDlKPmiacUq10Bk
EXQUQ0TAN2B8UADwY9wvMTlLYV4aCGrugVbKTsjp2kvGMArIHP88NFJrtkEgg4pLmizW/ob7+Twp
QatI8RoLQ7Y2Gqf/samqVM3Ga1C8ZVF2nycbs33xYpJJplgLLcuBQgTooUmn1xrnjKJtQ4nvsTkZ
NJpWe7K7o4AydQ+yPwE6beccg+I/RXEYThsMpQvT313la5h6Tct2xeieq/4IJMhx9UotospqBSik
eWsHifry/UVOegjhmQA/uhJMu3wex+O9LQIKzrE9hEh+PnmqMn0AEvIr8jLwbegxyi/x07hNRouM
68fhaH1vLGhPglSWuiTWaDmAgV2Y/w3hAHRVrf6+lLFRevBV4L3bsJSbiWE6q53iIhtIQTBfyK+I
aiFTUnNMHFgB3eexV45U1jVF4IYh2OjGbHRQl0fscznOfeuGQG80vqgAoeC4EwXIBW0tseIXzuJe
++NrqxnP54YpQFypjoSd6Eq5APLOM6a3LPwaMYUvnIqi6vgoxtGrfSdqx9RONA6hgqUBgUGBIu+T
7Md4Hc/2gOIRgbQMjMcXOKlQklHD39ZpAx/mW2n9QUJPF7fqlY9Kqnp55e2zpw3eCKXh7P/H7umj
GDG5l9BdmCLJknRlFBz01emGPw3yv9joDBcKto6HGwepg3KvATrq5vIeXZ0urbUQQ7dLGTmdotCv
PQclkjSjy4fX0wSkgACfscZaM0m9aEyw606YEjtLXPQt1Lkk/q4l8G/E5e5VqE2UfzG2VYDHnjOD
MY1dtGXRHbLOK2vsO5B+43n8viswgUgG9Dqj9yPvRIhjNBL380pKgBGxM3S1w+9kn5Uqypc19rrq
sTy/hEHJ9GhKbygxyXSUsxq5f4snVYg7/ZgeWY8JWUY3gyBYSQHonWlvXHC5LXNolRJ57DRYyWka
d5TX9KQvIszvCzu/2uYZpzkFqmuB/mm2I/qG4LljtWuwYYlAtF61Gt+8t8KD5da8wR4k9jsshjbd
DoTm/J/68m3dcS4DMCswUEYZE2nEwu56eBT9Jbgayp6TC8e5TQqH3HbjJLl981Cq6NKnOYbLLvvH
ZDDAM+MHG1SfF7u3dTSl77Diigo93GMD8Dfy6BqiTWdyjBnpXxLYbNlDY50yuRMqgHffCtm3YXIX
9EQY/2Uo/MJMdqPrVccwJ+7mLPDfrfV0rhZBU0vA67G3MBo7JzgEBwhL+WOwGeAtLBAHFaZXfu8u
ZSxc0DCooKCfinsPzJ9J66SrXmlMoENoyzciwSJWqId3w2yxsAhAARduLHRpVQvWOgqcIMfhEKxL
xJeuQk8yLVNzE35XZ13NMZVe3Okzd6iPe2U68BkQ+IEBpSWrJ3qmEA9sdfZAlyCkxxAoWqRQ/sP0
GmhAs2jl7TZHoZ1z2rXAfPhsbypRAFb0Mnsa37lbX0QKO8ZIucyOP3VCaCtRoJJEEDug40zeVRbj
g6WBu1kAnaTa9sGtMSuZPtFQGgGE17ffWWZFqDj3Ufpv3ACN3yK6G1tBstOZCKwXnvtTM1QOl1Xo
Hw+Ly3ttjd6Wn5gRhFKB6OO/7ATOQqepepgRreplRI+RTrwdQ8UA+xIFiXTEzbRjYt4hlA2jPZ++
zjBSdvm+Z0iSV99zmdU9BTSdsiwQj4b/kN2RM8yZ4qFEKP3pIjPmxXulSrmu+/Z8fe+rRRcWTSay
9Z+L79FLdXkKjIRnMmm6qYdzfoObuPU+oSyqz2xfmomOYVk0bZL3ywNCtdg8WeziFcciI9m+juJ0
o4mkfQbTzIXjokURPeP6cEzA35uL09KJp/IAqchcMAVoQyTWFiaogtp9UQkgemHQ8diZG4L50a20
kndP8l94rxxgGPnD0dw1Yk8DL1VWlm69HHpz+EtX1wShQUB/kgnMzCelnPbTjDrRyrfScWzwzepl
JnOmKrIUhLPHoZj/d+xGpAtVPNtz4uBUXUQMQSjISvNzD+07uG57LaZJTveL7ENCU0LIjseL0ESp
E+bj0JoazB1Aw4HjL5cUZHCVQ/2huk0H7UWN28Mrerv/NuOYr+4tHBuZ/8TZK5uqSt0y9muUUk8a
bTImJxyVC6lEyPK4RgM3767qtKAT/87FJpDDYCZW6F7gN6CrqvYlCMrI1eYgMwWSS8hGv/jwnjV7
4yGxfMteIaQL65YR69dmm7Qyf8svgeY6yLBGEJiZbeFMz1j1xunLTh2BWet0pIUEU+JyO2d4C02h
lpXPbsmdBvPY9bynFo5nDjDGvTk/la2hE+U8Qh+mr1o9o3RnVKls6s9bhl6j+7Sc5bq7wiMkiluq
hyzIl/Vg6X0cr5uEqFO9/RPKrTZ+T1AwvyfRZDL20IeyK5y+wvfJiHhagB2/zhWMptxT8KjT1jy8
M7WBkdEADwHP5qMXPJopkQ5sbGpy+IIWn+BewhIQUCJcV3pSC7mQ3WASR+VRfR8JbLcmzp4y989O
BP0cxL5xgug8dGxvfVODVShtntOk02fG83I4c+cS5p1HNL/Alq2cE4NEtYKtbK/Z+Crf9jpow/MK
WKP99wKC9tgfjA8Ov8c9UPbEWczrKn9H+zHgkBE/qT8mEsDUVYb0KX+Uvh9jKpSPz/xBAehBKS/j
qBGIV+sl9ehkHgqQwZIGlUdBYudahOPa/xitaqjbbZP4fm3grPlCt/RDn6czAPj8MZP1fZbY58WF
pXdRIenQjrNWxJ4ggWHF3+IKzPjRNjlFXg9YH6yUFeBpAoF8sQloLkNFp5NA1tfDyTQIIGM/P2vu
RSllUckyYuJuM1Czvrypg7gS5LIuKxveKu8o8ceHeMIHSOUxfN+0umz18+a79y2cauSl+lMorEMt
z3GsPUOhdkYp2ENYOqEo883+qD/Qw9OCDo4k+RePMhVhEAn/YnAhOKuOZ+g36fGiaUkQweb5XefA
WWlT0eS3NWZFFjhl9ojaVxL0kIviCbxpk3DgHixI0RWCIQeYl5I5XoLpthKZGYHyYbeD6HT4kz9Q
RhJdL2JtR+txAl5SYP8CxgqVt3yK9Jm9kOqb2K6NVQxkZlV4VHfvVvT9eLWg5Akns7u0AoS6FUDu
7CWDegS89KaK9B+QjN4ugSiMm/ofPq3bLV9ntbFB5V+hOW6Ovr5zM9Oz0aYKz2oqctMcVkL03DD9
tHSARr2SB9uTD9glQmPt/FvzC+SD6vKRGsAUzD93nRfFoGRLEMKhA5Pon0y3s95iAx7vdZe0kNGc
XO62izX8WJTqMXpnJrgsvYZSlp5Y42+DtigkjZYBzeojKJkvy+okvL/AgWPusSroX33Y2ARWFJRa
Tgau7o7WP5fTQcfALgw6uBSN4LqGT7mnuG7uo7swIr2Kg119eDX0wE4pEVCGQQwJdyn1MfO96jNj
8aT89RpA3hFf/zWur8UsMimFU+loJo3o5MGxluat68aRq7mjZNGF677bfInTmmQwAGC95WMEM3IF
PG4h8/gT1KoMUqKS0jZ8sZWlR+alYKJdoxgSRYwuBxMVA6oVuUZs9QWMGXe80fyPq9oachvi7OjQ
gHEgY0QgrkBTZlzYdWYvh4YyOI1SdsRRZBcEMUgjs13F3IuFQKbXgznDHnPrbVGnHABlOJPQN41x
sL00t3WdxtFPXMkADQshMCl8qPwrc9MqwtRotQj4vr4v8mjBu9LgJusim2j/tVmAKB/hpBUW2O3b
flQi4oaPlFRzl82xvIvII55aePJjuGe6MwLObgZAmXldBQEO3Yv7UkxctacetWka9UZ+5rmsxB3L
3PZm4DF6L84kgsWgYbf67I1vvwK8HKXoyDTGV2miAQ4+BA2G+VV1Fkb2QvPqgh7isJpkI7qNI0Uz
VJ22Y+dxs9vhOV14wgqJxxTZwdZHXHpS4+47+HHwRLQ0KMMq03GXJvQgl1pMFI296OT9LDG2UYbs
MVV0ZBjFXhnrJLq4tVHTLMT+2u+3Tur/LGFL2FsLpJXw7wf+2iNZDQmElIHGMUFJejVjr7nZyGlm
npuJYxp8wAUfHrAbOdK62dtFqD9FrH6yfP7AjqH8G7A2pZ9XsmBw4n54ukQM09lM55D+xjPSccrE
DTmLCRKxbg8clzM/3lw07nXEJPtVKA9qai9Me7VvlhqOprlBl9WENdJC/pVY1Ymf6cmExOM82gc5
ZOuQ/JWyq2x+iUkVJOqhHtyFNxH7/u4yocr5y5nNSZeHU9GuwWjezv0aYhegKXAYxGWrXM3Ljjyx
/2TVAxcKZBemimrv2Z4wzOXsfir7QzwC69fJIe2Lzok3YRhY+Gza9D6cjq4OfEWreDbjHAO02G38
ua2qhG4Dj16h7TEB0OOmSwE10gNT1ht92jf8+VVn9u8lANUkIHorE84Vz1BQmr8t8k93NpX2lgpN
WsmhY+KgGV6N4PPDM9HNG+DM8510Ei/fpqOgngMLF1vuFSaiRR/Fajbi0z+6Xpcw45Tw6g5MMMeC
MsVO4D6W1wesz6EPZc+nU7DVJPEC69vCvtOL6LPZq0j+bTgKlWDzvaC8hudMMgS9aXod+DinZOd0
to2IzLIohneuuh8+KyvYsE14PjpB4eCQvl9YuR5OC15Z7oR31eptdnjYQW46kYtAm54BSUarSsWj
4j0juWuTZhyGjHx52LxW9Gr55GhBDR+WRYLXG0VpEsWM+CaXdVW9FPJBMAEAtbZLSG0sM747h/jJ
c0KZGNKGGHdxkaBPDdOi9Ss+flp2sL7c9sijz4RPNgcH8792EEK4722r21fR+UTuD+mavFd8PxYv
FUzXfc+rEX0xmrrBwW3KelFcCBMuej8TldfjDbA4TFuLz7yzOsOAAx/cngi7Pdl/Q5bX93rhjHrI
Ecwsq5Jw5UUcVaLXHiwwKMculh5mtbFYn5nGviR2v9xMDQuB4BxoURsnwVTkpHw7gLYgAmiWF46s
OLWOtc3vmF+L3cjzm5Y2DR49bo7FZC/NSrptwx3ubvZYzzSm7gvNf5Z/gcIaJ0ShZKOPJ1+lL1n1
iHb1w2N1LRQcR3yYLj5M1RyrVUpOveL8axCQp2zvaos09Zjbu6o1fGNc7eHtIH7BjEBIMY4bx7uH
JN7ZoOsTaVgb/cy36Ut3pa9i2B6xW7J+I6UQ0jOOYu7YUikxm25m1u45Zul5etoo4ChbAZNBoAOb
2aPEYarE/qI5aguq4DTwGgS03E1Nt0ibninZPIUklrwaiutXXP1RZMoj2f+RixqZEjrllwyUk+C8
xOe+8Hlfel4tYX1/krQ2pBB9NeM1Rq06aHRx/GRW/optdyBV3JcqPI+xmOvbY4z60chxvZFlDlGC
rugdX3F7xJ5lggeiT1SN8D0Hg4JzYX5CsJU5+jLB0zd4mmA4v/1uABKJFMmxRXEktNvd16mK7OtG
jK0OfNC0JJmmurImuTkuB7Epu6znj8PXwYiUOX4nvzCrkdGLob2JV3pGLdYWQR+ZO7ehM3i0Tgvx
V02U47OYO0QThQHeyi7bXA9NZTIadAV7Q3H/JoYZG7GLI08gjk1s6e8NTQsuY61IwVy7kX7ljOge
HMbIfr8S1vFwDfpihI4VvLY3YyUOqy5PmcJugrismuovfrKVzvNPajY3V+MNiUAjw44/2GYeGruC
uzlp70GjuyVFf9P1gYDE7+ZmkgO2wXg8/icOXzVTsUGMtWUPfeede6scp130u44wJIKrC/AURSC4
TaJ7siFeGFJ4R6l9O7dBmSwuFqkBhnB4X9u9SZYOEsq1inPtKgBA0KGsLBv05Qtxb+DJswFnCGGF
g4BIID06qSAFSImD09371w1m09fpZ8LbbVSm3TrfpL6Fu28JWLvXAhuJ9/yiYjJRMZsuMl3lWOS5
VlCjRFg2cPphDCpHcNww3noCzAuifLxL996rOHMn8Uhl0a4Hm9z3ofoDFXLdCDlrBn5NfuO1x0yU
dPx3IybTXGIrFjilFKE9eRyzuEVC+/a7+nl47WbIA50MtXRwGzZo5Qf27nr9KqEZicRGtCyUSeAK
LuTLmulQu/e1LjzQhFF9SHaqMvoDYRsXsth0uUj/l4iL+hxd8fgNVhe4KDr5xs8jOxtkhLiNHTYS
Y3225WzwIh+9akIzTYe4QZgDdi7Zg3SgxJ8p0Yem8gqwqEAUKmynRqf1OxcauDdP6CkBAUdhYjQs
c30cQGsE/qZyvCFWVuc5r0cwUWXPLOmJz9zSVsjfgqqMlqb3lsGTxLVqr5KYifm3OOlrgotFI9fh
jP3bGFNTL580Ej4LImcxfzEsM3K7P3zcXLJQkceVOUj7Npr6jo34R8m9wJ+/wotTNMk7hNdlbJuy
G2nLATIr9l9qRQEv3ccVs90LWjuLmV7OwoKxOYXX4wcX9az9gvoabBqvOSfHrqxra2s7gH4G+Pj7
U4tu3MDuA2sjMYlLD5UNzd2ipsdiaT/SawcpH6vzj7YRTOGYr4Y4tOnYZP+xfqwA6q8yWnl6h332
vYif/u/ZdtwWM7Patz/Pz81jkpzoEDiIK1qF8b6j/ACMefRDKTGWvbbeyYGB1tsF+sUpcgzrm2QA
gykStBziBtxnGUUXR6FF9eypxBcUORCeTrs4Ricv8y6uDx1SZg4XaAQ383i1zAnyw8dM5Pic9Tgf
9wbQc6oWAao4wTdZOTESb5h/rsIfgluohvklIGv0eZuhFbj21Xb5oAMMUwcXIrOiGrnr99pcTzGD
4LUn7UY5TIT4hnz9ujP7bKePNRHBqwwhdWQyv2f8ef8Wuu3rPt03n0jlR3yApiISwEiGPSJlWiZX
eXrR3CcUOJ2ZEVu0xswMjQPeSJ7oLWq5GJx6Dv/yBMMMdcgAjvCQIV6k/39H7rk5NKpkPWX6UlWe
LCpoDqlGJXAilnzJDzmnpKYdrHt3x2XwRZMAmaxffDubMXNvLGgtDqKtoEQ354sdRYxQaZGBGkYy
Eh9oR/x77NpOLaXeV/vVW0pICy0/AJXi/L0UCo3VB6OYwWgmqDaZ2M2gnT4Jh4/aKAu4H0wRUlr6
VcoViwnA9iqg2OVGsutictShLUpNcu/bWiH8tz9YMiYz8NsuiPChDVCo6qwuYDjZWh5xhxef8U44
IJANJbG0RLAPbQ6Wn2jtnL0Bohi/LjXrJw9H8ck1uPUeA67gzAiavmMcUmD3d4/Y+FZG3kmpkgb9
thlLni9q4Qe7a5KwKtDX52DxCKcIHXliIjbF3GhYiKeJbnxTLtY1zsTuAUhaWKgDmjuHDm6gTsXW
ka9pm/fPWroTm4CofqI3elSxstQTQc3VJ+qdQctAlhXOy9lj6Oxu1Uj9GA45lKjq157DRsOMCboe
EyfMDhBdPuomlCWasMZ4f0kkLnikRoQDaXb71fmQtPy6Kj8s+IyNhZcLod7c8XDrffgmE31FQAgU
jW2+epvVSKOf/e1jB8YVw76xi8FwStC4WhvrVwYm/4c1IOWzDzzNX2E6N3nzEp6jcPl949pXd320
G2+wFoyV87gBMwKqeKWNw8302U9691bk3FzZZiZivn4edMLT3Tjaz4zMkyJWigkO0avL/yNd6LTq
K44/fg8PBX0c8Xd74V9HUer22T8iLUSRqutwR8EAIiFDdD2kHCZDLLb6tEuXTyCEZXahWeU7zHHl
jbtHypsEkAHKWTjzC97ff45g8YHEq0ovFY3H0y9PuKtb4C88vozQ1BcF709NpjyMsGhU2RTZptKJ
Z4Zr298ndex0sIeqaT/P8HPhFYIYfKSNcPWRneTPdQwJr51sWiMFKk54s3h/1FP8jhz2DnNBLfA2
RqWzYhRqjKr+RSI5KRpkiG2sX1HuqLoUcDEbEgvyvYe/KltnUtUD8kbYjqq/AXXjz7loERIjCAQz
Y/8xfcFfz1R7awlz+Mwp27v/v5nGa3MxuTjyc5IR4QnucbIHQR+cunS2OpCGaSlR0E2u6VIzi2NL
b+b4ac6zZeKmEgjC/kbZTY7164hYNskLzu8ynaX5+y3yx+EhuQ138wvzuqS6Lys8BZv9wPeanaBq
CuFQBjeyVbBg+BBxeiMNmiz8QV7+9lgN2yrU4RCMOHJfJOUuE4ZzKAaSwAHTXT9gatI9H9ernlSK
S2xz18S50VhqQNEU4WxBpqirMFY+p/1kYZk4REoS1OY2TfsyUHmdrICQiWV/2Bm0+q063KPCi9zH
nPxdjlpeM17qFMtPL3rYOMuR2cWw1Md1imHqq3XHpfq1ltDFtupDAjKWE6rUoP7P6pXAORXH24PH
uSFHQisNt9vkeWa2+AFEIDFjb1XkyCmJNdAsRM42qGDOrCR/IltMAG4as1VUL7ZA+z+4W75HPot5
hhyTBZHsfOB/Xta6rTxNN49ijHaU+kbYZZOE3Mg8Mh2qixzAoiXheOOHgnMYHOA07iFIcTzbRRwG
Ftw6GPYASXv8eVyVDRffrRjCRWd96aEDK/3LaWuZYbX2ded9Akjz6MBjjdBj5zpyQL3Wc9s48yzF
8Gej1rqYaLw6X9lTbq6d6fl1QvPeAxVWJBir/rE+uqvLTbVD2WQOah3bAOqnIlV8fqpSx9ikkcZB
C87jwU/kX41+bFJM1m7IJwpy8yj1DFjoTCesjacd78oAaz2XXMCxcxcBVhrGjSMxhArX9K9IPBWL
dQklRyfIkAM2IXsojke1iABUEPfcwUN+k1eOE0PFCnHyrve3Nw8l3RrZdfGL6M5xXd1MNM/1Z8cv
/vFpY3KRygRplVvZPvVH3+8vBfaW0QO2F1FUgRFiHtNaZEtYN7iZdNCP9+h19McUorhxpe/rQmwL
1A8KqCyiFuEIudXgGNtLSjH82m6EY4y/GCCM4Lej34861lO0hNZFukvSoO7E1zHsl/LtilOPke4t
GzUsjM14kqlsEeV4rmy8Z8zqAXLYpoS6CK1/85pJx9bFSLtqF39NtLlWAHrjQa45eZlhrEexjnzR
bsl/VQ2+DKd1ReH++VCuXYR3W/bOG9XBKXbvdwOw4m9D0DTKwUbH/9LVWucwbtRHWpR143woe4FL
hjhh4wckAs/JmXnB6+bsbKr+uBuV/a8+zpM5M9ealqwdEWVoON4srtyetHikWq0tHLUPPEHY2pfa
B+VU5/H8d4zM2/DoRI1RLGWM4M8Vfm9t858T6fQv0vwLZSC8eMrW3rTa27s8A01WPDnpHGRqSfh2
UbQ94BfWkDwQUacNsSghQk/0ki1xuaiU0vTNcnC55eoa5sZ7l99+L/K9CccLVbW0oRrQSUaRdlg9
93Q3E+4EyyFY0Ejc9h/+Mh1iKttNqiZhVis+9ypNQmzTYa9oob0VlaiyWk0bsdU8HfLZl+ccv7Xo
z5BRu4u3rAODWbBrbJh7eNmqbt72TH7/DAy+UAonU8Zl5BZKuKASLSk0giUOU+Tdxq8XLk+u39ta
MmVvHyR/dNwgSTO8xLuxfgp5iykZ/jv8p6ix2JJX2jLNy/kFtEcccMhVoAoCALO+PSYajB5bGfQr
y2adNja5tOpWoZc0rHD/fJXMoxPiPA2s2L5EJcQGJbD+NXRAet2jQ7MpVZN7zV0DVat5tceGRDra
LFOzoXJz8dquPfzyI6SbTh+RMTPUxFHWAsPML+/KvXG4tTWVYMsheLsqiF+pptTEGslwao73nzgG
43YezqUQ2O5BBwnT0Bnb2uqsP5aZI32n52ftHa7xq+5Qz44PIFv7AhHa2f4akv6+WVsPLDWFiS+P
9d45dNEP08Or9KaUzis7P1sTjunDDNPHKHm/3A4n+bB8zfJNCqu6CB8L68xXwhYCKWRVkcQwQzPJ
s0dQLYFGPLZJVHeJOxAS0bKkAAv0ivShpdtivRQfZVBeL7s968NU/LC4U5IkA91qikUvh6zTBPBK
PdngCfC9zbnxpxQuXw40zfSJMaJFLmBl+LRPpmCSvVDf6CcwiPahdUCyIQoVqpXv6v8BQd827QDM
Gnx1xwQyyI2FVEaO8DOB/x1kDjEuQTf2SWWvSt2FrpSbDyFusA3aR2b/aRZtM8wfgTp61WTgxt5z
VFin6uLVHo96vucws6s3DMo2gyS/H3oXEJdZa1yAghLnM0WEr5MmY2yO5p/NOKwMOaiv1eX1QgFU
GvZPJ78RZRIjjckCUFTCTIYK7AnVyR/MgG77842hOrA+UAKpqv0V8JIH2aBA8CewzL91RLcUzWYR
i+ixoALp+PBFqpkZQDFV8d7c3GOvS3jm3kAgoBtbdYXaS3orsQvgNrmYwOHupU0lpyro0qLf6Tx9
AQ7N1r6ltxhkMmbjwfPAgMTIH+ndhAdW0b8loEh6FK0+ibpGNz9oaAqsYNsDwEqHm0TGav5x6OL0
CHCrxS2+d4HO8B3K5d7SOQbBRSO5Yk/JLlndBYxSZ2Bz0NBgkl2BmLcK1Jk/CrLtkgp1SDTZ5EYw
pdDIbvlv7tbT1ocLD5Twtd4Na2S9eYJb1W4yCOytaRjLYVp+6O7Dgb/IYqmwHvssgcZ2rInoEaa6
I1MafsjSAsStyILhK8zTHwp1vVcKADgSR4phEcONjN03ZmobY+TP7vVdYW16nltF64qQXxY62+gW
xf8RflqLiZHpE+G6YNQ9KY4ZQ7jxG3JRM1FvN6Ov9hyy0pdeGyWDmfDQRxyhcjQ51EKN8GQPDzqi
6gGfktTeuv8hQr3oNiQ0E9ST5vVM5OGj4Su5r60NgeG3HulyE6blg1GRBis1xPREnElWoV6pd+w0
tndkslh/wleAMXD9Avwbgsg3jOwe5n3PWckPUOif34HzSh9qj9FN8BdtwxDv+4MG3pd84CL+SGcJ
lH4WsgYKBodTMz9v12xrZDJFBK02cl8lXDcO8QDpu1tsG+K73ax8/kq32iUfO8vYRpJy/GonUE4T
TdJ/za5HmSXoLZyqiYJ9sLBn4VAWhAi2aDtaTjkVHvPvJcnOQhdyyCMY+vEZmmSpLyJQA9CMKRwI
lXYHZp9eoMDGPdc5ore2W6aGSQmxQZrU7+hoe+7ivNmnlD8m7x7t7mZVC6ZmlCO3sgUw/uohpjvs
xTmygRGrXEgqWZekKpWpC0rSO7LK+5yj85mlYOw6EFoLNrEuPwrZeVHbofQM1o8o1Op+nZPu1n3V
GxnSMaFXkaA97Pc+eYff81Q/nvOfwt0nmfaV4403WYzmeYOVDv8ldASr6a9H7WAAhuwJ1zS5uSQ7
e2Zf+SOJ1yC2xSwiSbAfUvs7bhO+CVEkxoFJCj0Ai1Cf1yuHlGXrAKUXrl+1BqoeT5zAk9w/X7O7
j376hzxIcDPskaLilQMvUL3ocEnSjbXiPAJJ/Ka751eIMcBx1m6AXbQI75x0mTyrtlKbG8LiWbXO
xo1PIbNqlUN3bMOm4rSuoStgJ9WUcC9P7QXAmfWgFkZ4wRlM9b0TkGpGyejymgheZFZN9JZ5WF8H
2u/zeC/nLZqPgt3gtfMvwWKZudihX+ciscLjwYqL+gfPfW0OtEmbvBv+cFGcC8l9UvrWzd9POBq7
P5Xb48Yl5Fhy4v/BgdHO38HYERWOqX/wUTdwX9+F0Mb3DeR5lu+pvsIJTeuNerfZ4YXMqp0bV7jD
8qp416G7VC08DcFmrTCtoZot/om0Lz/Wc9DKxuPAVd2k46kVWKcSur+I4DWkZB741YVQGqcq/frw
43BR6WlFyr9OnC+5Pp/t2yP7B1ppk2K1Lr8xJpbczwT4RnjKTCGPWBBw3dYdaaRAkcBHn73vithr
dKdY3bhPsZQtFFxDDrCSIIXOlLFSJEJBoaFMJORts3SKz7vBoh0vaGfdThjLaECPq0bJD3ELBz0W
AjvPY4fP00DfUh4XNgZf3ivCoOXcicxfd4jI8D/mmyQBfs1cedCtj7Xzzu0a5ecgShvATuElOMK8
ZVzKTysNZGIGQy1pOGF0TROeynvD+w8DQ3IXIPmzHjH0lGwis1St50NHJMpxkFzYyx3d6Q9+I5c1
mgHIxUy1e478UYlaOF50IkT1Dx595f6NfK2fPUa7OXVw1MMVdDePhKAhCdcnXylLXqVSsT8fNGhY
xFPZugxewImswPoGqPaWkRM8bY0JsEE1QFZHFE5VuB6jOlVVEN4QYZe1dQAF44BVOyATJExinTT3
vEfo9e/fmxO+2NlUPWery29DWOv0fOX/dl+zQ9GJpHhWSWQLmGfG49HiIKblixBKK1q4CWBW14Ys
wJtPAPhrs8TKfK19fCJ9I/rrs7ToARg5/ozEAnBeYshdH5KSuFlpu0NgUn/VMzbeXzpFyp0NmlZu
e42n7WDpgjb2BcmmsrhVXa/8ZwvbdLlRXyx34E/o2Hv1OF7CT8I2dYHygXKD8lU/L+oPZHhrbniA
algZDsXIcGrCpqZLaoM9NWXUx2zwqXFwWoUgoHJHoSdeW/aBQZCYbJowoMr+GwM0Keqqd68QuKOX
E2FwO6gMD3kyEDfK23gFsNOFQt7Nry2ibMMmn8XcGUXWYv3bpYeSGXW7qRXtipoL3+L6celzd39Q
i3C/il/d+//Yh1xRuhO6/JT5VJr3a2I2WVjdTRSiK6VPfsPzbLTPrwSfY1IOS7Us1akZINALkkiW
olY/rGjQVCvwW3/MEzQEJeBryHviiMYwFApy9XeXgqi8fP+WWcMMVuy+8TifJOUjs4FwqER1MI39
pIelS94J1sCRal+Q9pYRpUuxxdTilBni5CsOVJMpgFQA0YBGAsPiaOR3F/L1D/4+HBSeZGd11YoK
xU1X4VdkJTBjoZpGaKa+6OB4EtV5gsHvt8nnA0xOyu3L4f5cYSUhaFqO5eUZjWC6lwz5KyfLsdep
4Vn44u58Df1136pszOWmYjXhpsxFVOxkDT+BwDfNo3xSCezW5NQ+pKjw2yYMs01J9qTHvt1hnWgL
oVOQOALL+vnaTVT7ikgXdM7KitDqGO4+hVBLk3UonuktN3jQ+FTyipxAMs98eZPi/r8V287K3Cgc
/E9dXiltadyXGFMKhrp4Q2tfVXLnbelaTTRmVwCQQ1+IkyptoODcAk0c2tB2FfJy3dZ0QIQqrN/V
ya6iLvwEquPrdDjGeNm836KQjtjBLTWmyXUDE33N0YNzeG40pU5GtTKFGhxwvfMbtoSfoZJpzVqz
c+f+V9VBvETxfFblnWnjuzmFSbb5tov6+PfM3XtkRN+HRlZFGlmtXgp5voPeQxOsDshzUYPfbf9u
dImcevaERMCTeoEpGxjuCXSYeU6srpSqOOTaZisfzP2FXHAUK+HKViJW2zmINpGfLV9pCTKqWQpw
MmnPizJLxLPJZERZpgZzdusoJMby6Kl5Ehb0Iqv41U/52ZsKZ0lREmo0nlicYGfBFjwmqKB1IRMT
t2YIylzPWKSeZdjzE6Ngj7EAtjiVWCvN+xLobsKNS5s1AK0rh2fIxqrAG/0VdwvFviViuOKMtERg
DRmTJNut/urrNHHMC/cnqvsie5fXc6FX5T1ujpCV+PoINFK5xkALuTxrEwPsmYR9G0XsCyn67/OB
0HmHd8wy4iCgNTeiT/8KGo8G/QXIGOV0ZqPyKd6JmLpSFLUYBeqoyygsHFS+EmhPPDa22BfF0Qlv
SoAgDEEdHlm2aV87HhfS6TFwDr9kZccKxdL3POEtXQgydlB8LBehWF/KSGq2YjGbwtkvcZr5pTGz
MLVHmhqME91DSufJvwSfzYdepSLVWS/jSpioad7Mvs3K2mFFz70IUj7EHKsy8mge9+YmAEQT3BYQ
z286hP6qnWOlKNs7hc2IvsMiQjULetGbsAfQrUmBZfaubp6jFzywZc2I2iXm2/WJq+7HvgaKzj6W
1yNuMZn03i1DTFuWOq0w62Fmt6KB6nI1kThM8vVoXBFx0893xtHhwaUICpHGjtHgglGu2Xf1KoBt
jaepmkG2m8AqltY/rm9561e+rFP4FtbBY4OI5bz5m5r4zxyAcNSjy7okTbjGyh88+JxxxX45HMhF
+/FX2Q2z1rgtvrRwwkAmavkbqkGsZnqCr8mQFCYHE1+D4IVA61Szos9esL65hO0uAQelgIWKWF0H
Nk31+Al5OJIijlcFrhoLmB2Tb6+gF3IyFNYa9U1Bo4DKuJXxzzIqMboFTI50H6rd1544ybXvgVQV
OmOMGcL1E19wnrsiX+JtBWbTZS/E6jV5qMGkLUJXjQt9/NtA4lj45RoHwJV89Bd2aXCiqSjZtvxc
BBBxZ3QuYENJtOgkcOFLCiK1ycXevWWrRjTXDMWaw1pBOYvqCEcGwMPUf+A3qrDWkOvK8rU+xHFE
1jOz7w1tZLb42M9Ob0+XFYxG5zDpF1jE3TyEOP2rYulgf45YouSiyrrdxKisXfFBVg6zkR9Wcrp3
/ntoZCXPwTYf26dMYE9PbfpphGTcAN5yieZIy5a5TSmD7XsShQ8jhUozAnqEvI2dCrN6IcBa61bN
Levr8boHudfUvEmmoA5UZQt75bnxHNuxetpP/Mi+sWQEVxG30gMbSLsbHfdIGAotoJkCxyE74zM4
84vAAbAiWX+zFGQe3P7yFqPQqced3b2TZU5JZxtzW9JsKvtZRnhlAGxteRUWU0YL1GQo0w+PUXTU
xJHn6E+iJpC/c4zkhvBRF4PfDQaffPxtJH0/LPICy5TDYeL59jaQvkTdOF+u3WmV1ZFfd2SY+dVk
NzBDpGiMbDGaBwGVYnitCLB+KPw4qY3fNUj+njwLlo9x1yISMU+DZW4TJ0DsZIpgVFqqNCl6Sjut
EziBmQLWQ4eYxvUF/F5zR+TE5vO+YxjECweJ2feNUAxx+bUQDHqu4DxvvvXn8TVja5/AwEEkFLTk
IP6psX7tnTtiqgwcGxrv4yRp7jXReGQCl7+HdvXj6SwhSGKLRqvcdDJwbIWx/FWAVoz4rqBQMjz+
rywYc9ZXY9NeDtfepkj9ETPjCfSj6+UKCwcmLnqnHhC5g05TrkCF5jSEkofXHvTRzdvQaK27nHpX
/l1yh3h+PrmLYCNs/+U/M+5cJiZIr5+qFJ9xcF+t+xev4OAjZ5ADT1GLdaLHEF4bf+ORgPrU9DmU
p5NWy3h7hMK/5jVXXvDi8X0R6EEeaioy++yd9pWV58iQG8LODO7YpLrA7vyYNQt7QQCkYp8t3zJf
RoBTKGj+/MZPL41bXUGXQ8lHH8bzzGHcN2inNjWWUCTRB5Q+w5KU18wo+WZim5JO7sRPD2WtraEo
uqfD5uAXTOtjXm5U/l9PY5RT9rzUO/FGFo5hd5lOpWgFeKNWsdyNFLx0JTKIeFR/nxelGmyaeOFO
uBOj2fLapDWuWAnpY8YGZ9W7CvAO66i8M7pDpdp+BqAlOsynVwDP8VqztTEu2bMfuRZz5mooCjNV
N0kv2sBZkYDPTkUHt5qBHLp/Ei5/TViKuuHtAkYB0jNyNZ1qT5WroGjwB8nUdhMIbVqVOiQewAtR
v/t3ahBXWZ4TZLpan1X8kiSGWOtFOXBqFeGU1pZXWtcQPjwR1KSEPx2yLUwtb+UNcuItrrbB9Akk
L9R5bONTiLZvFb+/2PUWjW2hRj4qKElY06u7I9y49QtIu0FN6o3csTkbRBk+ewCL5UJNGn2Fa7hX
YU1FUHY3FVnx27XCmqdigOaWSLmJkHjMErqWKUJZpnNnaGYmfMPAc5yvMXgSvRHGFYwTHs+DsxIQ
W/z7mMzziyWG+pbgZPRWwdsY7OcPoFyC4YND5xTHB7Lf2EcmzJygX3/SQI9pRTK1KBnoGrIOtU9y
cEq19CSUceeKEM+GEPi1zIgHjNrrD41zOtwtGIc7wQbmAsqsSsWsBjqlUdaGZZg6FgXcHsVJQf8B
c5P6gj2yvvveeB10S9XhVC7RrSAyvjuzvwmFPiSKb3mharD5FzyT7MbAS8to0dH18Hqpows2yt5A
8HIbjcL9hitLydMHJ86/sKJhF5ebMROKrhtuyDpuhl+SqNGMzpTvFrvB5ye78SllN1I9A7rI7A++
R86tzvhmgHoyP5E4LjxNEJ5GtevqRnb6P7vnHTPvt8IZANGhChJB9alVBwO4tL3zrnPDi+vJBS9l
Vg1+ci5G6qOQRqKyMo2XjbaXeRSPEiKSVFU6HIx/34yTiKulGXyHV5ZJhhtCXTJ81r3WQW1OW1xD
TmHGx1zneSxd+Q20f0XwCU3bIS7W7AeKph8puYkrZx6dJNSwVLaHRcE3pAZPuIH3TZtCEWPs+9zj
JOTWuuuBcIIw82xyGAhx082oJMrnMOP97Nn9EXm27Gx7tePHpM7iD+Lx1+swzpS8tKE2Ti2UGb43
pIfgrhwCUmOnzQ+c/e+VzroRegByizNR1l0ZJCmdz4KYOf4FgLDy+LrPQevYf/xkj2SnnJJ5XihU
zWWUvnFnRxSeO7Kuvrqbt+HpAStIjhwBEVIqkBAXZ+EcQSRjZ85A0rKQWWnd592dTuqDSuMQOPmV
MemsWorxLQsz+Pim+bYZaLoBxM4f4MK8xzls68ByQ6sf1GlMbFXoiJiibpyx248+9y/Rp3Tep0Fc
3E6LGCSyYarEtCvDcx60KGbG+g7tOscbS41SlX8eDzSOMVJpGrtr93XUOIKVbud0TT5vzqgnE/Wo
ADYepoTQ4SKx6m5OKeVu3NAIhc/AmNXvmW1inH9VfKBFlS06Euz+rkoQvNNeZMAXVfx2eBYRFdDc
CdOGq9eunL/OEgAlygvCTZFXD3OhpJ2rbFqYppMMpzSO1+hUKWgbDT3ntDwHhcdwAwwMA6ekHCxp
ON/SkzLq1Fmx0SNIoaUw1Cb1kyJVz33F/RKTm2vBrO5yNh5hYSA6PKpSyKwHCBW66YBWgiiglrCa
OLxt1VXW3G4rPwONzxL6dlHt1Ms5hVkcveEYMq72GGCYLBNcrKQ8qJcWgidiLymSAbssZwke1h7B
T2XbZn2mkmtPQrf2XDro5mGUuCG7WA3tVdHsncjN8djDVHwVqddBZXkAH2dbVhP+ACAMTJq0qlLJ
ctAAVeDDL9RT+71RO+a/PlZ8or4qNHTgJ+faWGS93vd/JHDrGR8UHN7TgWy67UrIYnR9CLXPCuzf
e79rvX5HqQUUPftfWU0tR7wCnfHXnNL28T52eGbDiGW9rBm09WV6tMD1XDNTxoMzkyeQDwMrQoWY
6JwThMco3ux+b2wNzgHqBJNvoEV2NY1C7EsX5wjP/3lzdseoQTtVdCn3S3Qu7LLSOjQNTmekffJO
s6jXur7W0EW0FpdoJk3X3Aohc+HogroS6RComQEERktxguxxxy7ILu3rml7dzo2E7u/an8sA/C4z
osWbBS5REYlwnbX7Zo7EMo7caiLMmXyteyS6PapGH57r7CO0CR2eGFfv8sSYfgDIxMEE9Raj8tpT
ok4lbWBHVg89rpG1byMgXIV9qLoVyDQrYVkmJnYJRnHqZBZSqV5PnzLd1h23Me1CVgexi6+dy6yl
EM6nXvH9sakmg0ncGDRXDVmzS2GycGMjOQPRQ0EV8Rj7Z6gaN010PJkXJt8KTrX5dvv/rHgo+4DA
6RnlYAt4+ORrPg84wTyrvdly+vrxJFa4WVe09z1HCi4pFZ67fB1kvJC4Xp+hjmCdDNVxxONtYV6q
qiNfBtJ9BP4MkbnPnokqaGBbFTXTMol9CJxfZ2AmCr1facuG7xJSebgakQlq939pJIp3QFR0aORr
y7UAzLx9wirF9nwjQOa2zLZTK7PwZdkqi/JJKwEPU2lUCyIVMHUmjeMG3Mc2/eaXPjGE/2CRptzD
dioNFoUxVAkbOC6WPWRPBMQSfdjrBhc9bp5Xff8sQFlK652fRX8C/bZf3i0Y1YMNLTiMWkqEQyUP
7gHmF2gGZ6zIGQb8EXbqotQ/yr6TcsVhGVmOgoSsjG92Wph0H1GAGVMsoauMmVmMZm3SCsChxhyD
suWQFU7obQpr4ip/wr0fnCGdv9UOm6a0kID8p+ia6Tsn+XQPVrvN6wLdvjD77qwOpIr6DI31hDFD
Pa+f4TARSyBtiywJs55lX5XcgUIgVWQoJFWxNPio5EeWbG07Kc8a2mcxTYJvaxavQZ7ZGPfn5MCd
XN/OAZK64BZEEcLQ0k1HEFwFKafXv9FOIJOv5j16exJG4WXPOU9vS9L0a1qtwTJ8avorQx0NiIZm
pbDJX7RPsTSB8Ur6PrSuihcAceiFp4sBQcSxuTqwvvXXQS260nFRlL8dMcd60W3PRbiWrUcQMnl3
2ryPA2VGN0akwhNekcOe1brawfxNGnPIgnpHCV+TcC4g7n0/4txtofLMjZP0NqJVPA3p1RfyXJ1r
cuGpNJars9QAwu6XyRFNi79XfG2cpH8lIFx8Cf/695FEdmfN4R2dEPQYe9MQ4gdwIMoHPlvjT+Ke
6daaK1n7psOOFsMwT099b4dnYwxW2lzRclSxn2KnGJHg0SLVQJdqY6l2+NbqoC7nzq3H3Q13Wdty
lLi7BWf9Ql2m3tYPqrZC37Nuj/L/tCbjCOcCH28qsHSimbs6s+TcKNFL3tYmkyGubt2UoS6zXx0u
zzvifrHK8OlBbVExgKifQ3BS9a7UT9U0LNGHbbTa15q8BREx8GKrOzx9hpYpS+FpsSKJSvg6tkwK
9YrLWfUt9W82ApUQHF8ply9vvO+gYhQ8wUKN1Ycvd65fRAIgTH1LiPba1dkIaVeecD0bRl/N4ErF
wNOVhUD0bh6mbHsBZ7wLt7LTQ0Be9wdTe6pSNHp9Ul9vkb+bNsAvoIU+wrCe/uleb1X4k+PQuRDt
I9EQxNclCxKJk3V+SGIIN4n5z97lkEOsPYouyYdbJM94Y0T/xKEhCkSP29HpWd/yxTXbV3vrHShd
k9ol4zK17iKXZQfalCTac96mBTw791xuP5hHdq/bq4c7fsc4+ae9zNpfzl4YMwou8kkAJFlG+j4U
RaRbvRLOFYaVRTsCfjGEPQPtgo/zF0d9XMXiZnr2uJ8C4CgYRthEtJ5ERk9ZpR3hPb6RYRr/6YKN
5lb3s9Q4UrMQY0nMvkqhaBjiYGsIrA6Rb7xHzgdKYKvkUXXw/aohHqPDWHQ6wxhJkThQHy4k0Yqi
S6DD+VwTvzz7h94P0aDywuI5RjpKJViCaliM7aqlozFjisdEmRsBddZL3kJ/RxVPYok6SfYWs3e1
kqFgxa8cRYRZDhD4GCT48hX+SILzcjQ4KbhA6jO95wFmc3ORuGJYVriKMONA+wVraEyLfeLcsIFD
O9a2wtiLRUnrJdO5feJN4IkA/fQ3Q5Q8Oe01KjWEB3yaaFX6NmQgEJvaZ6FT3TsXTyXdtb6fYWZQ
1jmXGxiwxILzlZsDMeQ9vBv80WhSVZKsXXQ2uWuYNxnMQuOwmd46bO3/I3Z7uNPxWtb7uY8xwXmX
LOBENk0dFrXAgcWht4XmN7rftsFaLExe4olCvk6N6eWR4BN9pxHomsZQdAuZ6c7gB1R3uVS7FIBT
SgeE0d/3zUPyg+SOdleJWwlgVybrgP7299qlkONvqXKOq7QQqcPDfKNE0Usgl9hjHLUb6iHMvS+z
wJs7bPMIG2/cVl1Dl7N68YOwlHFii67ZvEMnIlz/45LgWxH5EhojWbQn0jnyDIo5I61LSlKLG2i5
dX43z9BvTSSTpydEXk8AqG3+xkNr84MP2NlhdntdIkamS/Gzt7VN4YW8nRdUDp54GbcKdZzOfGb/
voXsPs2Iuv5QRHF5dYP4ZDYLhyKQIVKJ7nei/VglZrh+i1rcdr6u8vIWvWWyINH62tm8vTpjYAb4
Un0M7RcJ8Iv5EWbIf2uhUCxsjkD1AFpbuTrkONHu8rm8LQwW5qql6h/29aTF342Q/t9gsLBjTq+T
eF7x+WR1wY6WoJioLCkrh+CVn5TNtXbDINOfaC+IutldYaQgrNkpXpVwOCvy7V8QDgivcanPuV+S
IfBe7XPerxAVA47oXkZNGR6bBJKiYyT79XVb2B3GMOK4YbUrHr3JEcIRj4pn0tOB3Inl0FdBzwp3
X100w6C/4ZUxdhAd7L/CnzUM9dXfxWGY03Ruc9AzymCMYpO9TK1F9KE+gEu/QevVGSlNY+Fsi72N
9urry1KCQULiQRtVyxRe+LBhGPvb7eLRLZRkOMr6yqTqEclAwlF0Qhb9suU+z7hFwuLBQrF9wHDM
i4WAsv2sQVxZPIn1q+ZC4b4yGJ0WnOTBbbqwfrjYb7YdMQq/Jy5AzxH2NcJACFnWGRN8YfHoYCnH
3iz7y2Pc9dqQxjKebjfoVZ7AYJkx9E9lxhB1ozhJNrsDgudecJsU1kDX2Y+f38KycX1t+Rv9B+Ne
O9PUquyF2JGO5auCatjFZO8bx+VKHiRgy/b/b2bO57/bP+1QmIjOrssWsisqYqJKL1TpMZyYfMI8
iwVcX6d+G60BOTHaTACR9xGvVC4X/muJYJiQYpsaBiMZ+za8ctCsiLETx5C+noXQUM0mo3jaUSMv
wWurMiLANFwrm5lH3vG50hWkJktz28YF/dslcdPFw21eFi2iYU1c18cAHaKwpV24LbMXj3WiIGfs
e1Lut8YHuXSfmj2VMQjuzR6uaYM1j8BdKeYfHT1epuCfHB4aEemTiUc9R1mQf/r0jx4mA7e6UaSW
M8UMydsl1lXx/ylOzJi9cfnJ/oqu8sOHrmWJmybLZDk+icaKjy2FF8igsvwEwdfF5CHClHmh+yKu
Qs7EW4EfbfHlX+imIZVtSiVJiS47FXkn+wD2m+qcT/sxUpHoxmBHcArWURCS49rTfngWOdXfb92L
Cv0vYb/U1KgMfq61e8fpnk6wqr+/Jw6QGlJauP1VRMm4fez+dZNjEbs5SyJUuA1ejL2BpNftwRkZ
44SLaj4ome2LPZ9MoPXlGQt7RdJ8FMcFMAbCOKdJo6BUhmb1y7Ob4Tn+az7QhGtLTHCcs5e34s5e
P46jszcSmWVzmly9ywdYdOCaou21uyb15/2IsTjSVyhKpRmgR4uNVlRFKRa0QRi5qbRoIBMFJGx9
V+8Z8RUcweQAguvDaxXGY6j2kpTlNCqc4zA59yJjVbDpcWUwHZyYXXW78O7lghxu6yU3EEAB9ogj
Z4tzeBbQM3Jpt64uyNYLkFEMaaCpDTfmumttwxi/jxJIcLwG/ku6ycuKUO9vTMgfVP12U5v2eHb+
k72D0ZzNruXbF8Duac9spI0X8BZ/8Tyiu5cnEZloe1VYItNC41xG+YaeRterw4NaBGrNg9gtsR6I
yeonwUbH7j0DUJnS0o/Nm2pA6q4No1zUDKLeyC9dD0zQZrbEuzbhqX+NXrVf7aAxprwOFBYHcMmU
Hv6t94vV49WMHVf3K/iBmQAQ0uDlQZCXZZ/27nb5rvsW71z3qTbFFZu+YK/H9XRBoc11Owquatb8
0c9/atHnDsfY10EDfgy8Zpbf5B5HgRhTBXnt39VYZdVkTzuhm729+5ADE7MmYBBP7KvangCa0wNI
OgdcTXKo5LnWZF7rlSLjdSPUjRBFJ/8XlhPMovFLztkHNdYrkHPrCDRoRbkqYx6QSAuDONtS93p6
DONFGQTXg+Z1O75gBs5a+gbpEqqXWdildYp00VXPnmiFGoNpGCkg2a9BBEnGu0rBPPiduoOn9pUS
RdSWJ29pC+8IfEqpzESdOk1KvzpIbUHDD8Le6lc7+sbqSb93RIE//HCyR4qzGu+1ACPX7wlfx1wW
q/LWt8OuXJShNxqs7XDu5ckKbvyfAYXIJYHRWcSbFHJEMdPEH4lpsTG0AQjnDb13iiYehf5fmi8F
o/1PU89EyBAh9KqBM/GLFqe5wzfMMxvi5nwOE6cRo8+Jbkzv5W7/NMu2wBwhhFtobHUr1xCa5ql6
vB4BpUOmHLohKwSRWBzQPehR9yzNBtXEa9YVXEotKFxcx7Mp6btaIOpCsBfbLMfCiiF1MWCAuMpH
pZ5TdiLUMm8KF77srOoF0wSEFT/FnET+je0QS26if6/jaqlv7XQbXHYCPEP6k1PCzH+lkzYkHp8H
/UKAbEsn9x0bz/XMICq3ywmdb5Wa3Bj3o+G0c3GicTmN9tV7n6LbPPKsO5q/klK+98JdnG1bjsBc
mBZXXF5IwnC1OeO+xQeQp89KlPGlTriluoAIQXjxWoL2LSmLGCS6NTZ37VKwsC6OojORog2JTfCo
L/SCatNsHtplY0BlQW//hZsDt+G8nyZPn/wqdZp7+2TVNrrcNeRvQgvu7OhHTTfosDbHOn4kPrH/
rRJV/H64OFpy0LU8HS09BS7vXwgutffri3LpyCGoKFXS4Wcqyt6fcVGwudaQkS+aviqMRV+1P5d5
vTN4pdMtUC6i3/vwYMltNh7Xfau2E6bWAV+L1yc4HWW9m4ny7Z/C54mvqkPiOfEnGSvSP/1J/cNP
OD2NCHjaE5M7TnxvPh+ELW9ukCvIEzfbFnKt10mPjWLK9B2Wb+01L+qEGzZ0eY0CL2QsJd/RfDTQ
39nxSVVcZHG7YewyeCyAjvjSOnB2e662VdwmqdS5WApIGcqIsLRVo204+BhdcjB8DMnx7N09wR+i
B7cvkRVDxH2KvTE+SxzkSHLL6bQs+e5MKl6w4fGI0tuDeeRShN8T2QO3QRUWJCyPxk0mPcF9hSiV
2yoD8JoXTYMw0AFaRZxF2B9LMTATJM/l8dPlPH9oLIqN56aVDmfjveoxJMyXBCAfCLcnebNEPqWo
UmcZEWcb9RrQWITZEikDPrvd3ARMDhqS5KA0XTRq6Uozv000igIfrRivcZQP8pIK7qGhv5t3/kYy
C0J0qhdeU0AqatQsKBZBLzS5z6ZisJ3n7S1xv1B+rZP7fYhEu/mbstOUcqlpbYdSR2t3gGwuOrpK
9beqbs2MRB4YPM5BHBbUq0x7KLRe08fIO0/sCJZ2bnpzlHoeViucY4c8o9SpzdpybAN5aiKdBGL2
BxxIyDb7NbWGpRI+J4b2e7q8ysRn/Ta9/htVCl8+K+njUMxWI4kq6M0CPGirdJzCWFUfXAdvkDuM
a3pII4laN1zjqHrP4cdlTBKDRIPLVI+BB6dNez/fftOrC3CpY2kn7x9AV16Ddtlh+49tFvYKbtyK
Q6R2h4OWC3Pwnbl0slt+Py98lhuW83+qVA7pST2PimL/sz9/s1ZVoCwuGUX/YzkNa/wyqzPMQQ7I
U8u1iuCx35YqJ5fZrUbjosJ8uslZ/2hJ5s4cuzbaEQkrVCTy2Kb90v1cvNTs/shgbhWc22M+NOqc
cO++vjgTwZ5a5XgZY+QOuaWbQOUnlgCNMjYBPDqHtDJBHb/7RGxclj6YiWmY2pR1XStzmmwF4kCg
KHc3AqAsjXH7QTP7YaHNl8OtLr/WSvjpbNl+Kk+Rf7M+8blURC4hcaHOrjKNAkJJYWg3NKCPrXI0
u26MhpxL0upraVyq23XpRCDOIh6rhwINajfyOIDJDysl+/kwd3H+Tti8cBuJ2bropPxfGs6VaAvt
Aki3b2+wxlkMarPHpdVGJNQqkdDWudurGIl+PbnYrHtEK06t2mPgv6bhbgoDlxbhfEUQyh4QGaxe
nnD9KfmupxC10A+ZexoN1HIDEtCxRXBxDlruwGBBF43otdZ56Lg5H/TmV+9hBl1HuXQBHlrUcYvq
Wk1Ipo1h7mzr2iMfdo0phRl9WJGcWJtkjyMXJWbBVLv6I9WywnyGQSNOJPHNDgdahHvc86OUJT5g
Djn4Ipb8LIBUkdr63BkE89ydPiGZDohFKnMDP3/T29g3vsLNpF2erAltjame5+8VCdlpcgA5nSYF
sTdT4KLcBMtt1nmQZ5e6edB6pDmyPOZvQQeSLT/klqJV3TibZZx/B73lJvPYppHjApjfqYybfhEG
+h/9z9W+lixh9ILqmwOZR59vd7L85txDzAf3getAWq94mubzoYsxoeLhxFWG63LS+C4WjjrySJdO
rJn5Qe5KOQ5WEVp1+QgluBhFRPOPnQ9cYzXv2Wem+1myv1E64+6LNTerz0eOsTMPIrRUIYMrHmer
jnyxXJT/rf9VEXMGU/xVuHzRSs16o/ElT1aiZ7N0LHOSfL2u5X/rQ9ZpwUYs8ZhDPfvpSwnsd0KP
UsXBI/pSTnhryN2eqeXrBVwVBAMDiPgKBjvHpVM01nAOCq0N76KDtWrupwctOYoJSuVIzljJ0zHS
X56WJDqI5eNyB3BXK4yMXhn2XjzxOKJOGN94Tpz72yEnZcdo+YLiiwQL63uax0RSjzxwm+tNvGgY
6BnaDgQCrinqoAHQ5O2Dc/E8CYEvhx+LzMjUURy3DaE16RVHSlvhixV20IBoszlYFp9DgyQ3IpXN
l72E6l2kpwKmvVCZz4z1qWe+IUfH4noLXyrzVH3JB55ctLlA5p8f+MR5HxtfuITFbK5aZ/9/6Fzm
utr8h/NnwmAuiuj1LPQ255zGpArZQnqOAwE7NAcso2+KBhX8c1tkP/6bYwc09OxEJkLDyvR6Pqr6
WbmXEz9adWwFrCOO9S3EmEHRsaKeZ8famoBe5ikhqpzBjkY2/Ea9gGKL72cM7bhP4zfalwOYRBlP
xuoAfOO1gQfu4wKUUj1VgsE9SKyICxxKwpIPVgmkBPzcWMqQNrtoFUrUdhIRaiRuHN1XUEzekL+L
wewOxD+GZ/ZZvmpl4+uesoCyN3kAgkmLqMGrUSior2C+Cm4gOJS0x+v97DHVbQ7uXM3pdzhjzyXH
CtO7WjIRBroScM0Lfekh9j5+KL9hZRMHfUfsnqf+uhTno+Fpna+CFAyhbDd+EHBcTkfM7vqa65LI
uJwfVW37E0clIj9ENtj6o3qexWeWdsQ5dxh29ksLLgmbDvQzhaQ1qi/AuX5iFRmiExNlGbWscowj
KBXLnAuXM5Vyao2AJXVbAMraJFA/PCN1CZ7tMtnRxMeG0DQ9H5419BkIssF5OMEDXcLtTa/yugc8
GaFfdo4d2e7F1V1LgBRIR/2hnVVCg28MphyMNNGsILlRu54Ac5n2PhzAwC+9JM+Wca7+4ryyNDoo
kjjilWn9I4YUXg4clq4BMOFeP7yt0beMi7MShH/631/8MhAaoFiJO6VOOZuRG1pjUVtaJx9Q9/tB
dROO78qPl3kVlzmO7pouR1TMk42kecI4MClhx68V2UoaLUr2mk7tQDAuft71SPOi45ktDFT0h7ej
oXGOnRx5BfG1N7Xu8KRL4LG+zMxdjAxhdcmaJrqlX2yq3fQMVE6FWMDCvQ83cn45GHYCG+oJxzd2
dUxWLGH4UQ//WMsz/W9m6ZJqHJ7v/YgxnSFXv/giOHRP7pyn2pmRPCPU2PTBgua1syo0CPFrgQ1c
iQTHZDnmnpx7fkFbSLOQTOrgktXVe6Wyp2wtFplmR332SWs6OOSI9zXPZS6gApoZDvhO+Os5xINk
9EbUX8bURcF5PQWA/kcnLEesiYXI+gSrHE7mS6WcbbTJypwkWyN/N0PKmnjUsU6Dqhdel+MnHbcT
6aMwk9qOWQNDKQ6mOvSqjBjciarfQDFP99v390lNTWsLHgENCzkJO7IbvFMNH3CipFwfBsjZ7PFJ
cZlSG/4yZshWqlDu7cw7mw9FzP8vu5WoXulI0KQHzru4QdxRp4DrxEqKGT8o/7l9O5vhyl5l7a3O
hsczuCNBVOmB/3WZ/ymW1FWr6SXl/W5gJhlrMmOKoT+LkkWYpn/s8OpJV8KUG7xxl0EmNfcdBiOf
V1TSxGxcj+0mKywdRD7+iPBdR1Ujsu+t6FCx7l98wfVgCFgMT+mXoFdwipBGv4GxNIfry+wWWBcN
0zCFl4JqUmsWEz5Cm3qM9I3Xi5S4VN2A8z5/MIY6ov/hhCZ7X6Ur0ykzabvrXNwBrP4qGd2lbLQa
mc2s8bNgOcLz7EvsecTVHTtn5zCx/Q30TcRVeTSg8k/UjIHvV33zn1BH1NksmkDbPQA3u5Nqjcq1
BqD9oDR4U+apwQX7kqcKJNLt5RCt4O9NT/zwspRrQ4yc22FF/h9/CAcxsK/f29tfkDVlRhyi9DaU
85l/AfZ8m3959s709FsMiv89+mmFbeXrjYiKttP/062R+K8K/6AzfIHXQkHJ+hPtISv8ldmwE26t
46WEjCwN9yAB8mTwccFlGIJPPz7T2U5Uf0faT97RGsxEZWTrMY9L/hdzt2K5yG8ZAkDyOu0f1XXs
ccGF525csIp7PbBX9r9KSpKIc/veAwMNIa84ZolwQ9kWg7tvVND1gBqDIwrZFK5Wms4vq3CSd+f8
AWGUFxVAiQarzpaZrkhtm21fjvtTIyMrIhzSRMzkQOnw6/WEMIQE3yjUh29TBo1uruHjRl3Ar+u1
8+utpqYYiAjnQgUHjDNMuK1Jr1IEDMT3bOIO5TJ9iKw7sZQG7a7S+BSBTcx0UHIVLAgSoqrli3nY
M5BE0Qkn79zzcqnbb1Y9zPHyfFcnbWCsQOPfROEJumvK5A7DPO2beARHd0tejT/B8KGwFtxfyO2C
1W8mf/ucxsmn4Gr7tiusRKcxJAkGLD2rsqiuwpk4lX9naSD0+wMo9evd/iSnZa4p7tMGSw6EQmjD
BsGgZT/HzMP4sQCfx19OuApNTgFvnrnRmokzKZMMBYeFM+rNlzlsnIst5GtgUb9MKhmP3aKl6jvj
SWxnxLOIoEAYlNhWh0Un1RNPmxgFhECRq4hxwODI8BE86lCVwRwofkAHGZQYP3+Wbzf/RC0tYvpg
WsqweHJkinsYS6XY7InivIqM28kJhld9WdfLn2X+LCTbJ/ArOBH9BGfPabk1n5VBLB+llm04EiUy
pG0ATInMc43WO3pitbbDeMpkFFtOuUUy0V6R9wmtDQN05Tq42dOzRB0/MTwAS37vYAIAwMCJmTeT
++duq0CLjIOLs0qZgmvQOxD+xU5WN1MKcbolr2bbudUdO6HxgWVkLxPBwrwEXgUTh/FBykt8UPnx
yYooHYaAjhwDCrUIhCSjJ8LpCIEag+eT2wG5QnC1/Nm3Zhyhd0iJAi0e5uyXefq1luQXB4oXtMpq
l5Ox2aPQJXlRdfbclIjNNrJzGXX8vq9i6iplMKD7m90bsyeEj4MVIkKf7xCd9osmi5fkmGQQCReI
fvk5fkLMvKLL1EcG7i9H0Sfx+puZQTRv1KptWtv5RnrzJCIJ9zZhbdegkpLIQ9rfWSYM5A3KZCbb
8b4tVrSpOkLxiMREMAT+LGK7kQSPO4R0k6XWgXwQZJr3ZTKW5YxrIchKL6IczroSnjplK/Hoooc8
utbwkL2epkUmyTsXBP4A36JCATCEqv39YXqoJPCjxtoc42ZVL4K4GqhWbHPuA9aZDktc6QnEBFj5
3DKpxNLV2kNaqyN0iYwkwD6u2ZHMMB7c1In2fJ8otYYXfBXdBnkYC/FQtQQmHA9vsbpxRsOqvlAm
rKq4+O+EOyH9eDCPU8ogxEziNxGOu6QjIxBMyxXcCYx3uWNkWioCGfMl7/8fGwnJr0BnYvNsYAbi
LzC5OFaU/0jts5d3Shm/+JpCwsAD2gwEbn7C+LuGK6QflPYPSr7B5wpxS8I5NE+vVeZCZo0CkvnL
nx9Mcf0ykR2qL3hXayffTwfuAs6t17xP4CBTKwJTR0Folmiw4p5cYiJyCZbXgVitqwU1A4sBoAS6
+RomLyZyn0+dUa/3P01QftlLcjq7vFiNJM3QOOsXPtJxDIdisD+tIL4yULvybWemk547Aj7uTsA0
a7+OsCvO170LSHcdzJJvu08QIdwBG+OllRSEsJb+MQABJX/ylrlFEb2vAAd+fKd8uipAl/gRepIo
Xcxf14PjTx/IIo3JOXTejSI42/ba7xeV38ev7rIKBbAyX6vttFn2FEnuAfvSc0yzThn29b/ip0+J
kJiuprX84Ji7wKH7TpgGI/trUXcBtYUhL+h/LW9oGLnrXEHzoLrR1fLV0SPwBpS2ifK1avOpqpu5
QVOLxyNBhN3RHXdjNRlnTaiZdcALVAekT+qouB6lXuL//YwDtB+NYBxvi2e5TkKR/OdjNEEBRF6D
84KlZ8JfnEVh/3bO0utOiYimd9cebZBjjMsTPKVpAPoB6k6epLrS78nLnvtZWEiK0KKfBJKAJ8qB
eFjCSHZhdGU2zX1q4aAh7Um+BfSwOJA9v51v4fh2Fe0+Zj/cd09ToRRvecYl2om4ikcfxd2IltpM
ujCecwit7gm5yNWCtLvpySq6eY5GmSUORBslNVUKCtLKCFCWcZregtHYNp/wk6sSfKuLM+Lu/zVE
RlRc6cHXLhSS2KH6zHUQfc8/EnaEoYk1WQwjs/qCFUO7KJjQZabwa10Je4BcByRWAY6lX+kIFxJ9
aI6UGJk+D2tC3geDbxz1bwQMb1uO7vBAlmxP9f2IHZ6JiJ2RFdqXVmMtsVg0L8GZBSg5d9P7oC23
lrSin8XaBw5EOBd7I6FXaQUsF4o2aT0/shaA8PzeJHfv0P1Ou5CExRtN3S+CjmTRfoU7SDTz6P15
fh5N0u+utI+v93B0rVvBqjElEXEAT4Y6eL1+1tQYhAaa/qF8jzIDsa2lmr/mfcrlFzc/8O9MrzzC
86rgl7rK4XUi12NOzNVOamJnWbcQoLbY9oQq+L3sLyFyTeN+F8xd4fAQXY2+nX4LKVifPWTa90K2
w/WoJlEQDgnQgNv4mButf56UbishV1d3aC1IYgti9V4sx2e7tHNr7xtxqStXODpRK5zvzNqnyuq7
LrASaNMxZMP3fWsgIJvLtus5iNXmWDXtPPkquZr+JEkgW6Pm4sKiJzXcbcmj0B642m3K5OJYxAcV
w0WB6/Je/j4sIaobrBihEox6i9z+Fh3MM1GxSZ6iPkb7Iz/mgEE/FEt4iGveHhA+CxiBt0+vySUG
i5EDAjn+3GfbDN7jdhw5TGpG6wWxKo4BuHKFJZ5hCkLaZxm/s6VO/getbSzvP2QnYldAjw0/taAT
0fyUl/rjh6VXrSzf1ioNiG6FY4Eda1FeoR2t7/F6ukGNBEe3C+VmweexifK7OkXui8jrVga5u5Cf
yla16jJ9SMBP/ysu6cRHdjh2YsQS+6t5NOwjG1KL+WQGlZuWUK9SQXmbGAPkfLwe5XsmQvqAl0TD
jha2jVv+PX6VjvuUVMtprwgB8+3a+zBalqmX/TDq0ryi618r3lK+zuk1cjPBu0B75YJORzMyloOL
lDnBNeJ7sTAtrrzN+JToZsi99TXfCPLCz0OghDpCzFrpcDCYjAh5cImbwhDdDB6bu3sSrq9ZOxFZ
Ypbd/ZTRwtbyU8HYS021VMg04pmWqCzgN4YLI766yEYoEzI5wHL/VE9AETxlL67a3QDrqvM/3Q4F
njsqg37PFvSsHDzh3CYrfR94gJK9Yldli1kJwFWVGs5QfL/JqRQ7kKc8O5rFUdFPfxKStyCosk1r
+xSzYNlvazgrKnpJx+6KZc08fmuadq+VV8buydbrsbwaGRij06USD1pR6IDX9n8QTNaZN7AD+dAm
wuEzKuTrkoakDQdH5Y+KTDk8Se2sa0HyWIT2g0BLK515cZ6/Plf7QcsncJeqNlqheQP/gUYNR0uJ
enAcSftnqxGhrScvLS2KwTp8+o+yFKwmkiZYYtAEtuMUyRshQouEwMLleMUWxK7fWcTbpfJozD0h
LlsMG1Lyk4e07Z223e+zMGlcVrgmr4bILwVF6RCdxXYssAlR3Syx9RBFVgyYKA4dkrw3rsqiuVE7
OTprLRCgd/6007w1y9vC5BwdtjXWlagDXH9hlQBTVRLtq4w80DSsjkqrI+RkqyDgOyRM8IRVdSPL
2LXlAONRj6QnOfvUWSbOt8JtiqRZI4tqZR3BmTggNmiwE0aFn27HsHL1zzqB6L2ntVIHSYlfG6AQ
L85P35Km7m0pxmnBngf0YvYQxxNppNOwEVmnCAxjIC7h4ZYS3LmXdVAr5SGRSXpwfzObUEWYCzJl
YjlMYKdzZ8tKd0m6ZD6/nAIlnfn6ZgzogfZrweTDOuqczY6+2iBgFhf780JZRLCooMBt9yY/PpMq
u/Zqx5LXICoc9cJNTt2+PjNKMFSSou4BVmGw05g8z7ZS/AcNcga3XHpbEJ157HdwunXM2UW1xYqX
oNO+nCMwydArLnLUNjSfzL1ZQaQw3vtQKIJnxGHlWiB5HYyoBLy+Qu+E5tB9FLz59BliQdX2DjXb
D7jU30lvUTTsu2ceY6VYufO0WRCby2VWukzRE/z62Z+EET40reUWdVI456YkzZP9hbuuoM83kFUF
ph9BiBH3FTmeiDCP1uO8w56b15O5dDmSmkQtMkyLlcuotP6wKEFVyAvQIaUDBqISN5fLwKrOQSHH
3yqal4kQtPhLXNzt0HM8X1pNuGoqCz4tIbb2yQkRfWHr4DS08bCx6s4Y4prGc1fGhgnjGZimKXB2
/WriBvficDJ5XNjg0rHXudNgzpkfKisYoHF+gN5+r1JVy2y4DRtvxdcxbfo3iIWXan0zjGUT/fNJ
fJPOTEMgvLaCin/IsyflI7JUciSgjQp12ay6gcyyEgxj5mal5PR3pOwD0vAinLpiyPML65y3GWQh
16/q77Bbe9pL/13g/JBlvOXnVJYcj2BXpcHWnp1TjwPDpZSIm8TdMyigpawciy1pISaZ1wV0ti2k
OEdCw4YvhXYnn7/NuINgMZ4mbzxRg1BdyX7AiJJwn4TrsJ7TsGHBYLoJLxhh7JAYsQtY7i6Yb220
5PF1MzHBolEfa/NiUGnoTdSqqmlz8GGLjTEXjy2RJEdHbmZA6VROCNmkQDg2z9Q/hhGr8nl4i2ZA
A/cuuRM8CsvT/ugs2wUurqpkBKmFOS/xGzoA0SrkznCK0b8lyrOuQjxnZfWy3vPIpUH1khVyJiXy
tegyDVwiRfk8rAJRjjGtXqXMFRUeeXMDQ5xsDJm3p8++mfn3YzJ5n7P1c+NvUUwZyFdvNaLVcsFp
eVV/BnWgzhUxKZQu59Bpfdqf2bFGi21ZxLNuge9cqK3S9jIWCEoMggRtN85Qza2D93rUAw+bkS8W
arw0adG7L4qvArlp1WFjnHxMOHPMEVib4P6ckQDCwoudKrYVL1JKdWVjMi5eoR6k1ap27UL/S4zn
yGYgH6VwH4MFOfkphFK8wL7ySS+mnEhyhogsntvhK4oMx5mfZZYopOc8siwjIo7gYp6B35nLTV8k
1lJvswj+0YUq1M3iu6OGXJau2u2K447JT3ruqGOYCiU4hFwD0WykSpb0zw3IO1AUCqEGfZSM7EBW
C1bWNYDLftRzLjck2ekiXa+8R+MudEw/oGz3yNAFzLa4pOtDJHsowu8ijWTZMvRSHweH8L7U6n2r
C1U2JNBWl7+/Ld14ZQT/6oSA1NrZzaUeb0MkCLg/tdVrdS5jmmkM2aFGY+kJzJ9zJudnmnPZmLos
SqJqw8kLWU/CgqAuCn3etIklDmpmSAAzDY2se5bEyGrkYk9fbvv206La7sS4cvJMipnn4/dqJdIA
n/5tLdfy+SwSSO5w5JMBSm2LGKmXVvIaru6vo2r9ittj+sqcvbpYr6lD6HCd2uewv7gRGTXXG98k
3ItoB1FjeYPycqf/KrsbtYo9WacM1qMW8pN5fqNuKjS7disV6FHBj4rdALoLJBriMA2J/ZC7/yPP
p30QoUQLarAeHYJ2+nhHhY3+pE1lqFkmbZ3CJl95zilrB2aC0mzD7qQ/k0YnqkSHAB7I2/NcVvFS
3q7IdkBbCWwMKRapxUuj4F7P42OQHxdO8UmuoMmmhge6c5jhOC83yeFUTvZngbf0/OBgV2Agr0LW
1ZvfsCX8k8sJ2koJu/QBb21Uftr67ZYdUWBWj+dSFR0FXQCo1cVRkxepmOT8npB2oHwVowlmO4RY
RgEKmWOqqoVRwzeI9W5SHCn4A8KLc93W7mzRYImWkzm8OOcwP6Q/RFgAOZgGD7904tGktMYxUlAc
i9fnTEi7BwyGuE7MqUtJzObUkeoiBhwtV6nsdcxc8zQYizI3RBKf8/D+IOz2JGACsDSaJnjOooA0
b9qY7UHxJDye40NpaXSNrGz0tcsf0hDEct8fDVw+y5oxdYNXSmPH2kJRiNz16wz6dlPB8p+J0yh3
L+e75XK+JHsUNVuWn+IRWb7eXcqBRA8taC2sQFOhkTq+zqPyu4Y4LOiF1Z4x6WT/ZUCkjZ7ynbiH
3Jaw4oq2nwYZ/BDXV+uZY3uyW+huri5ZgxWSq0tLgSRm6tGze3cxBTVDqw/3CtBTuHdX4aiqBdHO
9pxY86MGXi/w5ZeUEtmc08Xg0KbsnS9hTEVDx5i0q6zhxAQj0+gPv+QBvWSxyCD832xVrdMPbKnv
c1g3rPvUfo9qotJbi49jXO3ylPwA94uqQiFoqOd3VUhnVxLBjSiXbmFEbjjcDL0Wgpmmzh03jRaF
VBCaAI+GMR4ttN4rU8rIQCTcoN08hFqTCauOQDkjGHvjTL5ClQk9LddBDK+OjnvBDABg/R933y0r
orexvMJNat0ZJgroLO9I7b53PxHprjZ5zppFTp2EuRHnRTBw0O7ju4r+NTHQFL8FNRT0tBsqwiqh
0G+HpkOhf0icC04nUav00i31dzRLtiGSv8l3arWC3cVgI7Bb4VBE2Op6bhk6NaDP656v+9McCE/y
XF3YwwKFsW7R6vO/6ryzOqj6qZJDchkY9UJK/nejBcIYJQLwpP6Yu74qqA5Sk8M8qbjpQAXRhWXD
0gJkdJ2zEKhO/jogeaCD6l0YsPkdfux4Bs8hoFS20aJIrnMxPPiTzDo1dUy+jACs0zuJlxyaka3t
i7GE2P+ZS/3AZw4lDv4vFLZLO5a4ZVzFkINphh5SzU35W+toiTeMRVVNsJHNZLixKfcpxbrJSN8L
x9vNiaxDRXCAHz2XS86+ulXFUMuu1ADAEprUVYjqc44KYLwxlY7tZ5P+Ylsr/8xy+jqlzsZZAeki
g4lALRMufR1bY6g3Un+yVPoHJKHPWztXqRaBM+TAF+ZbZ6gXOrPwOldG9c83KauAjr/yL6Bc3z75
ge6fuFB7lSaV5qZNx9fHwhLUVpGBevd7erRoY6Z5RETDcjZGZlDg650ZHt00ZjNMh6rKahuauTbh
5f01QO9LkAgJVjtj8oyYkfeb8Ri+lrGpjvv9LaAnY0SeMhuw1ePdLIZAYt4l8hqAFqTZuR9Qgdlj
3biXbqzkDT5+dOBSnTdZbdkC68+2Ijz6JgbazB2g65gPjBWe522QwY9FPIp6VIxC7SrmgzxMnW3w
0Al6rW640qt+XlQS9f+XhA0D0ZqTZWdIWgxI/0YbzR+XCxuQBUo9ER4AHHzLXEvHpuEqPXDxYHyQ
2JLIuuGXF1I5C3c2KH+puzwzykX0NTNaqE6SFjW5MIdWhOn6iaYPQF9WG0gX05q6cdYexny99ZSf
Miw4n+545s1joWfLbMsTau4v0+NHxLNIfG4rQYMJzZR7m5FEcs1oUtlVPVfLaXwczGNxiTTg6a+1
z+vcWYDhasstqjG2n8t96lJk929KomckOtDgvOBB7/mZEGuVhommcxm6uwJMGSmkbKtY3XyfHuLm
6W7xMOJNe4JeDCDxEJCrn1Z9VKJ5NCHIeOpVKvay5Ki1nws6Dvo4lM9TBv+8B8ajx/k+D+JrvJJD
SVBxHecfFeMQYZSevOFGRaK8HedwU3RCIKjRUr/Xw9ltzZpQs/ICJp8nIxngL3Xc6iJOBGJaSGis
bx6yTZLrTOIh/7XwIva0IusE7FPxxMQ5PCeEVKJNRlb5R+ict1NyJ5t2ZSzGO/lQLZY7XTiM0K6O
q0FWKYtXsmBGSRh4t4U3btGHlzR7k25De5yRGev6Ovu7IlsKv8/ljq/zVxuiAG8Bb5UvalP9GbgW
r1F3BIa2yA4RcAQph35UJHuX2Mjhl1dQ766py6RX3lr4Kz35J3EqaAFm3kTIfaiv7wCMa8J6E2Lj
plrnCwlDzeACvIvlvfWcftvxmoaLqSmzwRCrc/NFP3e4A9Q1UNI//dOhJqGBc3PARwfSz+1BCzJR
N8rQ/1eVQHNkJRm3p/3R1VhkRseO1dyV4/hSZHn3LYYKUWeBFP5gz/Bf+KMtQvYfZANqPMfogE+N
06H99rJV7Rev+WwgxFkHMlThOmCxrcWR9RN2uA/otyCHXP3SKhPpGNrLaSaIenlto2VVEO2Ty79H
klzbtOC6TXFYqbcK+VJGxFDzrS2f9y/yEeOhmH688pkYxiQ22YY55FgWiI9F3QjAmC4c1GztJoFL
Gd0fvfJQGTJD86EZvA8FN2AK3ya9CWkouFAquVOxi86Xru8dm6hOo9dAhDKEi08TqnjqCK2kUaIY
vPKtCRi5I+Lh+WfOuULAtRSRwGnlvj4JXHngCqo5uhOujfG/IDayIN3Hpt/HQBb9JYZk3k6EP+qi
A0k/vBrgdiKz4Olpw/8rvy2nAa7k1LKKSGN1z0PjiPx/VpBC43xDuolkKTYDs3uyu440EyIK+Xf4
iqDZVYsueGC+OJLxmlXmbPDyeUtpA4lJ1QrG2AUQLv6FQYFpJH8jfKBcc5IAlvwYk/wsb3fUQZwV
CfXkln35EngJTICu1tYu2UYkEIH1L0wP9Ha+5peVKsBJqSKvpp0PqJo0WyEnptFmKGV2h9QH5x9u
NtlfbG8byYI+1fphQbqsJBl9nq67vWNhpcN5Niz0VV34JKYKemMeA4159XxXWIxJoKlNJyosXO82
XxgW7Dk4KYU7qxrromHd9RY5+c5s2N/gaQVkICCikkO7g8bZl4nDRUhnuEODxiMSqHTiPAi3hBbp
pOfTXKvkySPpHcUnUINvoHEEUG+Wrq8v6VobdWhFhyDBQt/5zZK8tvc1XX5fCSrAj9wJJtFj98Il
0pvtuetNFqBkvA8UpTLmsXaE0X2heHBvr/4zhbSfkiASiDxrgkaZYGHQmO9P6g0ikNcYiqo97uMd
PzWEWsMuUT8MLCuNmtuBYW96zRddDyLeub9WplO8yQ0CzHgKno+TZguXxFPh7kc2YNyk0Bgm67lh
8WdsmTNIkrRqupQX5dcjEZAfaGqDL8PQCgVkFQqiSLl8EZM9eZtXPyGa5WxLPEti7M3lBvYznP9e
aWfsrrCySeQjomV9DSuPfjc/2LadK4KmtvAJLwyJjVU5MZ39sLG64SvCpqAewM66vs2jpp/gu8eb
Jklo5yyEbjayDkbd5e1bsRpNjW/3ayRTzWLSS40T7iz9HaS6BNEz8pUDBq3xvUhWwjHt81F8UfEV
ISl4bJ0xDzq/J8CvKAluh0t5xZIuK+kMPHQyPyjARiLxDIlhFPXnNg/06COaj22e+dD3IqKBVY6R
5S+6O1keR7OufWu5wZwU8llOU8F8UM0lEo+9evOkza8Jat486l5QIFdcamVRRhfSRY0mbZ6DZp3J
9x45Tj3RxyFKkGsBqDcc2I+HyV24sHtxIiVRYZmvwVJpxvZ7rBRGn2u7C0HPRPcDgyj66AoObSWU
B+OHScToGz53HCdxXvGDcnhfnGkMIB3nw6xBQUw1gCgvm8Jj5z+p6SIJHHmHocJxo6Splm3Ad3Ft
j6hsy0o3FGwwTJoMs+jQ9J/OoyPwsKrzAE8vrQYsFN9hgUuxQ8Edyu9c24EL2i9cP5s3CvBJpqig
KoC2YsJJh622C55OjyfJEUbEO+aICUq/gxaHYqVT0qN6k3H8uf3oG0fUAqx0HyjVizfTiciClcSK
vvgRRJLTkUfTaBXsMbLIdxZp39NZ57yLcYeQrfboqVeyQZG1NVE1sRjA9sYrZzP5071Ls68Gjf3Y
sxZdZsMAk/EGdLa1czLPdnO76ebyBj3hfadGGWqYfeOXUcRpbnSoHoYd7gDeaAC/cQ1aKQgl/ozY
poN/bjA7LtN3COB8QgQf/prCveDFoo9pjMIkc4PWizo4bCvDLxp291rgiCgOLfL3eUp2cni5r5qp
Op6AkOwKZIFRgL+dWhwoIWf+n88Vsb25xazHM6H5/IZSlktrjJTSflGAQf/uD+QKvLzwOz5FOzFj
3eg+t94FqRiED9bos+DfkcJ/DmNMpSJeNeKF53ZqgVvqmErxbRcKoqz3SQAUidx9IcRG7GviZJLH
d9F0zhqoWv7WsYkqiQvtbzwfw6RbvYXe+aQI5V24iH96C8/nEKFal626UOlkc+wOwSJIe6wC2jX1
Avv0mAN79Z8kn8CZsmYfti81Q4jxumwJLYLY1mgH+/EFJCDq3EWjoKA7WnY2wG/CIWGeHzWkQcqa
jWOe09CrmjY8cgZcZKPbFjPOnYDhqnpTlLdyyj+fViT84l2mJJAJBKrGluLT+frBS7fkkg5a/+QU
/CvJBdljcgL+YQI9rAs+s+eSJk5FSGVJ6VoYkUdp1bh2KggksrgwPCUagjvnQ5YZL5BTPnfUu8ku
z0eENCNITWyUDJlxKpv9UG3FTM1AuVys+KEeiNlimJIJewpX6rrDgFufZofLP3ehoEfE5HQmfzoQ
y8m3w24L9iwcA5eihuhtYKxHrTgGk74pN4H64qC2eFHEtmBRwc45K56QGk3jEM4fPcpeyAyxbC42
6GbXHVjeIfERWMvt1eUKTP5J9wFREx++4iEu6QxO+RbjTf4e+JKrBwie6fEOUW5E28GoU2b+qRs5
tQBNgqW3ecI2i03tu/vv3iPKrM76k66X0CvQQGsJgBKg/ns3ic40G+tcBS8hUzVG6yWFhNlrLRCP
IHu8JfrYv2xgkUYBygRR63RR0VL8IsqHbJHROGg7rk3M+ZH+5iEsMGb5yvCHPFNbtxqUogL5BVtJ
1mZ8ka6+cDso4/plgyEkTD9HVf3Cf7ua+RLpBMEPcTJJybZB+YXZPb+W6ijCMMwpnbeeWxZdP15s
njN5wYl8VFgeKKtnkxXosRYtnrGEqQvtwUHOjMC17A9f3q/8h+NyNArcRDsJTbplORBayDKrT1L7
NSguNa32WUdVCJdB4GOsPMx7nsMqvLFbb9WKpblNnUTTLpVjhNq7E5VPmtRr0zoyxvFqitoXRyzH
VboNchud/i2hSkhwcPnmiBMkl+RD3O4cXeGpRk4sd77qWR1U8O5+MHR4xO+LcERAhMmNa3FWC6XP
QNVWBvj4nO+K9ku+Yg4p3/beuxHGUtX2K6BfILY2DTFLdEjw3/ohUOkvTAk4dAH9WWmPz05x+Sdh
X94eHhNnitC4p4f3CHBAbI1BxHZIerCtkBnerJZOCkC5VLGoESMopyjzCUg1nnWq5cRVxaVGwfB3
BeAwesiLqDpIJxiUW2Taqk+Y2L/ijC8vcb+AGm8jjUR8+lqDTNxZBYXY7gZmJjaACe1MbErNXWq+
5wQdfpMCQ8ZJ5C4PZifMjyaMRel7ws0feZF1H2SXwslI0gpKz+L6ImyzZopw2sbClK/GpMGrveVu
Eb/inaN8f6XYBdgvZG78EozgrKic4LDKJwaGfc9yxeb+cmYcQBeCOTM696J5v4mu0VPBxVmh7MoM
TQ5JKak5uWNfxu682SPeHJUQp3hIhwPmvbvogFwzLCPG5IH/5e8bPeMDAQdxpji+3O6KVgAd1Njg
tvDMFOqfuZKVCW+99tVd2/KgNIY2eCvXGmXV/iEak7FNa71rhGhP3mPoXwHyfLZgXTDKtO5He2Pv
QiRVOaXijdjfl7vAKaFWkOlAtAnxZEGipN/ctuLC71UJpr8y6M5PIMKyp+kbsKlIr9SfMIMTV5BO
rUrSJIfKtyaBddneR/3v2vtymDh/lziZSA8sjhFArs511S8iHk4XmbCVYg7U9qDVl+R4BKzsQWEO
oUAAoAThA28Qs+gt50jw8jELffC9E1bSPKjQBAUxaD86QkloW9KkyyOFv4L3ZgZvMpLElswT3NrQ
6aZT9KU1QvzcYtsoqm2KxmRr97/1L4Yd/xcd5VoRL69CktcAFr2Nq+vZZXZS2KaHrTzIVv8VKn5q
r+KpFfVGx7EgLnAknU3EDqTvb+6CDA0HDWhd5daE+nSYytsF538KT22XzubutbWzlBQ2SMGxeLgS
RBtHpUYyb89rd2l3ti4Ql3dmX8fb7x2+8ES3Fc9B0qcg8Y12J3fmXhmEfJRpzqdo4JCwxsKtW7af
4CUmTuljGeQM/30An7MV0h8KyeG4nxu2OToT7+mgARdxGrlV6PqZarCkSLg66U4bTwoBhQ33F2sw
lXfVKu+CajI+BuHPDdrzfAXHspxY3+8f71IlqllL/al4lauLu8VRXxiUMUd7d1yMofz7aVmFeGFJ
F6+8fYZ+SLJiDjYqMwnAx74jX59BpxksY3EiR29qNxuRFBeo7aKFmVT79Xy5f0F9nw3FB0bzSKA7
sLwzpDjB7/DxFeWx2u687ctQOgeHpQphStl3rSk3PedteaAfmQTjn9myK+Rd/5hWpdkBeon8ODfy
pbJ5ka9j/ZfVQ83ATOF5dTNSxVS76Fxav+WmtrEoIiaN9b2E2oH1634gnposowWbP1TB3IfQo62R
P75pP0AC0D+dQ2LJkhDuNsp/UFePR49+59DwbpTBUCxgG0DLK6KNc77w5JZKz9INmq0w4BpM303p
ruJh0bScbMmPoXinXkcchObTnMl8X/9Zg8ftEaG/2XdFxVczz4er76pkhzP5KlqNbMzK292Xp4Hl
PsJ8M5iZFaxECErmYtLhAv4n6HRmeE2nv8MLF64IS6TWlQqRn1aE5OJDh/RWsmkmHr6FfSU4lpoL
4LE1OSIv4oeYnUINKta5psrhZH9PSRw/BEOg56V61fKMjUTKjqskY1qE8uI3PjlKUGnjSokPvhrr
P7kGUqq+w5dCsVfa/a58zK9Ih2/KUsoFYdYB7n47s8vZvgIPkvn4yPafYdq31Ghf94E4B+OK/JRZ
TBONReu1k/xvOgdAUBgaC/tml1AkmLMooeam5ST3Nqq9y9rwMv84yOdtZWPjfQfeF8oVwUV6gCrH
e+6eN51AJ9pFdFjg7LFrhr4IW/o6XanFFUVYYNdzbf3e2W1w25668P5sDAmsjfve+reb/NNY+4Rk
cVEYY98JKfxvYvvqGiMQrclejg3scyXGAf2OimZmKklmnQsKAPx8HiKw9esRBR7druIyFu9Wjov3
SXrs/ncdgoBY0EZdVQ9sZ/5zuK5HhfFoYRVIMJvKYDiWQ36S/YR79VgDU8/+yiveL5RAHAWRzCcE
H95pwS1Rim9BgS1FZG3tH6lbZ7vDAFOTrHIkENoicV7FDC2fXuxKznnpNVgwkt3LK+0we9wNFYSH
xhGq+OBHdHjD9DC8xGXd/lcBMmX7bniE071MBifbD0fYk9G3lDBDVh9uzI99urViZZ/ARd4MBv6G
ar36yOpbWfbMW5zXZC+5dawH3Ra3d+G7qcswc0vRBVlZzeww0x6ZgbA1yxZXZFP+BFh+qqeZQLoe
5sTnk4bnNHgQXeFNXNm2TAdyx0OFgPfhLdSTrnK9y/6GSSdz7EICMeag1fGBhNXuedBIwocdAmib
2GZLWSSqX+0U+BJMDCRhW8cmZYaOPbHp4qSDFyCkg3iK8MbiLtlB89qn+MOV2Ma4SelFZ+5MrjxD
qXv4TGDXo0RiCiW9mn3GanRnD+htnyZ14ySXiDkDBT77YLPUonaTvqoeogkvyXEojznYQku4D2E3
uJJTVmBQLapwUdSSUVRRfBsrNqrdlNqaRNaI8Pth0HuFKxxk+stMyW2wCAplEzlbynnTX18QrbZ0
AueUZEDDQ6RKa8WcX46FDSuPjPIkOVrj7P81eSJT5+zRwcSCOU8IG6HLQiAQGD5ODyfZwyvsnib/
3j70cqugkb6A4W57GGGLWVb7nAkZTFkTgj/Y3FeWC5JgW0TfFhJEHlAvd3XW7zlGtTweuAQrFWRU
VRwjpbIHOqyMWjWXWzjcQa+wxfALYicNT20ym+dQ4nback6H36NoHy8dLgFXzx99HPoDpj1z+BdG
T1Vr3PU9rQvcvqNA6yf9uTA67ZKmPQ5zD65u6L5QdVzRje4k3rLH9Hk/bmggUpqcRHUTHbuap96k
z1eJjZcPSSzhiD0webef/PljkMafXrAaJkUnNRvwmhHcwtDNL5V1cHjBCN+TTN3bydZ0zhLnMlJ/
UYb7ET7UzqpTcLR22OXP3iZJhLP7i+f+/0d5O2kRWYE6Q26yqAeF13tBunFX1VLlSSuG1HE6Kohe
ipxE/xK14wCVZHUuXovsUnWmQHkIH1g8Ghzk9zn9VLGe5JIq1i/GbMkjOQO53KlwLopll3/F/6Lh
3tx+0+hB3DIIKhp3jC0OaFab2Xzf/OAwXXyg1rAJK1l6Lnn2nT566zq8Er6kd8vbO0NGiMq+s0v6
dRkKoYDUQz8G1iuZUO/L9NLvDM/o7Cx6S95+UDlsKVPvmtOzC+eT7lUBIh0hVbJTBVoYPOGQoGA+
Cj3VJYMWn88ecvnIUYJ/MWvk4ZAHKaZatiGamLiGmXEXP1t/J/978ElaqXe8V8vOGN4btpqPmmiy
vze+bZZV8y0C8T6iGuJ6O4ix55zRPBwOijiBZ06Aaokzr8Z77ee7cf1H3Np34RAwgBHKL2COlir6
En4VwPQ7cUM9rD5TDt4ik/GjIsttSXHunU7GevpIyMSlIMEdurT8mT3Od6TpxJcswfd51y2KMT9d
ftsT/jEx07bXltDKNsSfkm4AkN4dV52sllverhgdwNmBEMd/2LiCKZ3rxHrFP69x7wdwZrAO874N
q0Rb900M193Mdf0XhnAeJmWesIlTXTvb/kJCQ/pbdbsbctEQ6MAsDy4ffLrnZRNW6o7/Fc5nFtnE
T0AklphAViJafBjorYuLCiAe6+M/woystzKp+wOGglm+BGtKcL0APbceAOJJ1F7n040qFEftc71z
Qv7TVSiuuVgCbbrmb5L69jcPnuJriOVuVJjCtZZHAG/BHfgugKOs18EnuIoJPd4N5YlKj5Hd3y0j
QJCGzAw1fZDbXOnF6I+SWG85OYIs23k/S/FH2VHbGYg+ySHm2z1kw3pOobXDmzzd0pfaOma8T9K6
jLyomrLKzQKcQJJ05PyTt9j+nfZAvBqm2vxunw5LApkx1GbX1cuWGeoahVp1DDp64a4EEuPNnxJH
n6CXc10/BrQWaswEAFuzxBJ86D4bNYRLVLjTgp/Yvu1fSVfFHBGF9jW5yDwtomfREXeTmPlX4HpD
t2bSkQkS2ZBbNhYmxnBA24Qo3pBOqVC7pCACxRoU+LHHvHLW6GKzpTeFUaQKgoDh+WPHKJEycQ9Y
5qnCgrse+gs+RiUu96+OY7cMKIAkVDERt//hD4LeBfyMy1xSzYGHYIVsoX5Ieyq1Nr2hD3amTiU3
QNPLoJRjtgb8GLccE3vukb5I8QU/LNV1q/3j9xYU6Vd9Swbe+s/3fBIsxgU+XKpkMqBLiAfQbpf2
SoM0qQlApanDge4kka2iQ1wiaikco9VBCd6GBI/mf1qApyTXMyLAX+a+mpsMxFefpfycBlpQbVdv
JYsgDfUYEBupKKRfoyvjejzavJqYm8xKCWDgxRvQ6guuH+1q3rFu6fWLlEwXfhwGa652U4lC5isO
XWpbFh0+fPa/uKZn9J178Rt04H1F73ww7Ee0CuQrb1TLbMYvAz9VuiuFHCx6nLzsVe14OofAsiJo
NG8Cjov89Tks/N+4F6B2zsBtkfdFc//5JulcOeL0OypcgA9mnfmwIG35VmcOPqwPnl59jBjSggHJ
+MxfIHW68h9WrBmne9CPX6OP/zvzSjj8Np5CPshyfXwz8dykO1kM7ZGNZz2fZZqsEkZt/VmlMqAg
2WEcGib7lh4tsbkmhg116orDYBOy3XHWiQxCIJevtHcKHjsaxVdiXQdrbnt4iwkMPm3+hl8pKXf8
qB5PAqgxUdKL6ASDxPQqb8a7PTxnrens7Z5BqRS6mcYTM7AaHHEf2a2cRGXjrNGDZXkJg/aE4mnh
JJo6J0de7PWoA6xM8q5IKaJCR6MHyi4oZVWfnlz23dlPsxUtrhEe2ZzCkZyUFrV/0iZ94hjtcy4U
7xuDKO0iX39o3GZczv/ne6PQEAYZatdVSARbhjpDGf6PKlF9HH3uiYQYP7ZRN7wmOAy9JndLKGjK
PeA2VfTpek5T0fT9d18VA4LjGzpTxQVQ5yRIj8QUj/DgY7dYBiepec1x5M1xlHmlY7vqM15FqUN3
5IQN+CW4k8o1ZObb61qILK66tih0biNwVVsv4ZUQEcSmCI4xjO1Af2uX19E6pFLA7hdsxyGh5lZS
UBRSvgcCJOLD8EeqliQs5haMe0Q6NaN1sVzS1QkoaO9XuXOo9vUbpQv+rm0Q/5Pq4TvajvNvRLD9
Sz+WeWIQq0lBjWgrBlLsTfbKyYKnB25f2aLSS22HmuGyuPViiOpe2cH0gFkXFvWKIu0ioy2YcQja
IGsiC/OjbNCCYVqtWDUJNtJxTbMbL6AwnfGup1pQ/1sErIqmDF3b5346ySqp3sJOGC6kQaV3x+sF
6VSkxVhKd3EOp0RC93gICpXSElkcBRWX6TlBWWopSze+HYpIZ1DsR2HWBOi+9A+c75UatG7Xaw0D
bOMLFT2wWt7BaZR9QA15VKqZ3QNjX8a+9XIKgFFy7ZDACfjTTuGBiKdL2gkcYKjjKQbMQaoIJNNl
xeJ1pwOcJCGXXBjHU7lzfX94/fVRLVQjyA9cr4aCa7+sEMUerPiunTMRGwjMyJ5gpydWodbs6PSZ
lcQXlu88m0EbOB4rhyNGnvjbTes2fzir2CaiQl1O49k/k/y7iONLwV8o7VzlqxyndgGNzdmvb774
gh4ikYS6r9QAZ65Q0prvpOpOJXXqBzX1xMFMGkBM2cvMPXcgsSBLqHEgTv1gORfUAomZUsIAY5uU
ZUiVb9B0ur8b/9ed4Zq61eC+eP2sXtGZb3LTUKatf2wQfqxFmxlMR+ivaYM7ekyxE6XPuetdxEDJ
sdeUah7ki6oDgdakohQSx2V7X4aWEIkGoiUQtpaDatEaI/6Evc3XGhv70pC9YhGehpn7Ts8AayI9
lHFLZTtpKnv8LqLY/A0ame7dPyBWXXwPpATsCiTTR0yyhr7dPwHr7t+x8eeu+U2UHL4hBBNcVNJy
F3n9w7uZqvGr/t/zTMmcOn9f7Miy2Y/3txiWr9lK6CGkjV3RmHCVBYDB+4QsopL13nirXNUUa7YY
wZ+3CcCeEEU1T1+p6GJVtPBaqTAe9U6u7k0xVEOKBm9pZhKYPjRxvpGsWYJT3V/+VkThBpdsYLaI
mahI3KDTffTvVB76moNMtXr5F/MGh2a11EuNaRDseDUplZKstiVzsfqzfMuJQvwgswT0iVmfMz10
PIa1mC13hNPAFs8FtOYoe987LgKOlR0ME2tgwm0wuy7XoQzcUmHxjxr8qrFuoH4ppY2jUtanR4kl
pb8CG4p6anuP2RIR4eDIR0CA240sfI9rsSFj6ZenyV9/nbXtRdFnD695nIkdd0Z/QWF842NqiQzf
aO8ZJfL3Ho2Qlf+cgyHlYSXsBgyNTmQIfxBICiPcJ5iRXtEhl87ZPBaLokuTH8RxO2R9kXeNEvLY
QmdaV3nTkLg3F9LNQ3xx/jBBQyKY00dBKipasbpm3qpb+fxFzdMZayWCb1VZKnjdZSnHda/7FjYL
zSK31fTxh6BqfgNbgqsOYhHHBMKVu+sBorEPVnQ3pzIAM6Uyvm/t7KsLUwJFTpp+5sUmiV4D38ow
ia7sYDmX47/W1FikHufAsYg93Pb3G0CkUJ5McDtn7sugvaiip+p/OlSo5InoCZl5oH1nWJvXe1GL
qxXhFg4stNRE9lUYUtyKQpw9Slchtn1D9XoTEbIe5thKJqvwDzNdjG5ahm04R9r2tOGQeyZjV6O0
1jL7rNZCgfBYgYSksUHrANgUVVZaOvWo0lA/t57/zFAIAQwuj22hPW0v4l6ZkA3M+fHI7KDvxUVM
wPegSHhk4ueZE0rzItGLgqyZGCQR88I07SN9p0EKhnLXvGPSYfxE6gkWmLmlIrWvx3lXKfy+Erpr
zCk/xtFhfwwcrXYDByd+kL1dd1dCxp9YzbTLCrhlsBGPOJF0H5pZvRDxCT6IjvRGu99PDu7vnIrq
vvyt8DniaFzEb3UmRotvp9rE8JZonQcq5hx0sq6xFXlSo1S3EaVpbvcdgkiqYAjYlecjzaKrSwtp
QF9gouMjOLC6Y7oPy0HguFUSHUj+hXKOJL0VpDwQsMdyWSd1vAFZHwEyYK7TKSIm+CXz/vnWA+uJ
7bj07PVGKnX4ypECEu+Rjcsulqk5IQsHoyBG/rlIcZxdX4Go8FFxFqH7B6DaayI8G1UTa8Cs1U66
4b+Qc+OvXEqOb0LNmAEGGG0TS6AKcCKlK7CxyyZHCkkDw6R0PaPrWjIM+GwLFZBf3jtzMA1N0dwk
GGZGd91yVvDptubk2kfMvYnBq4Yu/i8NJv3AvBQKQcmqMBW6hsSMDb9jnRijulRiPCXUMwjeYlnq
gVgHoHpyTbBzVthtEd2MmGsr8iVGcaAbIqaCiNhp/jGe83ikwAvrQHFNXdOSfsh9j0+akFDHZzQK
WtQdR0CPdk3E9Xg+r+7MCzBnAT/rkZ7vMHD0nkmSbMRcjgQSLwMS/q0MO44O49e4JfITETr2rAZm
JhdzmH1VVhzN3tGdXzFAa8oi+MJG0Sm1MtmxB1zMyrFq03dXx3h6Il9qazBlFpMPQPcxuBYhDa4y
3MCAnYcgPwxZ2y45eznSVk89RAKHHAKy4i4hCBqZW28hXOYya1RvjE4GICAhe1e3cQXRSGKQn19c
aCmwhDfsIxvbHyYvXkqrwlVETqsg7ZRnD7lrWOamjDKwyyb/0G3PQwgsrPDPcxc85cb7heUm1g+M
e9Msij4s8upzeC1IcPQUMvwDpEo5qeXezMZS2kE7B0D0rT3Sm3MhWk3MltEPY4Q+u4yxPjIkR1i+
YtcKwTw288qngkZYiI0jOIZBD89LMmVjlgo50GX8meWf+RS5xjHZsJG1hz05IAwvcPqPjo54CU9E
iLSr6DnXqH1kTwK/WGn/DRzgpM+3J9Bq4TtX6xKtw8RBvP6dwXq4pZW7vWjOb995BvOcQU81ydAM
t8747PSSudnbM6L+EN33TMxP7ZutrpBJ9+us/B6f/gwPWRMqHiZ9rD5aW2hZidWypBhicSgOgKiL
6vlplwcHI57GTJbMJkHkNpb1nacLQ58Q7EglUBxKJdT0o6Fxd7nPxLkaFznYRLA733u7Du3AcT4m
ZYfPci2z4SZtZ0pDbksXVI+W0yKlnQLHCLdzj4QVhPDGtP00Ef+DnecgbriUYKCVyT+1XpnHcAAe
CUC2K0pffVX8KOSFwlGISjK6JwUGVuv+Rnjg1SOsTV1lUeF+m9032vG4OfzXFDgZPA8yodUs22TA
+Y1N7zSEjY3Wx2cOinyuvuJQ/6ZxxoguIatGOBkymLBcBqr/ns9UrFtjMmoMb6vW2cc0MEZNucgQ
Ui6xuueiu4HmwSYOG/dtfcJ+CSMJ4ILLNYeViXrFzstPCUeVVR0nUs5G7zWfYKl2Bk32S43Ppvru
z19ubRZ/2VjWlOF2QYEEYePD1slLPrZYi1jDcKmi/5vafJTg5Ur8mL8m+/1OEJiILE1Dg8XIha4+
EJLOVig3DLKqYOw65FeEHmEA6THNzGBUxdypofs9FLRZ2ceylNp5xanKsjOPdcWUVrVH61sbg5x+
hI36x4vTKo1S1BstLQtgOhYCjZFAL/twIXtEdy1uhItJ6hmxhsa8vz31GddFSb+s45jl4PT52OtR
cheKWyW9Y9JSu8wN/Wq3ZGaeV+fWmNjSe7aepcPUVV/RtwtDHbFzk/qP1DhjXL3AOJhmVVAomOBU
4uWUTw8PNpW7PjgNKSqXMG9924GL0Np8V1nW0GZz9Uz1dVIsbeo6jFQmAIcE2yRf3rA6HgryPyFX
eapcHehA2F+Ta2gEN5CYk0U2TdQcbvL1ILY5bYWhnvLimWlNqGmuxaErjSHnbphlKyZhV3KfJRBq
4P9HFYWulmmjH8RHQrbt4rJRk/P7rfW6BYdL3vSgI1keyr8XOW7FwAlhPVaDJFxWmY7eeoRxdoeA
3tluym4yHU9ny/qCs/uFyDg66nEaFwNcomoT6rzL1AerO71SDd+zkMzjrCgxzUrm3Ns9ssGuGLbu
3AKBXn8/vMmXjkVbYFk9OC7IUkipYKQo1GSucTCTCrJxPv3LpFTXAVyh71k11ZbiPqjv/pCZd//L
9kEoZBTX1E9gKH3Oqv67yjjLQMSlCLULOaRo6vZf5U5LKT2u+theoMddM/L7AtAM0iOMzUdrpqod
/iEACodlgW4bhgsSx3RzEevuNQLkicEmghQVkXCJqYYeLG89yj5YbIvsA9ph6QPpiHXXIG3Q9sRb
iAyCuHzvlA1lkdNwPRUes1bFrS/AbOznfg4LGwq3GppfMIxFM2reM5hdAfqOKR4ioorZqDZwb8XQ
HZqPvgztrohdprlENjykKhQ9BFL50pFg/IBIkMk+mM/bBv1WSxtRSx0Q/qN4mgkSF5fRebHG58MC
l+7JStJ6r6thtlH5DXBOpDdgWMrKAiINxkQuYLKPrjY48ItO0smFJiDf1EcJcGfLuKF0ADOsrsRR
W65xQ2FpIa1Reip8fJWzI63qn3PhfuVzi/9YsBNKzTb40GvkXmvUa5Y4ZLFyDhx5YfexZXwa9R8/
2Wc0t+mAn4QHsywAB5T9TlBHiApFIE9jvMLA0W4+9es/acuqBU7VUy/iCPqej6h4eCjtrcuuhKvE
GAhrEMf4apNkiOJHW8L2MqlwdBpEswAPTcnZ6kKe4OP9DEEa7sE81Dnu9YRA3iPeKpK7FD6OY4gA
KIrpI8ki3dfSuECkd/SryBmFPE3zCCTiNviA2kOJ+retOiJxD6EhByYAV15ApgsrRS/YC+yC89It
QdS975U3mp6A2xMG6zVd8OwUWFbBg/BEYq50AZi/PbXTdDr9XcIH26ZPm3svZLF4TIGMrS2nDObA
xWdwifLLVWzybQuJWepmwVyHRPUX9mwZ6ypCDFZWLrJwV4US+N7JiW7sVQnmRQ1BPT9mAbrtFdRL
mszVLv29oGgNEU0Ow3Fuo9M+XLN7dJE4O2J3w6NDCCLAxkLIh3neE9FZUvLIERFIB7iwgsK5R5Qr
/MuOWe/es20zHDyH3XHjruKhjiH9oBSc0xwE/QSjm51WT2q9mGON8SMIjtccUpFVBxAbp+TBLHnP
YGszbTMoDtL17B60CGQRE7ORhxrAhsdVg3gU0WlnuNl+lfHsNdGSQptqFi2R9ICRKKTcTE076Vou
u3RSSXYKXnVauffFAogqBI96+pmfdx1IpgBL8lZtUtL1C1yFD707QMjdwr0v1fmwcogCGt1G0euX
KHDSOakwIQPWlaoPgXrNRX6HNMgtqmbHMOAI7/lQW7JDfcrLUn2UBnm4zw/LEbLFv/q17qPdXUyN
FVWF3yBQOTEaXZR5UqYtBhj1w2njaSaXipOjlKlWwWcvNEv6HTgpQ3ABlf9iuG1XZjgFYv4nEQZm
2FDZ1ki0kRLsyZpxBbiKZmPm+fDVG1dMKxyA7NZvyy1HPbKAaG5jO1AtMZECzSUIAT+Y3NQs8sqj
dCXhGzA9OEfZBNOq8s3VtsFoOxkCG2jPwtDdbjZKhQR7BZbkr+9/KDIieTfWq1v7S86l6xHB/6LG
AMC5CGuaiKVCpQOx58/VUBm6UOxIRQtUWVJnY3LNGW0yFutsPCaBZKhRSY1xqC5So7D334VzABQz
rQ4AinFNZ3kyVRYuVLBrXnGzwNzQAbOkvVowScSpNIR8M4mb0DvDiKX2s85uGgC6f5kRS9cFCeKN
RLPSBmg6BPEw8AHQVUIbdSWUJ9mRcXpyB+U3BXCFL56jaMc2q4P9ow8CkSvSpsJaVDqe09t0Va0L
fgrdsoTs3Pe9yDwTLPfufERy9cpprHNn1cr95fT4/yvxTVNvM5enbfS/tk/BJHmRauVplsD8HN5Y
9vU6JTweC8sgO4wO49i1Y1q2eiKWty0adwcS2Ecdd7at6Vb9E7bAWxyn2kp5PaOd2xJIn3JwC+MF
/CAuaBZesP03QnbEGcYvzPHir13hRbP4BMgQ4YZ2LoE2Al/KJgnWcAQ6zF9ByVG0SIfkIqoIANoF
pBXhIEUTVvLevigKH9eLMdXz5w3G4nCOxLYCNazoS1XD7o7JUD/GucqweuElycFUrKHaQDKQOedQ
eBkwU5JaPIe2QGrrUNEUcNej2Nzq9bNXcWazFpdpGF0RJ5eDdjMoNGC3WlMqb0RTHD3i6zcSF8ER
1aba+bwIzZMhUKTYRjWqcCQVbahhQbCr2EIzD43I60pyiWAHVNQW0hRpYfXqOU18T+h9CQ7a4w4b
issRI8QpqbJkSF8y88WeyW1WrUlm54ucE9FmfmG3b0QeztsqsEY2MqMsJ5+9SdVBSK/aHMLI9jeS
FoDixwaVRI1rwQYBZGdLw2IMmkC/pJ9zByON2AUdeXFWnwfpyKqTkVGeO8C9SxsIUxShKQ1yKwQD
+L8ACexSsMyEhEzk0CiEi9rgELpjo8TqJVzZYC6pXf5eNvMabDja2WtuAOiaj10IDL75NUeAQT7i
IiXefMU0/5j62iJUpJlosz5JziYm2UA5AYYCgw74hBWNUcjEX/xYtNDGmAZ5tPYS3vd6Xab9AH6I
ObqVc2XO4Z5E/9zqzrDwf7rU8e3ww7SMv/AusAhncKuGJUAg8p/gPJhh/eAr1eUASuu+V1P21cj5
wUBNqRXQmrnFaSxrdjrye8oMGQmHoMXai05q8ggB4JhfLAY8BrUXhSY1CADtl782DzpXfLSELB/a
Yrb8bCULAICEGOTpbHSr5R+66X9uPX7WIEqL9zJFd6a5VR23ylo+uKHdQreOkjLIPtDlExdPe5zP
ey8GCD9Ebn6XUE23rheDbj8IVUDe/3YyNJWmpPsAb427flcRzlOdpCCa4kLdZswj04LS0vAAUq2/
s0AYkdyudCPjjeCWh4Xo+bMLhUkj5mOH7UYA395CuBEZGL+zj35CfBL/bHADQYRByZ+HqEM0/sQZ
YcbwrBUPVyB/zPpigxmCLHkVt1x2mTKZS9bYlTObyq88i0dLCIS/4lch/kaMDQul8RuXpUg0HfpP
0ciX8uvCeHAbbZogqyJQnkwDj3sckPCxKngNrhGVQAwWgbjBDvWt5fxJYkWqt91Q5RQsfFUDxw2l
AcNooqpyWzf2XjgUjFPiJydmDpb/JI0H8xh/yy6rXjznINYiITTbZOs1z+gDHIxQvlwTd1FEmU0y
9keGj7AAMGIwbL5Nb9ic5wSXhC7ZkR/SUpSFPnEEoILfZB9e9Dn4HGzraut7BSlsgMjVOgbHD8SM
oIoRGCQSEP3CZodBBAgwZIxqWT3UsDPxEJsBRdZavTv7/GUKBCsI5/w3QPefWOvjUAoBoX7IWSem
ZrQh30ISb+UdVUTpNMk7Qt2257IKxHr4eWASbyLQAxLWE7sdq96UaqYCXjZreAuam15ttLGLnH20
q/QNSWb09J8WXJi597d62xwTHTvagXsHe48KEaB/kQQtHhz16euIyw8YtlPb65YkFF9PuWzLxfQ0
TI6WWzg0sDcArGY2uKyTUHt3KA1lJStnPBuCh1upFMy726lDNN26km58pNhEeneHTdf9EguUIaC4
fwoRMsvCjMM+sj9VAgDOETwBoIXdptCZ0rzFYNKSr6hbSxl3j2kD/5BBDu0amhTXXgeIMjRD18wQ
jT8KGxXudkxzdggiIUkWYfygjyZd01LIacxIl/+0AHfYUTVxZF8fbGxQQf6ZgUaKCydtbzdgpUDh
k/fXujtVdTOYokW3WaTQpxKFzxMrraPZhNBxpEDfmR/jKI2F1Cr/TGWAWMpJzSg8HTLNXNYDgyXY
xpeqC9nYQvZMXYRMRF+vE+j5XVFr+56ReytLtrFz9YFG+FMopp38Ou+SMnM+cxCUSdK5gRc+i4tg
0sgtp6vmCXezpwP4esP/LtN9h22WGePrjnGJr5a/JdYH+wBdsFRbcn4uQItkf1LkNXmkYLVAbytS
TKXkriJGosU5P3nVCYBohV6IpgJMlJyYTu0kiyYZp/WJ/TQUI7Uzj0BcTzhC6hGJM5W8sxZTVQJA
NHCauDI6ypDu+pcVFQJYUO4g/kz6cOrdjXZvB4bp296tUc8uj29tnPonMBUn/p6A2mj/E5Ve0kP9
IeFnGbDGsftypfMaAOv+NgfMEpzCgjMSALCQjYg7Dmy8TsmwK/zrzAeIJc1k76tjaN2RjKYKrodq
PEMTnmxzORls2L9GJigXKj+Jv+8FLfvlnNPmiekCr+b5UquNyYzmpjPrana/Mk+nexZdoXOsBp4m
uHizeSCIneRP7oA4Sz0rEX5MSt7/ZEWNhUIpp6URe8t454IE/sqgmJ3ekQFfO7JXKwva78EI+DDw
8wzWqVCODIB8Bk349HKSW8rYoumui78pYyOxuvBHCevQ3R+K2lNwRYrtjnu4L9fMBfyYNNMGErXo
UpKfXGYUgcPcsCP1ZtPROtMuX1B/egKcVzb+hZ9s8XinNEwUwi95mUsyIOF0TURdsXzFMU5JFNEB
oSpANbG4cLTxh8cwba4As/2r5f1ywPj2//baz/NP23P/YAU3e1x5sVabt5DH67fXwLsIzJrNwt5L
eIuI182TvZxvH7dYXa6Y+m6QLCHt+Yun4EkJRrxMN5pxonkcNmaQlXKlyp0mC7rSD9Wo1MwQlMT3
Qw7a70knSp1DFFWDHUCycfimeq/N7FUi7PZkL/V8vGdd8vKciz0VuazyR/ZSEmvczz+jwqbTGHgX
MTOOoalsPvgqK6inNIxJCSumOUpkTRhUH2QoReeUBqoAovFgGgL4zL3cBS81taessy8tRE3kVxsG
bVIdciThJrie/hyOawbDKsDNYI6z32NFVnakakUId3GgORgAnsVeEIi1wYh+R7/RuRuJmt8hAZ9l
NBAk34R1K3P6UlXWxurpJGkeiTKUFgCzLQILsVLn2dEcf9K9je06fHEOFW5TbcF6TmtHvIh7CZeE
+NQ8mCr9ZYIShb2q12lwLxcXOMO30X0QdAQY/g4C1qHXAv3M0dNEYhLqBr6lVmATiHazoMM3dvg/
bxLHNUHbNKIilQ+4xhmroE0YidhS8gaLm3dR0yoJ9k2y2kogx6gFIy+x6q13jr2UO/qfxhOmAn2Q
AuTDUTMBHwFv/d+U3ddsA0t+5r/B0UoYLa0+RTIOoeX6l6NO1RZrTtQzYZVw50Ajow1MpwfIR1wE
41XRgf/5feIwJdUAC1vWVw65lYOqvFdgVzL2L6VnmBzz/+KSvxnNc+3rrssU9i9M9wuCMOAJK/6g
HvoouhZd2Am3Oy3jyjKuXW3HMPfISQF7xeOEpFxuEKBpHmq9Gul+4FLp717GkZ/NYiT17js1MgZg
vf4IWpAk7LulGaWIY0oaZwWpmzQfG23UsDsHMM0B13p8oCWOW8P51cGW9FnDEHeFVJTbEDx+3vVV
ZLSIczBGiHP2O4RM0RO7Y6DsySEWoUd+VP1UC0ocg0nbTkJ+1iYNhdBn+tk0+3Wjh01kZAZZqeK1
SEv2S8i9yw0mk8pXTjWTTdp3lVor3v3WNokPR6TeSWlVRjJYF8QAsPI6iIY5The4rTQfs0hTyZVn
TRYaLdyLQ0L0jFMZVnJRYm7GdYzZIlIkaIgUIC8Jp+RZ0T3PCTrG61WsYcYeEZcE/bmjB/MPEJ/i
s+EBvImcX5ASjzj7I9eM7gs0CD5zvulKVL4N5t6SmZY8/AKLTVtigRj6591K990h5dZ54G4r8FQI
D6tYMocbrtMuAaOLSO+5eKz2SZuDB5VbtCr9KfHaFUe8ydYhj9YmMtjSayEX5/p9kH03xRGeMfLW
+5v+xONJULpcbNCwZpGj6OJElU0vgRjAeP4We2TY+1aPVGze31paSJLSp6KF6ttZOmvW/s+OopOj
dt5+7N4vZ54dAGx+HagCanZxfnhXmxDSAjM4l+oOGbGpVrBstqPwqnUoxPTN2561+iirYrDjaNpC
mvCfWZtuucRk2PNxxBNzuvsV/tn7APWTRvhZ4x/QH1PEi/5hVjprs7v2VSfBw5/7w3Cv0/sXl696
Cgbcc1DzHkNdbePj6HeUYAA8RWl9qJfhnWdWF61pv3bHsULenk9t0iFA5JHLaOaYcwtXSweljqGT
y4tpxR+8js35TmUOxEWtxPZassQKp84gfJcVTKdS6mQsoca/RXvyCpJkkpmUvBYFBRf7UP174LnP
xs1dE6rsQCIDxtGfxdn4arb0zBFhAC/8C6NiM5uq+oBk9vWZrhod1bII5mCg5Eb/5DaL4wcT7/2u
8OmDaQ3v5HpZlOwsve1+MPWqK5fDTjtVzUGIbuKVFww16o3eiElz0nFvHOce+Xekl/Fv8plJltt2
3HJvbotHaqEXqo6syFach2faMN5oN/alA0vkdCWbV3EvDMDlUUwZxL3BmpEW4o5GVLeyYqoU5Po/
E6IS8MxjEwWDK0WRvZrVp4CUuWH5p4F3mBp0iVM22EQXGN4cUSR4rjNM+Bo5pQshuoZbNH+teUoE
9RsJOyo3AwQd/ua6dd+EXc0TA2PEyXTt0S7P4r3AzHe+R7C0XKEVyb/L01wVWyz3Wt2l7N9w734Y
AAiSHnaPLHq59syaUuzLt5iJNySO4C87CyuIVtAFqnkiAOdfgcvzyELYfl83gzF76elkD6LWaIR1
xZovvObV+/v61EQ7inQJq0TEcICIIQB+I/t0QoaOdPwhHc7LrQ2YTZKtnvZyhjhjBWxqXXGj3lnV
ZnEGj3TVwy3H2Tk/xcqjhWRnpiWc9+DIdK1/l2dkXZ1vYTd3r60wEVUZXbddQL1PC9IwHmECBB6f
bms/tIKd86coSsFKoFh2DOoun5zYsgMUMw8mczcEeldioXF7PdZB6BR4mzskrxfqGjXdSnuvg2io
QxSBS+IMk+tR4UY1Tp/G7zHtUlu07UQuQ2JNbY8QTsUnAlm60TI1/VOnaeFqD7ipkbmtPsKWOmtF
ljS3CcQYzzkj7qIVJ0O5kjGWv85aUABG0IMxl5Pg9nhsc0slLIUHakt0xb4VN1rJK9Z0D4FfDZy3
IT91fmZnCUnKW1N9dpqFK2h2kOA0cQ63guIh5NjoqMq4aT9/UKRC4VVRIawjfTxEam1fuVwZLdLR
KF7STCTUHVJ0wk4fSkwvlWMaKZ9DjJI2OGA9RZsuTD5vbhccMi87SGatMWGbC4nnVfz5cf+DP3C/
ubfq7szc3QCmZVjx4fjfOoTRI3N7GfBcHzW/rPnEhrUIDFfrM/UuQO5OJhKPtr0DheFLmjb48uVP
MeCcK/n3DeApHoihB9yW8J70xcN1OEDSHGDWL8Qc6qDntiG22UDdy9MaDmHk5IzcDvv7kn+/LAqp
wKSHatDtNfexrWgdjmz/Y9qWzqbGVEZpbLt81Jl4wlR3kOyl2VDQrHX6S6pSaP1LhWexTMxsgB9i
2yERr35p4lMoD3Y//HVzA7jhDRZoH7wTneVoZODyiyLEJjWWQGfgd0Pejy8krWr5BBFh1+DbCog8
RG81kXiDTTHj/dtXJcni+XRLcOAxW2v9U6qv+hnJc5uxeJKeknPgwKRUPxK5WGRFvIFh5Fnf5KE5
+6YCZZBNzRC3bWM6GDML4xh1oAFhdmXUb5oEW19Rf/wmMkjwYkMtxDFHfo3u7hOSwx4RcWKkMyCo
aTlV6RBsnre9dB1yFW6YgP0GIG/mk2ukYXI/j/iz0Wo1AtIxD02XqVRVlSm7uhkqiSadXN195FrF
K4JrSD3scbeISCyqyummA/tjtm81CVYs5w13uamhCAgMgV2pIG6PeYLZlKJNBVyivuvsvTmar+zd
ZgKd9Q8+FamciNHce2E4Ry9JXt5Cj6xzbVXjnZlZWuxDmkO3y+YPYwUXJ5UQXWGmXiIrw7+1LXWP
vyOY1cxNPxbIR570UR6WY7aSUNJARqOqjfTGoWR8pgJMshkIKMBILV5LbgLMRopT/LNfYbJLlerB
HEDIssfAFSITJjaVp3MxMkk5C0aRugvddaWf9nuzBH4REt9v2bZKZrXAGoTBkfdmVtfY0Kep0PhO
GIjud0GON+vU0RmFOkuVX2FXaNiwJn+DXoETWEoJXGfWqayP1BpZP1ZDh4+bLJb8Tv5yd/sPw+GG
8gflyT06SGs/rYGiLrO8eN96GYM+lsHTgsNzZ3IQjTkiME9JeIO9wcuf3Op+K2uwoSDIf7jnkSs1
KTUyLwFPQR/paANCg/ro5+ikobs/Ew7eSQxAFxkcvFF/XSB52oSIAgEt4dvCasJBgWP+CxQIQ9VD
IoTtTQFaupUZLml+DuqOZxwkx0EiLPSZM0Cbgz7TYYgHQ3nrCpAxF1TnpmXKwX4pAW2FdBTjfMgt
/NgnZbyYJIzFRyJwvIrQRUJPYl+cV8owKImw4kNe0tqEpxLVN8yO69kqIfftkC4a7vrx+0YManZW
MT+d4lk/Np0T7NaNLo3KE1gxdU98HQcZHvTiyZoKJJSVSabMLYo/fwti647NZnABQFdofONnLTFc
qczP2GXdsr2j9RkJJipTB5fbd5JVDX4uP+Bim2FpA1CU29g6DzmVbC8dGiz8w54D4sI9gQBWktL0
vtQw4OTccT+dSZFXgBoKIhOZHD2P+xQeSdj3b15iASGRR9jbWDtbIeXyStbpHbZx3aXgWOITrINm
S39bigynDWS1IT/MZKMMTwNFRrphVA3bou8sD3FAbvWaa2LaHNSTsq6IseXus06v/C2eJf8nY05W
d0pIoTXiV5+ynHETB6Q47OLVUrJWs3ltqDnD+4fNbHU5hEWRln0Wn5abvBMJE6+ZdhrCoFUbyQ8O
6TmQF/BPFqmapMDy34p8wEiOdpJelD/Bxo20OTaY/JA69wAhg3HZ3EdBdmqMZXj9IxmJxHv4uSom
H+RM1Z4soFZwOMf2yhPwMcVJxI7mLz1K+fXljg1rByvMac4GQQKRd/V4VEkSRlG/a2ZpK13/C5ow
1PzkEEHRnE55UEjt+GJJuWiM/w0lenmjttjvm4w/dkurvOL2Tw7cff2B1a/7qDgOkM4w0KPLpRbs
bK1DKZdAzhBMq3Mh7qTYcSN4H0TsKKApjg7RCdS2x4xOtVjwyPx2S7v9I8bWQP1xLQl37hFFk2vK
VOyz/5q32tPcS+bSv1E/bkQDbPSj8fZ5TivVVrnPQ9Nh+Qa75u8y659reKyTpQMLC2RCRIxnsW6T
oZMCDOy6c8/1NOacLRMOGewmr20qmpqDfeoT+KdkL9owdRfMOcdaCrTtkaUObY+Z3E63Ylm2X+Pg
ZQCWFvwHnDh0IsyYkaohlrkYXWZw6ZDjTJ686UvJl0nQPaCMurwsAHgufwrDC3RaQmdOycSfKeGy
ojK0+FDAcCAOiH98C/1Rs8xXnwQZ6lnULUZUq77HQHp/JFpuxBoeHev0YSZwJyV+ILbL7wYq19FW
XXa8sCr65NxFTFG1PDqcyhhSNwnIW0tWGgeZPpHYkCN1U+vlM6Y2C3gCCrT5vSLazbl7/ZLa1QR/
XVy683aiWBBCaqfhBCNwUSGnN20Vua0LKzHA7I3YzJjmneOVCaU+rVA8V8U11CISs05JnLieON3S
SeVEy1eEKj6HxTwH4MPXnWu84vUEjVR5K5yLCrwRYls21vheoIvgbN6vgg4DCEs6ZO03y5E1i//c
Xu0vM46VtoaLrwZQMz65TLUmSb9SRy7mmzHs7wiDDu6/mXZpZGujKZFCO9YhfUDGnISWyWPV+IMY
RgYyXho3r6J8b6wDcybWwcG1gPuD+Qa/talMEvco5oQON2JvCbViHl4CcEhUBUP+QPT/225qLtkZ
rS2b+I6BahGTCpz/jqucefeZN3fQxrLcEVyJOOJEqnRWNPoHr1/8qb4mzjGnmMcyML0/wiPSXH6G
YTHyJgTfVaq+k68FzDFXp6blzB5wd5xVdd3yv3ixiVqoiY+aNIAnDkO/6GbWBAh3rXYXFgGWYaJB
bGAkQROvdFlVqp1jQAdknNq+8l3JK7hhAzEhRwE9xr0zXEkd7HaprruNs6htFUuAWiOUWCXzgBTf
4m/cjrX3sn0Ow5rODC1gViqaWvSCbaff1JjptaloGpiyiP0J0ZJb8PSafm5oVDstRnoHUQuQAdgu
q3M1kQD4U4NSz2iA6Dz8WRZyfYaB1X4nBRteY2lkJW7Saw92j7rSesGRikp6kEhiLOpb0o5ZBPX3
ZvaphNZCUyLpzGrmxERAVxEJqrk8RAQ3u1YUr311Cme1J47bJIKSEFBsTs86ddAIr5/aJLCg9SlW
KAbnjKBmEkTqr61N3f1+iMQOPB0yhXrigxTO330F4RZUxRiS4wPAwQgQvSp3RmTN+FiXUtoaRlB6
olEEMIJmuSm6JL4PNmXDkL3xDBtI2WrQ64rJ4cX5hIFcsMjc6KF4fY+CQzqhHunqYXUjWRqz3um/
oGobW7Nh++A+yQmKC4FpzdjfrZ/Jx9XFacte3dnUwG5Gm5EjJSCOizCxLz54o6DgpoCUln7ouBHq
NLo/ReH39IWAHL2JNEN0pME85KP0ShGOiyCTXavtp7ahF0PmsMriuB6r1BTSPpvxpJU4r2+OgHkQ
17uQIhwM6mCXV3V9kXS+hiX5ezh/n2QGqxQdfBfBqZvF02AuLepKFPjECmmc6qRX5969uhw3dh0c
EWkrjmTYAncv4BRzvQb/+x9HsisB1TNOdtUI4a5EqkRUr25IcI0j+jjzvj5F3QtTYeq6UiPQzXg3
62qCLsG7un7PIqWXAjDj9m839MeaxC83yFWu3OhzL+4NdkllrFUeFGyKfvtUfR3b5e7Ne+NU3sKa
3q88V6YU0vMHSfU2nu/2G5+J/NqXCga0u7HlFbrRcmfuNWbjXx5jh885tNSmk+Quv9Er+cAfpiWi
r/qkMEf5jmUmYbImGeC8oLkR+IX1w7p6xwkJ0Q8AC6tYorG6zKfg8cuzBJxj4JrusQgYxjiXQzjV
YBwFN6IofzPSo4EQAf2GNyESnGdEnozMXLvcgvkHtG5ypU7ez0qiibLf6anDzcUJDsrTLojCYl0f
rFaEgHYCF8namB4JrlkjR5OlOZ/YX55trPROsEDCbuA+lkuKYnCO0KJNoDrF27ytaZ4ksuQ6ATCQ
G1TM0un6XBRM2LrhCEEbFmtvWX9BV9nFKkeUdUu9xUlKSjejlBsWS59wczSvhlgeaHciuI/SJOfn
GybDEn8PReBNXZjwtzXJhwcZ9Nzs/BbVRHapc1oqqz3L9jq/Kvqk4MWgIgkIeheISb4g92cbzMgS
aGoR8+evqVGSumE3TgPrBdhVplxhHc4gp8hokSeur1YV0DSmR1+gFNfYX5e5LjRlze73EpN2xVpa
pfrJI4wdt8q30rp5GB8wOsYAwi8mrwby/zWrLaLVUXZtyC1TbYKqeDUygYJQOPImZO0LgcT/Fsid
oQbGRLBI9veYOcU9K2oOtcWrEpRlxmGqqCgPUstyFgc1X+ub3To/x/89eyJOw+rB5RytGaOJlhfw
6eoX37+XcjZZF/j19SbRneQpv/3ByRbGwZ7yN9HFDN6KOOAFvjn2FvvHF+vtK4at5LolKVtTzLtL
ykLeIXzdFfDWmA7/u+qXC3/T5HF2T1dOGCIfu5/TRxx5ZiRPe8OHfTZy9rIPYfzVinblTdKOboXi
PUhWSM1yMIysBo4P9YByGB4he2N7bpjO+MBxhEz1oGV9xFhTaIg2qFrOgWRZBO8dqEm+bcxJ2DGD
wuB5nHbd+vqazkdHLTnLIPVAPiNBJxlLFcqu3xkf2XU4F35dGt9fjzKysOVgN4laT4OA1SStsoZB
6sv0+/bbOC/4B3hYC9hk5P4ZrQjtR2pS4kRLAKdRcSDGhkQwixLFk5QsL9SmBmjj6IbTlmUhTbz9
A96JIsCODf3NEGvBkZKdpsBfPLoWAVvt/quhade7w5FoWvNrAtxvc37lNW3ZE0j2yPbuYKWkUp4P
OIAJunL4kMKag61HySofZpns4OOsywvKy4cpMYJPQ7wAZqM+bUk8RGvzxaAz4jqJOMg46nxTMYCX
Ak3z760DzvnW/cy/x0eIHDvRDZ029kmb11KeegpsK+gO8IlR3i58cjiMCTHgBfhofhXJPTfXhm4w
Cz+j8YjVD47W/fW+yEI8aPsq1LMHS2WEZYTCqDEA4LUqiE+XqwK2o+d82m/2ATzmFxSsPHYTSCwW
LQXTNa0R1cbyyMWgkqg9+oDJFQqfotJRkHggM8Z7m0XIkBwABw1B5j/v6s+/YhwpWHjuog1kVmFs
AoQXmvMIkEf/6oGoP/vp/5x5QLY0CvyB4cfvvfiTxdutxDPbcyV+vmpzydLsQ5Xw9fmparCoeKuU
8mzCIQdMR71W3FRfi7HHzLUUcORD4yNvAvp5CNuagAyo0ikBCd+oOlUaf2LtGJ+Nt82quPcAVe/h
YplyKpUTaXR6xhPdh4uLmAGZ7M3j3RD0n13c77Xno81+Ltd4n1Uxe5T0W1EErkth+uUvj4OLq5pq
774Dg0nbVELrhGpS1pAMpafKRtkDec04VqyWxg9OigevJvJ1P1fyJAEwgyJ7ojMJA6qthXCN7DFr
C+yQmY00aejZEiHI3XNBwdny4US7nrrf3u6flhyG329++D3dXaU1qCPhkO3JnatH7K2KNv2onKcj
oTNpzrcAng5q3kNZiXAHX9DdEKEcV7IXqEyxNLGViW2k1wNvb6VhJgvSmSKur4hcJg3HWvM+hDuJ
kno8VhGmQYlUZgZUpQ/nfSig+f6kd8k/zlCRQwjOSgEXP5GDIDoMi59rLIEDt3YNp3SuS0ypoQ0j
XFhYU5khU5Sa9S9loJq9rvLHX1x4LVOn8QOxvfcqqDLT87VSkxa3SO+br2nnsvHKTYMFXyQz0Av3
JRhoEv+h4GKOPAHtZo+DYa9ufxhX/Gm5fgkwE4mOFBHvOOfhwxWAWq3oopnYdEXU5f+Thq8Jw1Rl
/UtR0ovxTBEEb7qWoG6+e4YRM8L4fhx5/lCIkRxdci/ge6Edx3MiFJMwO+qcb/lStuxatv15QDhw
i3PTrOUkYeas0dW/VvitTF3gPp3dIyEH+hLdhW+KWbxdf38yD/GyFticgtKx/GRz7b+7QYUpeK4b
ctK8UD191lHcZ4CNQbmM3KCHXoQ5EKRZATvlueNbzHZZy6eL1T0+BmKGf0r72ys9+L4MTHbG1n6i
cqn2nyaWh3jgnG7tu4jNV9CTnW7PzrXzxgmmE5yIBuM9fHY0pedZq6vQvEPwUWuFgsbSbwluKkKS
YUeFXd13wPGzMuOhST+plTPzmhx/zIp7G/SL8wT01yvbT/UwENP0+wkhb/ajeufmYuBhPSBhq4J1
azuBoY2viASPs8fWDmUVdjEWi7hyGL3LIp8sRJ71aNoHsnrbpPZgciRkp8GF36D718yD8oGuEhIo
8pyGsnD1buXwq6ImIk0JH9Ane+hASJkHZE4nM/mq1q2VTVy/GbQYmH8gysjXWWLFubTQ/kYnYFVe
peM1jcw7NaraA7gRnRT3s+E+l6NeYFUa3fBxoofGV9PiL3hP697BisGROxtbGwvOp7YjixKBbRP9
uSkrxAaCcMjrBFnUI+B2EKhf1QhjvUZ2yA7Fbvbo1BzcV8fqYgPkigooq5Ekkbm0jCBG7EhTdbnp
7ZnlekfJM8vw6QL/eOXWEDOgbnkdfnBVJo87o7tWwZBsZTeRdrXF95Z+ZTqlNGzdTvjshlTGpB3y
xRs6Xb8drp0tFtmJX6PAzLub2612a1liyw7TJ4Jk9W1ntB1WZO7AzMwu36toThdiW+HABrns0OO8
U0H7XwQzVZFZ1bo2fgcr8PIOMJXc1OvSjKpE3auN6LYpOl52dG8dDVMXpDhd/PttRnwl8UTEB4uy
kV+eqeIqa1pKx6QeM7c/PGawzfb3qo2uZcGvMuLY2lyT1r5GDDw0vdPv5p1CcaAorG747+Rrhuri
YzjAUiYrkOT0Y4sg6ezPJqATr8pu3rMNTnm07aiQuJ51w2yiYQuHeYDngr6PqBpzanetfGU3CJ/8
Cjc1kxj5/d8SrUOBD8RhhX34cK/nsZn15HYC3oWRnOkQ39wwP7pMR3zYzLcyN9pQeMXHmYo/JOQH
vSXCjOs9cSNYahGclZPE9u/kYpdROHaWOgRb+GMim0fQgyqw07MFa5nHn525VZVYU95S2tkaGHqS
cTd/a90Oh59sqINV61UnKsiKShBjL/XWk8ubBd/Lkl3PF78VYVIJ3Bs3tbC5SKUBO1lWUstyt9Oq
tJe05i+pE+Fle68gOsl41hsNIlE3+hGr0UlR5tqv+yREanjW/U6TSfXfq4PPnR1zXtmKlwyHLZx3
TP+AWEQUWynO+P1161+U/32W6E4Y59LTwCCkyinfrI5fmIv72KRF0BEqKBsEFxb8LeeQv0q0zt2i
vxiw14PJBQEpjX4b6MSBKBVX70ET9qm/OONkzaHJJqKmbbN3t4TgWnYHmMKGnCf0faXnmE80btlC
2CJ243iZSQQ1nkfVaNfK8hf/EFwOyvZtN4Z5/2jQeFv8AlYcuykSKAN8Ct7BzOKjEnefNicFxLxp
goVVCv+8k+1/UysgnwYHlBSzwdO8dFizFIohzxVdwReJL33SpvXgLYMTur/hs70ckZP4E1oYUzru
qC78vkDOz/riUNBz+7tk4taT/lxReUy9v0f1bNKjn8SiuEl6QJ01g/9xRFZjThHexCH0aaL02Vzm
/LRqXpi50LMm9doUM0ETvW/SXjABerYktH2QO8NFeeN0ih2eORZC4ewn27FWr33f6eIdBfESagpW
Whv1VTN1OoubCaZrmmVyAu5rnpXX+4oIkDr+uXpcqmYmhJu5UouPGtKVYFmtnQMgQ33aWQtIw1g/
NfX4zuIngVje1ACbkgaSuSR0hL1TFyH36o0Riq8QobR0VOY59KSieddKUYjAac/QNrEy22ckCvYH
lqa2zfiSK1ExbbWaVidKgqBajq4LTh/lpZsnqJOwYw74jweaJZ9jp/RP9lIgrUZsmvVl8fnpeT01
Ma+uyKrMVRDPKGIkGXSXwzWacQozrqorKcvsXfWCvVD3ZpWJxglNh31VQWibGzMbZnrLVgXyTdfo
6YGFgc5HFWkYDfJbu4lxDnWu3FWv3Y/cb8CH3PNZgXKZGElVcBSN+4Lz0231QqCVwQW75IRUT+jy
2w0tVlOMh9kA49+jmg3najV/JnptPvd8FY2C9Dk8voqqhVwkt2erQbg24inAiZYIK8A3sPUHhK1r
9oY+ek1MtvXnxLo4L35MJ+2miqeSrBt5iXxZPSt2TPeZRwMANjy5IfbobOcAlj1l9hxTVO/zZ3Zi
62zjPWOZhZ93MxJ190MVcL0o/e+YMkYI1GqH2sGHMDoGAzKqb0la1tjQSatQI0SFup7xEBIg+gZN
4Z6Ql9v01Ck+btT1EdtAZp+ciJlr3xNU92OPzWYlxVByeyCCxQP73nL24wiv/i+00Htmi62BSyCT
2kLuskfKF3VNeLM2wyNR2FOrSz51xhrmt/t+9shKNdn2yH+cdbEN7FDv1+dVUaQ40PhKmmpeRaE4
n53243n/zbeDigVqkWl/NKKkw18Pudj9b/nAyuELrmdpqzSwiY+Q+/jsRb9WGh6l0Y3mHURbZbeg
Qxu8cCuSRj+zPJkvBnwl626ho4LNvnEcHXuYt2AdqkAqF6/c6eSL9b5IUas8EQ9JxqU7eavN9oZO
EH8EiFWS6Ir8vMReCYLvlZK9yG5R8Oo8MSoVw0t28lLjNOtnOk9NyZUL1AzTXpDTmgu3b3v6UW6c
PK941WTgc+5XePvtv4Cqqj3YY8zCx/R9YcOfv7FK2F+t5UwL5NFkV0duFwDfNE7AXFk01WGcl35x
zynOVXE3plejai80m+KPxcnmOQBTxijuzFxHrzkUj3OfDc5xrlUU/rSHoFOMIYISD4RU02iznQnY
QNN/3+mG8ubTlWg5Hc6zvovnub3bYzI8TEi/TJ1mbyAfH0oYJCRFx4SdGAEybDjfoCn0DqXzWA7E
Wf8gHCa25qv8YeEAk8dY0OcqB6Ev6UjuFR/lge5Y0OQsliQGrjB2yLugxLpuWFUDkh9AENLxF3LF
z0jiLu8iAdGB9dm2f8xLvfGFgtMQ9qR9GThJTUJWJxux8jzXfACWd9pAiduTK/aFDU2PDDvv8FPD
uwkZgZQVMnkTE9JvcuYSLANgWaMz1dLSccrNZbUhDBntxQP4MoWImbOUEAtlXCzoO6QDRLaTiulK
JLHLYvWMeVrQ7dxQnQXJQ3peDzwCWjdpWwRexoYlbTkhlt7eSWDlfwYYRa5dIqUn3syyvFEBz5vS
2RiHU9IG4lNCyQaKZqwH9BqyV2WQqBKWlZ58p9XJuYkW1cKDRLtyW54F20Hnuko2QgrJ1+jfRIY6
hS8zbvz7+TAYOUQHE/+W/2crdTCPiVGbNpZES0GaHRvm70VtFL6QzQOwVxK3XLGFvEbYG6D7lC2Z
LV2kTLwUyi9BpjanF/Cohf5bOpFW5h5gb5QKWkm903E03AeqsFOnRqWxAeq5LiYxgzL/d1RVeFKa
ECiiWdx7yBG8tN5N16mjiXKmM3/htbPfds9dSdocNPAv3ykYbRoaAbpi+NX8a9L+Nq0lQmZBBV+G
29DhegVWXmh4oANf6934+qwMke8afI/O3XkXodkR+r6k3ZrtdAMu1TZUFUrEE3QyrHeH3ZJLjfrG
pxKhTQsZclD4uOqT/tx5DxYbHj7eB0GVowM5gVd5hHIG/7SKIeTCgcrkA8IZTxZxrbd54Lh2e4eo
msYOBe2EwjkclQncO29OUPQpVUhNIyk/1Zz//vffGvZifwSpNaZuSgxShJNk8XK1p6l3qNE23ukq
3PAhAggB2r2qpCggc5716pxyNLlP+j7XTWWWO2v9RamNOJQkVm+Xz/FZ/A7+Bwjdhm31GPnH5OHP
FvelKN2q+NLlWHWLOpKwGV53wTPtYM8WsYEBcGb4+eqdYSLNBP32+eOi6JPeNdQ+aWortIAKKsOP
JRmKW2w5wf4V7V3vV1r182qmVTp+qVKNPAOJ0HavfnoWbk8MYPHbKJTw8rAP3yqX2jPtMP1X2arj
Ok4TpJJblgvqkqVVPCgWGZubRyY1lZ+3uwtqzv7gKVhe7Hm6QIeifByyMD+HnMUqw2A141vDx7+u
oYKjF4bq1xBjejEKoKcv/NfqrryijV/dmwbd3wg74LB/Xb9l019RHeghEgKe0DcCC6fW74jKhYye
bql0Rn0CSVD1AMaJ2/RCNSu8tZgZi86ETTwsix7ZXSmrmh8Khvi7YIk+UY3poxZeiY/BSk4diPFy
1M+p6DxWUmyrwzj5+mslW9JwK9Za4X8KqvyDIa7eAKi0dlj1OhxZsSZodUCV/K5ESzYD3ptytisV
mpUoaKAHTlGa5yxQlTnSvIgAz4hb/4PyM6MpI47KzbjF/HamLmdk7bWZ6VRsjAfHvktC+sOHCveN
IqjZuGZQ0bo6oPV7zy7ZuZu3QH2DLwDO0r+sqJpl0xI46+CrZwKnStG0hC6n7lCR2rYtj4OpeiAr
+fFS/bFs5TpDxsgrOGewfDs7J4UwzVqnCfGWfGOxm1i/Re0elt6GcrnQHprXJbDFZ+qnWqnow1kw
+IBKFcjUys7DnrOJYggUSjTe6oI2NQiwNKcs0JwsxDh7FT+t7T5ir7ro+00swC2eE/49uXZTkK5P
LMzBg3+4ishn6+7iYyjEd3UTclZdTKha8Fu/THzlWM1dHF8RW4PLJfUpHQ0dDOJzA2WGyBM/Uofi
m3jwE8wZOCXtCgzOht7VUIq7XIhnwu+HxzEUl9cQFI7FRK/pX29aaqMEydLIrWxl7rVFWDZkQPgJ
oPCV29jOs+ZoIUu6sl5L8VO+ApvcZOUsS41NZK+jo73TxPz7WsIEbpY78/6z1oCPQnu+MXp2Q82F
yhzzUEQaO2Nju+CU/iB64mxY0A5twj7OgwpQRq3qI3+BSayeBAnLuLiyxWohWZRBWNMQgmWdrD1n
SzPAxegpUMITKm0AJYplQ5BrN74Jgp31c21nDo5QRs8qx8ccS/xhel2LFKQy3jNLFOXgMg07Aih3
TYMrzh9pYE5d1Zvqlx0J69WBfcKE8S7lloUnIoSDh6G9Log/M103yP2Fx3P1pB83yjZDK8vsVk58
jp/oyy4RPWFpShL+9CjSF2BwrzpxUqm7Fx9/dojr7D0UGXCE9uwIIKGRAdFUrxXeYIKqLNilwtS7
t4maAGogBdlHEJP+2yyrffBGWqxd2U0MUG3CN3B8vl3NNgILaSLC6Eb9ZLvQR5gZ0AARzJKNi3er
REV1u7cNA7y152AenVQfrqg4Yi6WfgAINSFB9KOwrnim//ZfGvfV5DF2z6K8SvtyfbUXaP7q3JpL
FdMhUMx2zqFAgzhKexh20Zju2TqeE1vtNlEZsurcaVjxTlph57ggdDNB7oSkNXXuiQXf/asN46Z1
3a5QtAGEmmmZHdwToxVzaobEd3RYWRvFm1GYCgCsyug/gdxUSh2UyEhlcn0pnCBO0iPaUTuGfj1k
PkmYQmpB9cZ4/hVvX+APcHYzSa+6osLJ6OTdDfCscMl7OO2jW7M58Vbmd3Iy8fv3XlAK/5R3OOxL
qn1KoP31rW1cr++k2tIezbHgc8Xwlc23538P5cWXgKJYxbT07QROyLm277vDrLipguZtC8vWcsrh
CiZlCTRBd5Rowt95QLatDDKWgXWfAxuaHEpLg4xt5Ue/jwzZJE/PPGMUPl/GK8+6lGLx38ie7vzn
oalgpDIijgzkY11b9qmQQW0Z/Mw/KThHLKpu6terZ0D9zZ+PgOQ6GRLpnqKXhPKQu250g2avUoVm
5ijPqDi+oM/JTpY6wexus9IkakZA8ty7dQ6juU7Q8kPjUvDSQfNe9q6CDmmxb0NM4+UTYcL/O1ys
4S9pHaI7Mqd8HYg1OcyqgqIAgqaPv74bL8WJ2wcrUM4uIA93h4tsSYMKNVxW9/nUXMb8OdcXmkcX
6P6HGs6NEeJ7N4W2VUC3M6DSXEGpnDBuBIXTHcIVQ00NToso8GT/NjT1a7n/fbkAc1vdDfFnc5cT
FBAo4NrluC7RnY3MUMcDip+r/wHKh5QAZc5RreDIGe6GNNzJm+RnTgxDJnPjW7Dfbr4S6pHJykMr
mdd5MCZQqwwZppU8gPG3rpK3Rpt5ChRxkZZ3co//aP+lpimR9bByCVRk2FdgBXgyo9ViPKc6ak0o
qwtsKnXqOCiN1msg3R1YKGRoGZrlSnPiAmraHBqlxLRZTSVRaZmqTjcGtEtprRS+NCI935c+59yx
1SeObM74dLhFSjfkMNTtGHQFWC/JkFEHagwNB7qXlq3Rdl45NHMtuIn7GviA0HjE3yV4PoAMpjvh
LBD0Oboq0eTJttS4mCQtuFS2NjciG4W2uokbJV5Uj833FZl05D87DP2DyH34PG9sntG46swjchCq
ANtNZXsGJP/xdj7y3sh4Ia3ZZm4I3SMjIvD13AdYdYzE15qDABMBZIBNG9trybf9M5WCIytLGeR2
Yxh1iRQL76k65RPomZcHduL2Cp3aynAJXS1UOYxmWenbhJCGo8hao3PGGyFRP/uqun/J5muP96GK
x+mRYIClozr6dmxvVjelltXYmb+oC6gp4BuMhmOThaWaHv4FGSaLHO4Q0OelZqxVYlUjaWv0Vx8W
Ola51CGucdtpBb7ZJcnwDnXESO6iLPeaTvC7gj6YIVh0VlfoM7FkjHyQ/kNd17oL/FLUas56B+DF
Y0WuFhzwPXQVQYy4f4KTvqOKdmYQYej/qxWJLjB9C73xTnQn7fdnsInbYlUqiaYC53Hq6tdoflLZ
3mqlzr02YPDxCu9sVnaenQyyNG4/zhW9aaCJYpEYGP/hCNuzYRar8QGAbO6wDijC0mP1uHSZNVhD
ofkigM65qZuOGiQsdWcm/b+VQYRP5NY3yoYBP0NrRq6DFhXBV83vCLzungJwIXUOAf3NxC39Ne46
jtXLKOJlypkh9sZoellloz6Yf7nPURlxTtKW8HhSMWdCxWeG3rz8JNfK/jipSsyGqNV+5WJfZXAw
Pqd3d5KbCoZNEN/4C2sw0aZ4LfZGNj5DkT6zYgIM3d+iCI8M1a8+UId+tyusZmmnb5vg9Wa3nos0
N6PyUMTgCeD+uc6XZ29y5Vh5WikgZbBKPxvBfN2eCGiMxhDOEDvtRSGtXSKt0wterT9NTlyMqBXG
ITzYyR7sd34qHot1rti3NP4ntHmsTmZ8V635bKlYVLgs+rs2UDIzhxUPCx6bjLFYdrEAb3dGuJT6
2ierYato7XbHuR7fQlK4tPZpr8nfcnh4cFMy57DOYnxDMwmUjRXs64aMrcBagDlZICh4r9Zm2xFk
NqFmXo0EpxQGuL92ABX2Z4WnaOcaGywVv7xjNJ3Lv9mNLq+uU2mpuz0QQsoZhqt5Cj6IbhJ0O658
Ps7xv1b/gOQIg1vADAR8tDxWMIeO5qSgG+H82xPIhfkUJZ4xs+ljwObGMj5Jv7qHgeSkqeKTvWvL
q1VebLjZczq8H2p3IZ2BhHYSep9ITn3dAWB7fbyormG/G8mrOKQkfA6b5B2CeY38aoRLDfdcU8OR
Cr+Ogp+PHdgSIZ7NQ3TJyaiS/EP1YDy453AEmkvr/Zr0K1MKfxIccooYiGiYNhwW0hC6qRtbuejV
Xr07A9rGkGRuKLuwlNPakVPnRk4HPQHSke2AR7AwVzWIksoIDuPs//25EmSwFtq9vSUqqCwvJFsT
qucfxHBNjw8oHUow4tl8iQXgu1z1sSTld+EbyfmAX3ytEUVQwdmVSYA9FDSthSn8mnQFnWyK9r/N
LfUkc7EQEASKuuD5y4g/U9+ok1Q0x+gZvOMASi/+If3Y41BPmmFbc4BMnRA9Frdp31rB9ODYYXqb
o77CjkuxCORnwQwTtJyp5wdIPBJ63LI8e3vfbFV6wYR1Jja+p0aQN7QJOIW7dm+rjUY5krcOkJPl
vWHgK3qfVfHotpZ51SiGu2emw2WZZM6b9LN9qkpKyZUwvX1LZUkz4RTi63m5Vzh/TCyj1SVeO+O/
XiT+VIj4A4JN4LzgJLijenZQQu1nes6up81Fw0ie5cG88S393n1BoKIUSlvP/DPSPJ/jeycLnDCQ
b/yRgs7sSGOEodyKKNX19j0h3aQXO9HXNz88Tey3T7vcUk0TyCEeqH1RpjqoVVdbHYsYHo8MLKhR
4COR5l+IQomLVvYeGo/51FXvu8EBdLsaWY/Jz8FnGVAv8zsWwHYQb5kOZMkQtIp//0T96Vbkji9M
li9QW+KnWpK6CPNlBlUnRi+Uc0AALxLhIu/nH+OfC1F6ydYx8zpsCNFs+Ww9N7BwfXDuE6OrTSTd
bPaDw06Th+Vo3CvuKcImzUEmqisAKUMMq0VvEERnTRZPJ/jCquwsrexZrDJJDrMy0Pl5dw1HmHXA
Dof/AJJsBCwTGp7YL7FkCuFEh7qlDV1QczxyeWWima5bxvA7DnTPTIzbxN1lA7l8KtDP5j5UpzqT
pjnJ9DeNoAvAN/Fo+76LC790Rp9/shAObYCY/x/EmbwTGRHK+9x6NI7hfcXRJFciy8XC2F+sz+f8
iIn+QlFIPtceDyRQPL5Ou82AuC2Nwe9aVx6rD2nrb558PA8bbYX4TSodLFq9u7UxLUiq7mowfCwC
IHKU1bdLmb01lTI7E7W5WWURyraRco2S9rLhYuYqhDuevlekAybzReYojDUiBd8PDz627RjSUKHS
yIeEIY2TFhwA1fSvX3XQKtpJQ2Svv0umenZazHxQSmpITIfRKefXk/0+Xbl6ffAcDn2emxs6AsxU
Jl/0GaknmJsL/dmWJGivUNomOfJUQvFEI8InmKJaKQIXGpV+r8jL01jhFy0YqA9uSWhMrIpGQGf9
pjrD2ADXS416h8K9gozllxoIFyg6fU1Thq90+f3PEnB7M9bGOvCFbXlcfBTUT7NNoEAdE/74c3vP
DkAeESOzPpXb6k1GmL2jNssJDPLuY2+bpBdmVYt5sFV6mr0HaBDUuivITYUyWHFa/fTGnAj9npqr
XQU9geVWYnMQcJkxX0hmZZQEa+SuTiHvM8eVYUF0IBuVARxWiC4Wq7cjoHZ40keeNz0GI1+MlgNB
MEVxGtUbHckGvE0RYQH6tnogLifxwVV1T4gts8jesDk5oMnjXOHLuf/wKffX869QpFjJfbIKeGXg
hYz2aY/3y6TfypZkWo8QHxSljCQH5zZmmPlO59/PmbFwGjw6RgoZ/gf6pVfFGFdhyfZ0CmW760bG
0l8hFWWsM1BGPdZicpycHa51oVGUptc211LFz5NLyikwP7aQ7PiDKIAGAIczCJt2T4LyAsOpwC/+
8NIs6SkwrdhIi5SCefmW08h7OcoedrACSbHVk9Ig6k6vbff8NHpwUX2I+J8OVFZRT8orx08/lngl
OMWv2DCc4vCx13y2pGir3mdVzQP4IsLam011VpRdmGIgkV5Sk5E950sbjxupuX+aE2OPTQvqzIoF
pp5KcAK1xQV0ZJweGrZJkFskvcaP7yn8DdXhrKmiiqVOBdB/4ndLuqqBAjKS3XbSMTS2L7ZGoppj
BdfBA//UtBkDl9r9i74ICgssiJovhhZPsSJWn8HMtCJZ1OkG0M36WEtkYjyQqpEv41rz4aH88UGU
Y7o7OMa1ZvGkIIO++GST/3lqwRSIqyK7gFURZ3TiETP/kUS4YtIhjomZaEHk1Mr/6o+kY/0JE+N+
EfHYqA5kqDW9hBYbgDNslG4jmOBM8DnKgr4pbxEN0m8Y2RlZbSq7UtNXYjZIFBydRDcOk3yzjHpM
blm0Ad59jBLmNyVS+7dcj79EAXURKEG00z1ICbruD9J3XkhJ2iP/cuyjBlkVJFn9T8leAgubjlIQ
srW3+x5YXI+lrt04JCEN0PVeysJooQO8SgRyXFpUBSKvcn37lE0s7axYiUjFdMlalinhGrjnj4PY
/Z30liNyghSpD974W1DW2EW/60D7tC45XDsK0YJRAKi4ZHn8OogbP9SIs4TUE//JShTXN6ViYtTY
1f9LBYndxJp/5+pRSUvPGv1EWjY45OOdTHgz628sIroXjswYoWK/29XBTeccth/E+FXNZ3DdGZ2v
eKyElxrCqj7Zbgt4RA4Gz80A1Icdb29kPL5msvpKS2YjgHba5kEw0Q0/q/ObQj4w/Idx+EvcCKEQ
2x2sA82QB8KdwL05rgRQbAIC87B+BrScLDJQpLbzLsoMek2jC43/8FyhcPgdpr0e4657n+nBNjAj
wMSCpMrAk52henIeUpc3yG28R3tCJnn1D7eZDBvVw9qxBBl9l+6fjqreB+ebM+QKLMPI7uP2bVlL
IOvpZSqyW0veqgdmgYc6UJ/teXVwtwsLJJyj9QcilX2OOL5eK28BbZV9nDgZsWVaiEgm0lV+f2fp
htmZVQVzeS51jSTkS5PkYc/71MrevYhgR9FmvcNeKKNoQ/Am7zWLyijLdj2mOqRiXG5pcy7MuJ/9
xML8omzZK/OafEIp6Gy4/MMl/qtT/pjbeAKrmZnBoKXPXBC22WJBzb7qMiYWPLPwVT93FYDzlRbw
4+AfaG/2FYN2OPI47+x4cuiFwWRNw+bqrCEVEHqsuJZVrsY5EQag9I/gMbjoaf/qiis73gorZu0Q
xGE9tso3/6LmX7u8bD2QA8PdO5niUNUEpLUBoW3u8V+Y8zrQVncYWRDi7CDFkykVqK2v4MkNUxOE
aX0easiLe1vN4o05Jl5pWIlQOcvE3nBxVOxdZmoj2vQpjSiqPnYvVnfSEEsbz1UpEc420j9FbfnS
Hu1IkREAhjNB2f6ZpTKFi20AR4TUDbyN0wU/eT6SziIwEnHylKZE1bORus2GOG8uLVRBxTvKT9hv
sxdHTAQm/owbGCA8bzTiqxarayf87o3XXX7Pl6KbNpp1KLRqVX1jkGZnwobxm9wO5g5y3Go21W2e
XzpibHAYtCl7aO8bhcKiRtFfcZu0i4hXDtfiyCwESmSIa75zK+RIHogJxi9Q2dnmaDY4jqNjr+lQ
Rc0PkxwjLUb2LAtUq6mBtmvkW6e1+BuI2RHou9s6U6FCvR+RAdmRi2kj38UIq06o3D6A9+BBYAJz
S24JwpBgXAd3KkmKqWHBngm72vpD63CL+pR3Rtj9jvUYEIDm9IWH+O++EXRCUsEbsB/j34AmJxwW
UV7cpr4IS3w7wQr7oLJXV6ppp8ExDEBSqt427RI+ZCrrLzKdvua9ysSbQvykvhBwotT8phxpX87s
u66Fy6UN61/+F7hWxK6m7P1LqK1f1UcbFeS7pRR5Sszy6IK4r8W1dzrqcVCqW5BjlVJg9QH0Gojf
Xu5Ph+u7cb+jKdsYX2AEnvFv5sPLmTV6FgoG+RdwcjddjW4H3UalVpR/ws4PS4BSsLEG/Avyztqs
OwK5Aaj1SN7aA4J7XvnceKYk4x/gS4ewaseq/14xg1eHgnLRKFW4hzjCYTVjm7mJGP1yWe4mO3Gc
DAoVy+20bIbMft8dzJsamf3M8h21JZoI8SJOCknHqgEvG3MxC90CpRuSGgcOL1bI2dXOOxhlYxRC
nl9NTD1Tkq8ocehdeUUc4fpEC8FWp8ZsUPGRDWKhxC85WVISjFFhj6Ds4KZhAV8v7aOrXz+ewdMu
2HXimSNZ4ak02OAPS3zl9RFZA3gcqpNyEtrQ3TzphLPXIGuoTc6CCtpKzMZGCyILXIR+rrJbrOk+
dG3/3yVPf/bQEOMYgUjBs+6f64ipA4Ey2qWf9/wv2KZsBaosGIuSVWHPzIVcCwIf05yCW/YPN0ET
09jvhjrQBZk8ZztqBbt7h8rQLhzEFAC9gcEzKKxscnxz+v+aMjFuLjI6AlbztRunloXg71gcAgZW
Vlbe162oY2BGDtZdE4Oi4fk/OOlzh8ZVe62iaR948H0SQ8kvIS3L3ZbqM6XvEf3ZPbgH4fnxIngf
Xz+CNbpxt6K/Y4QakKsJ7vEQGKPTb5080fZ3w9G6A3oIhOGGVHvJKUmGIYTMZnlBrxs0ot06eL7s
w2O1GKKjLWCI+HMY8KkgEAdMJKE421eibKTnNXk+wp8gxVBfcJAyLQWIL7jxKE42jcEOc0buKedA
a93L45pbWfv3dcOwEk6q6t44XsfwO9UhwoBo+AHMb3TcjF3K+q33GbZsQVJ6b+fjZM1pP/6NkrG4
4Gw4rV0PPEs7ytUi+I9Xt27DMeEFf/6whAE4XuspBN2kxCYd7lgJ9/0Im4LhGBPRv1C1Kum6gjQz
QDIjlZh53Hu0xkRjLnswH3XbyG8fmP0DMBc7IRXAQ3dSVkG0C0Qo+S5Cf8iBMCXEKLFz2cHdhAGO
x2fn8CdbOKl57pxz88Kra920hE86HwrQlQ0BTA3Mhmg64M8sUeFYweNVPQN2rQZMJ+zPGhRhejkn
540yqey+3oXIKhnovmqIJIRILeRPYoc2Q6mMxpVKdHaEAgDqRkUTDqT8qy2cDwS2Q/ROoqzV8OZ1
EFuKyfd3R3rAld0uBNEisTDusdXCTqEYhDYBAVQBb5KzVttlaVQ3RiHNpXjFRBwvyz9/95WrAI5N
7nB+wZUC0YmGSke5vWW2opagqrIBvsxStt9HTuHa4AwY2OkFudyqE8TbFW9ICGGhedzfxhqSmldx
YU/N5Ld23aNIPfDVSBS9a+LsvUbZuqOjhl/FLCWO7VVQe7cHKTuqPEIckDvDlK1Oeduk+F02QEAy
TbelNRoe3ckWLCXMUN7biuaFsitNr7PHRSjFNM3wCU19ePUcmp3/bBj3FwquSz+KHGOMjp+NPjvl
A/mzquI9x+9NmCcQcuiOWqLXvhJiwkyHWr7dTispn6Hw+WsF0dp2uhJ8MYTa/H8yIe9wr2lrvjVn
EE9ipYcduzaWojNMwHW38qoDcA/2OPX2GvTaNLibzanqrsuGkUdYFYi5r1D6Ngs1lHP1yH6f8TsY
ga9r/wPajsUH86vqShT37tsiGnIv4N6ItVQm6IuY1HQtvulOZfkPPG8jTGxlCXYr1jB1f4OgDURy
CYdKK+uQZ7JaOepHJjrZzoWRv8SdbjFAVsWEfX/g0BlzcnRanpGan0DmOfaLFrVXGYCrEUif7lYa
WrJZ56+rCGqlswAWub/eLHyilc/Sv+tbRqCRQnVvoZcURFk1/Roqaum0LYOUqemFLgh+fHgwrkvd
DsMu1Dvq0IuZ9BmhgAgifIXIXfJ/+Wwc6hCe3FDofacNhWO7LO9SIP86NrP5Jw98aB8jzMY1TrwC
CAG42OZuBhEbT3hqM3rcWrHzsUTwoyZzv4n9SyOxzUmdodGEFMrpTCd56ueUHqYCIWV1nDRNcltG
GoNjOC/vi1AGdmmyjlOSp/NA/XFM6NSrBvVfTG4Q1iw2HOSnpFxkxazVmZ8MtE5T6oY4wZCBL9oY
HksC6b3+h9hGf4G/bYTVI+iLcuVA4ZNYsalnE+ZOF31XxWLIUUR3tFl30Xi2xWxtAjvt0KsnxUaq
QVJZjF/eYM0+rmdsk4R0vL84ZI429M3Du+UUkPCcuDRU6x8hNb37RN4AtkEXw/7SBa2OzQ98GpQZ
Vobf9t//IEhIETuWaO2/jTrimHpNlEfpiFt5OeC2F8OnoAtwqcj+FZyQfUdSbbM3a8oP4fOa+siN
dujJEbBuNsX4wfm3DgujrYqlLBvOwje2lQTd+AJOeKPrrE32QlyZ3ZvIjLA0tQ4RD9zAwMsOXh/7
SaruP4wpW1r7CHHlj/8jH5poogeiZVMGoNzlHs+hDmVu3QDVQlWKjYFg4AW5K32USphb+8TMyMBq
qRhllRs5J2DEykd4Bw4UUlSUrvOZ11JO1jb3oq0PgwPjSBzXkPxbvWtRJwfL2IyvJf/D80zFocnc
bH9EdWkhXYMQ1+M4KpqSQBhXW230BN8e5u0JeImooLsB1h9jaM9/EwYll1kJqrRO3hLqfWxEAIrE
zmFNKGG4mRZSehaQlbMoq6seRHAaZss+M2CCBwcznErmO9goy6+EBkmScr/stZ7Z9OHd4R1N0zlR
WiUdVrOU16meRSpvIGVm2L1PNF0rAOonDTPTkekiQibGbDXPxlb821Zpwj0ofkkGRpc5qvbjJ3D0
6hWjeAA+wif2jkY8EaTK7kN/P7qNV3r0tTGvAkMTrovKmO+n6WBJ8LISQEs1lEoLb4r/671s4N2D
YCuen+JXslmUlsErs+pR+m66nikQq13YN63HFzMU6JEP9KvvOjcJesJlEu39C0gMlYILXRBRyRV4
Gt+eMSUCIuwN7oUyn0uxcpUH5apOJTyNvcSYeQFQkqCl61lgiA/sEEuBMFEaZoYDRajb06A3dFvB
UhMT32Gxlr9WA4TZlW1KkYyYAfy1LrZKVFiVivUKe4CUGFzG5WxzOzNQ0VhKzoh6PFBg327coHyV
gc9ETGOguJZE3WlryuDL5Fx2NjzWiIFkLJGhE/RkVOAtRzePcD+ZKEkF5cUrXTFK0+w3MAkQusfK
0h2+nWYnzj8oEx0E6GHb8tEO/OH1q9ICv55X7s2j5lsQYtJFMNDw/MeoeJv9ECZDWGb1Bt5R/wxA
unOYdPaAYDMlLvgB1kJTJrlegq2BIYrGU6vF1Jt76wrT/81h+ikmP+wWACEurmyZTuZVvSqOwzsx
pHWTa72IC8tKYjLAd6pRadeZJhSumNhZmxuBv+QNuUdXHPFQDIF+JsF8ZGIjTA/2dcjDeOli7KN2
Y79Ufs4z61Nlev9lkE3k5f/pEnIfYoNsXKfQQvGwUTDkfdzLIX4OYXp13uBc4sfEALW0w9FAopW2
PlyvdTIuEfo5djrZhSM0BItRIjZllGP5qG1buzLp834b9J6lf2SegAneO/9a2wmSTZEM9wQ4osui
flF43ygAhpbjVhHAMgXzbPK/KyAl/ERirvYQXmA/8YOZAgEvDIJ8TceL4ppHoEF/IanUeS09Sgzs
AJe2ruQj6x1XC1jTrJ/Al7Ncpdwi/iLqAzafxtupwzxqo4zZxAyEKd0ZmgL8bU0Sg5/PmEl6jG/g
mYmCh1RWMIlHj3XDC6XCqMN/KSUZcNiO47WJrALgAWGKfsGtOagzyO2hXKdjANY6wDG0IvUgOwsN
XOPccK3lZn8D8MIddrCLQ5u2YiWaNfQFyfpzN2wK9B6YxVBlqOwXFWwwv9I2+lfyoWg51il6nigC
4lgtAWOFY0kP5y8lZ4SUIi9gLVYa74iZKwEB2fGGcseuP2ocQgx26qAdqbaKtuPioX5C2E7T9Afs
B6fpkIZeHpaYr1rahS8Y1psHBWSL2otj2jgZuNZ21ic77tJiFOiJpVtAmhsG9Gjy1thf1rQ7KjuD
ubly+HRl67K9NRJ0oyMcu0J6h96clU9A6ImuT58i8K0+47h2uruzXsEfV/C6+rbCkCbtSmCnQYxk
ruyuTRpvBAEbD0h1yECRe5pzaIcEcbE7x6/5Ad695xFyMFLo10Jr8UosMaxNpGBhxVibBSarEmqZ
Q/8MX87BF/HHkNhIQ5tUhP8cfluaZpY3Rx5INhLOIsobby1xVFpOuQyle9YrFp6PboPG53PeIduC
6IGe1G3Y2mNfjJJ1ILXB3T0Ja+lIdHKHiHyXsacGf45S3dpyC7Z8oxyCm/nt216KUOlLmtMRLush
8rQIEMkRp8dHkc9pPFCbu4cFcgU/3RFF3zrv2ljGmc5sivfrPpYJSO9I5MEjwpgtSsqVGZohheNh
6qdt9RzDlcpm0j5VCBopiXze64P+s0ZGeX0iBsWB6g3ClzMsq5PSK8bHz7vGwKtP+hreeDmjmxNS
SO46poBsRFqyuCoLXxGyVV7F74cziszRq9xBxHNksPFGAQGd/fX4TzCtMlDy2WZJbgl3pT/tZyAb
32ZPGDeF3PdvTq+R9gO4n9Huld4ZZ7K2XY2AR1t9+/t4KGBmGP0WYF3P+16pPaJ/VPM0fh3UG1Z1
DQahissGpfKxXlv8sZGNaqvLc1s55xbVjsx6vrRDEdeFuTLpeHBvGA51QYvnYUv0f9mQao7TnzFO
MsI5xbZUurnvXCGf0NmPt7KgeLg3F2/Uu/KwOdx6lepS5HsWbUEmblrY0YI/HfjY54wapQNTMLii
XNpakL8ZCwP1qlWynoEl+4Axr77JGX/MqYDRMsbWMq7eTg9umfKh22+HXc8H1cPSmaItu1UR/yOD
H4bORU9JitatydIoNRBIxHiFD6/Jd6bxUt6199GWTK6p1ZWKNLtrVFlj38eW3e4auqgS8Tr1gYi7
bXLBDOWRN6lrgPymfcEPq88x8YSmI9kdVhJcq01oJmOrf796jLfHiuCCR94nO9p5AcwH+OUKPrz2
ccWHg6rMhviE46zUo+/5rfcvsnGQdpVS/2sMS1XZYBmrlf963HIzBH53jdxMP2gdWHNnIr736Nyf
K1bygZTGNmle4YDtic9eknw5CY2Q3lmuExpV8/V+Cx5mIfGOiNgvy/eVp3QKr0vZ9LUxfTJuaO3q
106lkskLK4ZyfDsbGRTT1PsVv36pl3A3klEYaHaRg6wlSH8eQUlyvnJjK4SqbUhvWsUnaXl+49sl
OtF8OQl7ZRHqDEMXNmeLu1OBLKU54VRivucG7NX5gvf7MVClrvGZnAeZsuf4ylB9L8dcth4sxIPD
4brQG4bhwYeCRH32geI4sAhhpcfCCl5kUSmWuD9NWYJJ9vO+3RNCDWbhnSwci4WLtr4rlqODm5mY
jsCMlWbrxd+GLrnBtx1llsNxDTbcLlg4qUZ7Av9n9PMhZBcDWmo3MKLXWzUip1RHsJzKU+TgLB8h
2HTo6Rjho/ma5ejoLLYViqQ9s1QQMDIaxShkLE/ouL4FSJAvpKdus60Se14hH8mPhjaUWSvl4MRR
BKRv9kdIXtA7r+mFEBXHucZ0w2Xlx+7SbnlB0M651LSc3e2Qfuae3DGrHW8KN4y2L6xB1gK5EUBt
wNApK96S7+HgR98d1rDM+q8UL0XfvDNgn84aIKhuife63EIXhZ4rjiymuXdiApR+4QbNR2InMTCq
oBPFD4vDwbs8BorFWaFoYnisfAQe3xUaWUO4gFcQ6toUguvN0HiMe4rhnM8ecFSVB/i4DmNcLwG1
3DVzKPr+H/ET1vR1uMR40INnxHAlxeBLS3zXY+1Rb6W4tIyRe470Hyix3k9XpKraYglIcfJLZyTw
DIyn+u01RkUn9f9ZZcR9os4ULkgKvJNoljkKbqfBJzCho9ylZLrW+w24W5FS7IpMJNd1zHhi8qwE
uX8iR+jI904dlIBvITBK/A8BJWi2by+bJzW/IlC9gJOjC2PY+7pi4lbp5BY0XAM8ZFHj0uTFJMlX
Ho5O4Jdq8XQkSI/QszTgAKpqjo2ndg9dC5e4VPzPi+/sQZaIaiPGW/pW2cL11W3sEHQhsV5sox8n
DlwTYK0QZrifYCjXA7NmjR2ggNEEGteGCr6tz1ncwgBdW99z1CsWNd3KKzE7CvFB4jlu+fXnnrSW
5Xp0Rek5WBkwWttg5ojZe17/03ISSnjIxHSY8TE/Eabqg1h9IEtGhgr7PMtP2umFQ2O7ZY0W3h9w
d3mSqtTeqtVDSpyGHS/1LV2G2WOW34xaFnbmpNnkNDlojKerP0YZ+zaa1wEhj41zLji6QIFBNgaM
0JoFbI+xcvrKPErpy1E7FlhM5xEDYau4PVfUCyQpbxfemqfVvBqgDAkxbM18+J0X2r5XRF5FMElt
lghUDRD3hVACzXyRKLA0zp6Pf/BJZFjbXmudKb9v6NaEfvh8sqymZyFfIwtI0dHcAFBAttU6gyhI
k92iiCSBW0VKG/Z/BRqsqhLbTD20eXid9Yu4ZbH3uVI+Mt/8Zr8ZvMMcmJg4+9CCJASRmnPJkg08
tRnwg4ReEj+MtB1bBd9aTOUP5tRLWFmv7n+SiW2d518SSUVw2d1TNwMOD28lOvcpHQkoFxnqDZRe
aB1iOwIKQTgll6X6faLPtKMBWFmoJB+1wjsxKLnWvVPXQQ3i8/qHAsnfzFPdZrBiJW56MdjjbJAy
Ckz27McpVJoZLLw1h5pZZTX1JLhsNwYS3xLESI+vYIZgbM3UY/XP2k6/Aom6LLR24wmDxN2TUly1
bY95jEzL3t4k99WhChs3tub2Icfkw+8ey9WTuNMqiGpmlSNr38VWEFjjI0AmeAJsAKI1BFi/63uO
htjHmSG/UtOKe7feTso2gltml7jTdmC9SgQxg77QYilEPejBlVKsnnRJKRynZpX4XFB8lSOOgHJt
JRdTIhfQwSXQTkcz9jX27M7sau0LG3ALdnx4eEUgx7ogkoMaUC0KotoZVcHwVMdHvPh90AkwBDvC
ewfnXK04uCnEf6EUXxZycvmQkP87Q9yrdTaqWO0mfEwZAJEYnliivKMAK1VnXIjB4xuUnt/o+emY
ZIY77fq4gZ4UjGIU7dTmZr0ullO/VkFulZdoJxSOJtigeTTr2ZdL60ZD4rd3rmUwhqiHUb8I2kGr
AKGak/l4E54MUUDjUFbSByvggHT5yY/fpYylGewHQ3DCoOX8GunW6QSxuZvXCMG6+dFmBni41q2F
f+IPkjK365xtftmElurc/JlTkVUlHYKySjPCGF6JjpWm6/CZIMk9Slj/JnEfFS8XnKKWgJyNpayl
25xCcU/F8BruGpg1SU98G6g1/BSehzHNNgGzDOLsONKdyRy75FIsHxeFqOe+EQYxqwAF5L2eh9qr
Z7Br1x3CGcaCyzO3i6Oa83+F7RiXeg0Fow4xCY4VT1tN87pjGllc1Af8ttt4+6XcyDnIPgJpz8kD
DBGhLAzbYLhvoap6XcYQQs2Wc0IxrJYpu1unfJVdib5SJJG30KYndiQIUdSJMDbtT3M9gpxT+fEC
CuMPr5FKpuNG1Kp1NRyHyxM8ebLUAn7lfGPEJ5hzcXs7C3O7V4QNHZAunPHp7cvC2JrHCpGJOO3R
4ZqTJ793a+zFN3d6A6tJEphpi+GrOFdqcvaCZHYbx1cK5E55noBiow8NnHfbVxAa9kPBTLT2Vb2w
V6lXjFNInuM8HWe64Tix0vMWOqCqcn4x8VZbs43A+p33xzBXBMdCWznIrr78qtMr9fLxSTYqqOg3
yaWvgsq1hQrLKd5rS01266fdDxBsKxbOOncv40QRQ1ZYwiS4k5jayyvWwKzbIeZfCNVqlkIKQns3
cX0r6eMyNY2eYocDjdH73AVdMLJL8zifOvkOukyGBEGOBOsV4wM5xNfko/ceh1918YBmDZuphpb4
+M6ubiZz+LtmfxvAi1yWbmgxhIKF0aD+3tQFWWTHqFxD3e/S1rIzB2/W9AwsR5vXP50hk5Pl8tB8
DqYxZ/OExbNnmXig60NV7cwIY2nQDCworgxP4O1C22qsu2/f0hy2tdpmEV1VBxh5d3xA7yAWAObs
/H5AxAppiAS+qJEYFGS8s0GTgrVFxuCDBLDUgHWxHYthyMMPn4OfQhQ8Am9PeEi4WGtWGKye3MBX
n01GXZZydijiFpRkJWW1EJy6R7AFsA4isBRIiaFjtLWMB3C324jdWWGFNouJfafA5JYEwbnQJ68H
3x4oOWEp7v4Yi/pnQdv7OAWAmSqxXucqgQqvcUrUimBa3RLIa9megVstbEa0Y8EgQLmSZgldwx22
s4PgKXNix7AS0SwO5qoiFkfAJ7y4heJUFC8nHgSivyIdwrOC4fn6SC22v/DJJk82lmNaeKbOP6+z
tw7cFDRRG17gyAgXm+CY0hb72hCz7u+gOIX1XUEI5QpAgcCIPaEsunR/nLYpGLoub+3h2llVLMJf
nWjvVr6eHDK5GKrsRh0ZGdbeS6hKxeFLxoFdfXSuRm3NSXAxk/GrB4ByG2aFlAhFIC/5GLnxYvW6
Y78oUai8UZU0cQ+6pkfidhnA+kc+0zAmZgwCu8dvKvQEuO8Cvz8txgNqAn4YLYtCXhVxemdOW0OK
YI+F9ycDVQYmtYLn5khKX11DXlszwQvBuPCUUECkj5Nq0PR2thzbhVfdc5lwDpaQZdQlfnFj/5CX
KT7N+IAtcYxqAoRJYgsnRqHp8hhfpCi1frXWAfm+Cg5VLr8u+UNbdxGR8VdaiNuEOE/7nF4qtEKT
QXAxI+vruroDCBC6X3cjEZlKE+g1mLXZwYB3gHsigdxwMw4X7NBN0OyroLJ0iJOv0I9wc0oZJGTF
uq7JO9bMYDoN+sjupyde98cQ9O3DiU2+NEl/1i5Td2Vq1qzhn1k6sTwzQyGDozkBG7SabCwSBwbb
h9oHe3nSSd5t2Ri3jg7EXfelTDVYVXVv4rXrPbryXOA8PRNog0NU9kNndO1/vbxVSesDDJUl1BdQ
d4LqzVGga1B1kGL4+h1LDti37V4al1ErELB5wOWGyJVs5hxgTZC6welPXiy3DFsV8ezDMNVpL8z1
QgPKHOObufExWSg9qyg55nHcq+3WEPF3aJFyLL/T8rXPzsxLtdMS0B9g4iYX4DDDLUi03D7ZbK7y
l6K7Gx4HcFhqJVPVfJti50Kpx0NIy3wapnscPfy0KgefgG85HmqFmcakTML/rPCEqr1w0t7pelgc
80H0Pqwd9P8s3hl5KEgOKSAW3hOIqWmV4qPQvDppBoRZ/xs/ey2XsjAedqIbheRbzQ1z/l9xX4nz
8YO4Vqib4lsTH3mF7oqYeyZNtD/9+sp18Ku4y+uqda6YAw6yE9xjbmUfC1Cw0Wd6LhsqDxXi+2E2
mNsDURs/DxhjqeGFOFuf53Ij2EY+qjgQrZYtxbCXIq2s2kTQgBsxiVwCWcv+agCsEY1dSOvwapYf
/4gIq655iIyWgg82ynJpZXsONdsmtOBr8at2ngxvIKiXSIU38zBoIzcEz19JBHMcLAL5zjZCH2nf
r3/vO7NiTAuHDtP6V579J2GnCS/DJTb8XgE5NNUCcqwPQd3pAbNlpSvrMPoAK9YpVtUiikDQ8875
Jx427++9lXmdh7py3rHoD7ujbfgvB8OH5WnwmrsjmE4TALSZ4ceJVh1HHPIAKoAFYkgiqlwnqwub
cjf8KLbadlTgt1F/GBTSMcTpdtTT5mY7fasysvdZ8RCgaMVTxkBUrxkVPplqNzDEiKfHbY3UYMiK
SD0T7BzmLVFmOGqiWRCXamEZTL+NnHIFdq2rddx3B8ig+jlXIGPHkkV5ozfBHd06Ip71GeyTvPes
WnvKcYsptbso2DWMNvqFgkKdKgiS1kgZGaQlOKoMFh7Cur9cpLj8scQRfbCyG5mg9x8/e0i9UriL
MaFzMtvfV4ETw6nQsZPaXzn20ouL1NAW+1LJ+ZpymS+gw1ux3uBzc1pG8YuEfwUnDdXebAT/7vjf
FhLL6IiudvnmSs1EAw7kKMu05Vv8gP5oOlOOcyiatcaqJiEUejRDucVxPzETB2LVBmA8FWb+ivxb
NQb97TTBZls2Zri1FVj5DAyq2KSrjVGAQj4jNNFxWepmUWq4n+1p2nEnEs/hoU0OhZx55d21OxKl
IdwPdS0edFXG19DA1clLjrTLwDv/az7NxDyR6sZi1K44acZJEMrUT7a9P+mDsaOH2Iew93ur7Zl4
DCkRb3Rsp7bcboOIRKwRVhf7H58anrv2AdGCeXEcW5VyuvSIC6fnnpUWILnzXSyHWzz1W+WsflcU
4IkpY2MDDGMkZED1SAUiEzd//0zAfE0Ibi74Hz2/6/COeTRqshAeQn9oaeSAgXEupZJt/jtmsZmS
bbBdCCUasRYUfJL6iRNdABjmvVXA7ecP4z4fe+i3JlxT65c8Rv0QJRiOMdSXbYR3LSp+0dXZSZkT
NSdwqKGXoalggaRLL+wblsxgzkWofryDPWickTK4wfHDdpkLo+AVXGFIbZAi6rKoCgsRVdz4Bqnq
HS3i8RoYkFKSwfGlcACvXIQGKGjZyp87qhaKb7MtudS7EemhhIpv2veynihnQ7qZAQYTA3vSL5Gt
g9rB5wfhTPYfn7vYue2qoucN8qayRHB7pNYUxnrfaF5vh6Et1bADMA1wzID+GtlDCuxcNYH5rZyc
QzJWRmNJO/ZXv/jMYZak54wBj/267vAXBiUHYoBRydzgWS3EJ2sL6IDOeM/c0vpJIPL+s9tVMe5r
b7oL4R7miSOsBY2aUDzh+4fnRZjPfvxo+S+d9vuGZauOEOqGoEmzL/jslDMyyChSwqfeMFqCEAej
LyIumLBZDtE2d6xxrxy7cFqlndf+incGz8JApCfxVmhHKBbKcT3b9aSNzizw9oLtqVZxih1y700C
YznL/NIzxxlnuTzQJMUKrcLWpa2OSccs1vmF+YwTw8q55kKhN9aRoAlwh4UreGjRZROh/esYGdZ4
e2u98mX09V0hJSpXPDH6T4DoqDQXGe6gsRsxd5lF+C99khfXh4Q4kEjLEko9eCfdutiG5ZuofeYw
ts7hwYgysFxP7ZHbFZjdJIHa7A9lRUYMU4bKvy4Ju72jENWtu3D3m+kZGnDdXhSdbP4Cfg14JNkc
Sow79L7j1vA9ydEwwNGwtOagW09hkOtS4dXh2mstCHkl0kXh6p8XTLa13NIHmx9QfdniRK60hIUm
856zBSxndZ9d4beFMRDaTF5ymMXavkZVczPmqNOH5VDWCNieRBsF31PmEBKO29907InfpmECbgcS
745P1EADg26WL6raxfSsNwmAEEGbp6fEeobB4wDY0+Tqu0/KDa19Vveh5ZJUxZ4s7suqlkld97kU
ziBcSnT8phKhtUNdaZxxOy4YdgNQIMUV7U9mvEpw308R4iOJ39cX/SvdGFJSR4AYevoWhWZ7+3xp
MeWA32V1DFdY2EOyaQ+aLPCNUn6gr6i817W6AgYb8z63E/W9sK0fAXKCmxfMucWEsmqSDN39IJgk
rtLMecjou8E26BKjbNctQLtkEKYttRgysuJvfyx+FyUe3Vryl313SVkqCWDstOmeeD4oPXqSbcnu
viNBAJCDKFXWno9F7ezuBLggBN0C0UufLL83DwRb/OXzeA5mwFMyvpoSwnO3QRxWxwzEj+lLFMiB
1BbwiKPFyACGojsz1OQedcXfKIDg3JcfNrSI9f/ANJt18AzRBbKku1ZdWqGrRtvj0w3po9kDjDEJ
SCx01qlSUF+usH/PrsE/664SKcnel6Ip2Dria1TkQEaOdM7TiTE88huJfF9hzAWKJCpM91AUqci4
WvYfCD67JlPJBVFYd6sNyjWD1G+fb1UZbcm1NSSL/04ni9ZkM9A0aZAJUh0GuCWzc6pVAMsh2zfL
BGuZQP9hgbRvuoRqap3vk3AB7ZRQHyJgcfGuiFUtPv0QZ18pRN5ZvJxn1e/+PYsBRewXBOOqzHF8
0erXnCFxIIOB6FZGecTT53lTPyIG+xFW7IJORJlJ932W4EsfsgvN3o0VPCexM30DyhGZQ4gcuJ5o
hpPBfy6zt5WtaRpOmU7YItBUW9XPCroF7m9MYZJOQ00H84l4/XDt0TxJHE84H9Ne4jxJjQlJHoWo
ENe/r1xuRWXhZjxBH2j+vlg7MOWccp/6VjvA0aLnIdta2Kn0o2t49fHBLUgLHBtORwQXj+EB3u2b
PjcDZk7XAuSYbMqgmHfDQuXxS9sVUqJX9MCWzlu7BQo6v20p0J+WpcAiqQn6wsFZPEcEvJv6QYd2
058v3J9zeogycMk0iZJtt5PcDOsBXgI6/ATIZc4tP+kihhF3+6TtWoPiLtDOquGbRgZpA+lm8+/R
8p35krkAiA04npG9b6D7Phel0eO/01LCnrJr0CQD6US35AwXKqwof9YQCovZoWkrvCub9+GbZ/eY
7wR2602f4iRpXw77LXh5nK+6rZPHQDPM74nHwcTMT8LHJgK8neAC6tahMKyVb6vNIQgK7dCJ8L7F
odfNYLE25rRB8SuAtlWnZt4cZRiT1tEK9t+2qcm3jWHWWlt55OPBvARyth7TlA7zkBO9fXY1UykJ
yS/u36ezuSkiywQ9GwfjgOr2bqBhD1zz2LPP+YQ6l1751uDIXUukn6Cw0ZiPXl1/M47f/+PYU7mF
tp7Ow9bSfoTvq21iHXFeD58r7wUO1iRU7AbjSAejdvVNsxKdzerYasxPWKKcZ6zfgRsVcqrVDB/n
k74Pk9nuzgXgnbWbA3jTswAVhouWd7LcGP/4nkUztpPmdjARk80j7E0aKs2JMjKuqsKE4+J9T4+T
QFKf1aXYPkE/dRrFYaOZoBMwQhbTwSdoXwwnvTXU/BLtKc5Pha+3h21F7C1GIgDiJREECdfmZV0g
yCBbxQxiXsTUIgMGrLaer6WruMpbeFfqFWHYbxbA7s5nzgKAnxGVace1+WDnJOoGYjicMaQdjMEi
DOJEB1UgKCIRxFpMXHWLJcUZtsRgQGO1zKmoc8j6vOnoRD2u3Wt5e9A4ilQGxr+M2OXK+/NHyqKB
AXzkxvsQn/2i+0aFtsssrmAFUtV5iu0t9lXbsm7eFNNi055MHyYCxBd7O5IIzDNPxML3b72zjbV5
xg6cAoyiUP6IbwdDl0+rr+ITS0hNlkH7UdDS8Jh4Ta5YH2kAsRpdVl7nzEuZ2FNslS8tYoY+FYfC
eDTmDylhC3qx8R2b9AT1PSZRAtOpcQpc8P2asyUIq5sw8B5rBqY5X1hPCeyXjXBnMWutSAD+CRmF
UikHSUqrU1vhWDjxsfSoglm73BYfIGbOmNl9MgMdVp7bcHTjomRAGuCjDcGUfOdOmxHEjNpxCcI/
yFVrz2jWnsUIuuHixRgmR/EzouFqQ55xv4juiA9BmdUp/96hCm3OtA4wqLwuO9AHV0nV3uTBIe6Q
yFD2J4sXP6i/XpiK5jEF20Z/m3AbuleLRxTnvjdNG4QBAgHg1cfgR5a8oTmYjU5WNpYPdq5t4hz5
sPOWjqEjBfk7zCODZ6dgJ/WeS9rlMyYMc2eo0qaojxLdOoq/VZEWeOR5dY55WBLQE455by/aj5Hg
5tET9NvlP8TGKDKoAgf4rnFRZcGK7znOHj9PLsa8BcKcgYlStdq1KqMdL0YnDHpB+cRaqiNhEhTV
aJRWG2JGuT3DiPyUo5+F0FUKTmf6gtTBejr/ln21Wt0zDkw9hv5QOwKROqBeKypox1m67QkmNRl8
uK4ACEbQm6MN6zOLzamtAXnCxmiNMDmLEAOZM58z83LGwFJSQCLV9Fn5z/naIQ2xFAnX+2p7jzSI
oZMK0Cs/2uz9aIIqJxFijFuT3itkK0e8jOXF0LGDHDyIeTv94OeNc/sxpR2whIEFnI1RnOpBu1+W
GVYoFNKZp0eKWaHqF/L6tFDeYZT22iGJ8eSM78M5HGozPlt7PzhN4c43vuqbZOZRQfip5COAhMwA
hOvYeji6JeJ1aCZoCtJSuYNFnlYJn2GHzN1QWiAdkW0xFWKSNdtuC7eemaKLuc15frLuThBlnheP
zB50JJm52zUAPuKrp0bjZip5gU7BrhuaaQ3rpZ4EivFfpZMy5OpDsosLc5OeSUSHI9I/wPfyOqAn
mb4Chnal76GZ0JFvPF53ZQQAgsF9UW3xf3XzT1kpKqB/0kdC8X79KdjqEC3C5qNbaRxaU8MBmats
yC4LOoPtuMvy6XgiSQMbeL/cwK6BWPbU731uebJE3fJK8Z7ebKLDEBWmP/PVg9t0AHRjtPmGvj58
ZJ5RMxVflE7pSQGsb8JXdfHJ8SgeLG3B5rEKbvz2kICyZ+bdGrlGY7IvvcJmnEW/yqSM5QNkxvzn
81CXst9f5cwba4/ZJCcQhD3lUY9MPmalhJ+TkNdicGwrurOf7qs/wqYqQklYM0AbNGx8BNdtV4Ag
Pt5B7MkxTjFsgmJ5EQDM+sQiyzBQl+DnIUvT5ocfa7f1kzr8+s5LyfPMcCgUACBwMARP+sS0p26R
T9X3m150QIygKPL9Qhv6xzAwdT4NNdZ9I4THplyX9DaqvGPhU1E4mmiBi7H+y6FMBTowZdxqTMLV
XGlEAlXDogzHD0sEvf4JHDGp3If3Qy6zcJZNIeWMIu0SOabYcRgatt9UGEEIS2UkpayCdw1EzpRT
0Wr7Lamxdvb3rI7iYGKjIHujm7HEgl+yX9Mdqt/55O25OWePPE+wLdA8yk2SVQYUOcjc3kdmkgNH
Tstj1qLPPUZRTY4bhBxykV7KspFqnJ178ljS8U9pKGN+jIjzuJ4vdf2E2psAYUhC9FZWdbulTwIb
mXZFBGm6sLUPp0BgJcoQKY1GjOGBFgs0K3YeBnsAecBCeRrcVFYbWgT37jtG8NCkAkul4xICjfku
X1A4vl47kmzgGC3NVEx9AU/AdAzTIrq6ksBm0lv2DfDjmRlGvG3bgkr3TjkEhbw4YFQs3/V2jJbP
FKxlu+i3M3Iu/nwvB9zcSxpn2u2aRtr4+zxjLGCkcTj4vPaqW7UQ6OG36Lhgx2cGlxY4KH7eWgKa
/235dYWT4laPLp3v+QB2SA3AhaYCnLiPrBYz2c8/vITD2asNUTQXz4Xm6Qq16It/VDn/z2sNhK3R
SyNvK+AR4Uc06/r+9tCTmQDvg1bt0oCTovSTGIXl23M1z1iZpgYxleLjBQyLhA3rLFeqjiq0i8qG
rrEB61yi2fsR6VY7k48asCnosV57mjiFJNUlQfaj3UuEmVZkyVDxITHCecMHzfUJ5C4F8VXPzxrQ
AGYStNpifgIedtr54Uc12bFLJLpQGti92FnWDqMmgyu1+m9RLXL7O2+h8oqb6mWoMzFUaa+YZuVx
4mOQtqLL2IFLiXYxLQGb3F9yIo27F/Ul1rgqCymX5nIflBdOjYvZRsnTI3aFC8fexEVGY0wVV6sQ
4QkDQ2Vm79WXeN14sRtTEBp7Y0R2Sy2TbBK6CpcoTfvRYKjiNhQFwUB4GC9AtkskHSuXV0QL+NA6
iVkPtW18VwGnY0rlefa9UCO3Zz9uzTc4Fu5Od/mLdYF+Sl43aLWCYNfmaYmbV/AFBliNlTlWHu44
iCDif/tmWX3ZpkBO7T+iyEIEI82jQX9TR/el33nbkhFvwoe14cqXZDQiitYuaq+QiHvZLzKgvn5O
ESfJQm5jWqX4LJzzzt0f1pW4+qIQZ8V286WQseHduHUaWsOm4IsDnGOdNK0NWP72yocrUqTfpYfv
XIsOkcbc0c/h49N+a7GiW/mfmrrCX9zU3w5RA+8suzuzkbQS7BNjCAbC4eo9nRR7d0xigs+UQghy
2NzRUJL8ZnqNtu2/t0oECX0+d+qlgFtxy7tqJ7YemQMErIk32P9SOU/k7Xs921t7MxlfJ7jwPLwO
kGvhqIT/YR+cetjJF82o4Oyfb0N5W5QVMrwCxeFw4A/WNrOTM9w0ISoLaHCrFFRVvzQsvUfaHNUz
YoKpyH2aQ1XFcQk+S77TiqPEhaApHPuXsLFTq9eHBtcF4j+WJho6Ua/Mq5mw/bHoZCLIcnUVz9gS
AGdd+U0as/bSxIVJNp05CJs4OqgxRxZbEWi4F3JqUM2NrldNT6LJG6K7F1g607M1dOdLS1gQTC4J
bwbfbDr5D1Vc3ZRpWss1GPd8rmehgvQLEK+OrEYj4Y8Dp9/99AHIJNXlrRHvmFrfxVskEP7X6+4+
1O7Ccxd64S7cE0VtmSynBsSw+/X9Uc3oonAXmuLUG2CRy3E99/4+DohleGYX66rS9qM4JFWeUn4e
KT9CEMTXCaa13jssN0GbDExb0lsLJpAS+Pdlc0/ogryUUKhwTCF71d3Ds7plL854tw1s3pU8tq0A
VOz7/gzeftfn2u9/JJAZ4mHi9t4jODXdSIscbC063DGIF4oOGwYy8KDUhynl1J3C8X8zVSnAFJnr
dLpdEW3H233+p5KXG+RFoGnXR6HjgpUudj8m0G2z70mLzStIqjIu8Lvlc0jScJwbehRE2im06chd
9TdSxlikjuDAzZr6iSdNHxiOQgFhsrdh8gRrvUqP6AjDHRlI5anP5OGoHpRdDpkYS2m7/S5ZpfZv
yTbbkGbnQ/pMKRVi35yDELnvFO6xYIu8js6oe5Qcu0fMw/HwdJvUPqa+E2R1yX2kRuo6H+F/LjC4
DWVGfBInh8jX8NM3NwGP7+7Cu/nsEOQ79cQ37Jrsal6767c22XnPn0QkZ/CGpXXkaZVVrvW4OFYj
WKj5EPbBtuTk2xIdcFhlCjnmN4eWYvdTVidItCKPoX2cSL0ill8RrSotF61DXcxBgvXLVNUfWAqn
2A+qW0jaObUcl0clBN64f5/QX9RYqEszZ3/q29xaAPbmZZ1Wks2iJX0C9L4UCoQUa3mk5e5VJhf8
beaibVeYOrPKI9j5criW996QxOK/93PuuJggVF0m6uiaavoTcthUGFPC6jZGYI1eVf0idW7pGLpw
bffg3v505hz/DfxvNhSuGoa/LeuJI9zjKBQIV1c0CZzcf07tq3zv92wacUudtmSVE2hDfrDJRga9
WoQmZxk2gBWC85UoKCA6SucnxcArZktVnXwRtIlp0agMBMBLIR3U6Gwbq5eUIvAUe0biPFuNPKoS
badUYnsRrEF1SxD3xenMFXKG+9dBzZuys60mQlsmLvIEwxOMnKoi8UI4RQ7cSobMEdMLr+EoOPgT
7HnG46NNZoBaixuZvqVXTtNm4/8zYWnrS4jAZPFvASdEdXmI5f5bi19afqya98W7cW/S1OB5wsXq
5vlIwDWQaCX5aGD67n0RMR3k1foLwn/64X014aL1y4NWHcaTHogjwycC5fAB7r6e2Tu2UcMrXe6H
RextmHsfkgmiaXhofWvF6gIBbuuA1od2PXHldnDAg4MRzjKYyrCDcuox3UF7WfcRUg3Ap4IatPfE
WAjJuwEHh2hg7xjhNmL3CpmMIKqJHu9sG5kH4PE9Q8MCiXx8o3W1xKGtAQokkctj7fE+3A0lar3L
2MPObRQHKsSxwgAqzQ6+mHUHnuBbpJHGIgq7DpgbWCTAKS1QyJ6oOToiQ0PuvTc+kdbwjFpJWQPS
9O96dOpROsAai/lf61e97Dab0XRAMBAepeIcsoAg3VOik/o5Xr66mBOWcvO+BpjtukJQSr95cLKq
zOgoQQqa9KWhq1xh34CgIitwXVOaV1/NbDP2SREJ31vaCn1IsdJxNJ98J6Nu1XmqCHyn0/Apcz51
wqrIkL3TAjIbnAmTWhfDhPuWCEaDqlgAsOBai3leuWUKRSmOKlGn3j08Qr6MO+4TTIaArkh/QXOc
cXKEemnND13PkHMjApT1BfzlBVd4U3u+Oz16vQ1TNpTi3PXlTTcrfVQkZSWmnVWaKfoOgryEwY8q
FlKmcLPNHxlzR2f9XbllNqQ8IQpFtwhIdrvXxa2C9NZQ3XuPLZzuH6YBYCV+6zqz4/LK4IgI9IXz
mDf3VhHE5v0M17c/fUNfUddnokHZbYv4hO5am/mrt5OZVAtDLySMDwE2lKhmsxNx4Ve3DhcYvjrl
IdVZ2x+gzCikHFGi/4aEDDvjDuDifMDHsh2jsm0AAppZigtJXqrQuuBaRvf9MKAxtqNmLgGo2W8L
S7x0RT2j7JhpUKvpnK1qDmXEvfAogdfb7CQJwJWh0b+LxtckCOyH0/cCmIGuHIK4SYe1KLrsnMw5
GZlkgKJvaKComJzw+cTGN/wwux9XY3hg2NTWCXEKF6QrWnqRqgpzqP7mbY0dZXejvEklJyIrGU99
rhGGPgcAmmltzEMWIiP5sT+sLFd51f/aci341LNGiwy0FC7RFiIjMjyoj1ZnzPjklEbrNCNmQ3cm
ZR1WiIpl2c+A+h8cUGv/uCsJd3o8A5kiZ4pJo4TBF9H7UZ9qT8eatd6UzKj+wxGw+t0Z2MH5rQhZ
RsZD1erKr4XLky41kYIveOSFc8wlPwrUs9p0moeciAr8SpsO6//pcUtSKL9xDB8SJ4EFtHfjJuZ6
L9Rdw0Xq2HXszjgWejbg7oG4WJxerbAwmzAM+3ofeW4tdfKjOoqD5zWbBtimCVZw7uqA89B5Hnau
EpIo7MbWy5DjeqAWJMCkh73+w63gjJSSCvRV6XvMuzV8zo/pHi1oJN8gXMwJz5XByKlaCXZffnhu
GP8pmr4HXiiaNvVkgLslwXtNPjSEBi651ySb/moLL26zuPNeFjkddALy0L/c3L9YxNgxj4Lck1Sf
3cM2kYIyXjOwjZf3r4UpJIHLNtcjEmI4Ie1XxNrLy9Cw/udwRxc2jWxMCEjQRLMs47v0uxIh3o3n
OBAXKslWBOYuh99KvdUFeTE8njXEqlfPOhSrPwQvQ4h3blCyNYWXQl/0RBdj28IO/zpYYbRM0WXj
H/UvKapS+47T4n8YmUS7ZlvmcrGh8jXIC039JuFXVgsNE2Gta861IdopNWx40bR5M2463E/wlLdd
iTDqUCuSFCNIOGCA768uoKB45oeRNJANoI5rxOF7GbQeRw01oOB9eFmW5rOymS4p2kE5V3U04Ffx
ETK86dt8mJRtmXfg+2THCmswBApq4TjzC3U+kmeJwFd2qbrh3Qxxe1Ua6bjrXps42glXpocs2EhT
sE5NQPESVxdtriKv9/cwdli/e5jxKIghcykYcLguSBgqcKchGwQuNUKnlzx+fgFbyUN0Zb+RmQES
M0oasc2EUGaYRac3Pz0dlCfIg1eXLe69Csl8D9lgroa1FoTR/S86/0mHT+yz1R3+yyMsoYbbybfd
vyywBWoVnhMMF91St8KDoyc1hDbNtueCaPOBle3ExPS4shbpme/EC4LN9hfqA9bjTWM7u2Unr3Q+
VjCSk30CXtojIku4FT8SLF2ycDaCttGCYoL0O+g8C3Aw3aAtO7d2N+FTNUpkGfCb9psEFQefJZgD
S970hjQ1s9ggLnMAYSletjJLKMtcS2pjchhQjTPNd9N/jUYKuUkBjQVZ1Bo0xWQeLouMNEAiFBMc
dYUnGW6Hw9CFUJ3awsfVSVXJg472Ti9YUOOOxog+syp5XCeq+duDs64dPdrCSr6VFwU9nHFJCL27
VL2uqsh59nkzY+0y8YiOm3AEQ7gh6GzMJ6tveDSARNBvy5hCDU/1bVPlJnWDG669pJBevpFhvsC/
TZGeK3eO7lqy448nFMZhXpDgdFwTyrg3nByX5Rxscaq10Wt+mopak7U7Wrs64ojN5KXvK/Svewuj
R9VLSwKJOk4NEeg3Ao+usdDykDFlZouz2CQooir0qeCQ2OvtLevgdxTwfDjJYgPm7/0s4Zhe7jo5
Oy03AvhxXEwxxGRltQzckTBFsv4A+fIFt2UX3nTuGhbay64+uN66Wx2Z1qw3D2FL+1DexJGngOdD
WnbYiGId7ri/YZqbDSw8un3fSmHPYwmFmPkjnqnsHgbXxFtSTRnIi0Pb9HmbJKIS4olOJaFmiNxM
OVdKeBoKtOAUjfbwzifAfg5OkosJ2Ter8SQOyIbhXg6a6CDvrWNUNGbRWOw/7fCzKEm1XCWJRzGi
lu81FwmDL3/OukG13wU+WCTGEPtzrCPPMCkxoLq2t96iiW4orR+yzW+sUgRSkC9Bs0UZGaaOo9CT
5BIXUX1s3pRzFdORtEvVYk/RGFFfmPWVy/xEKMiVvj4R0cjuft0ANPdmnYZaUXyC7XxqiZk+qGIX
5ySxQzsR5vNvQcWJ6bPfVkL11sDR6HXQ9pH16UZIuobzKa8q06+rl0uyfxYSkrV0rN/GJa5S6ApJ
pOB06c/kfKuDbO3mC/VUXgqRInkN6ZcWQbvB13b18BDUnMw8UZUZ4NmtWu6TjLMRilG/OAnhovqr
x6wuMfP3dFw1JNJuWZX0bCAgc3FLC9wbBxPCow0P6aCeM1wl80A+lG7ueF1MA3YsEwSL9KaQVsBo
1kpmOW9HyjoP06iIJwNjy9SKRvCIEtKWGwiIuy9Ugra5XTSngH/yWLuV+YinOHLFiIpfVYoXpQW4
7czJrqJT1v2zi8W8cHDrDtyg8W9hSSAQAhs0+QFWWUBySrKXMfb1k06K4+oxdYyW2lLucBDHTq2M
aBoxrXVPUAStDhpk0zeJnz07uPmTK9NBa/HMSkX22qt6GyEKUaZUXNZ7pCtAX4IbzUErAMezmrHz
FIpgJLuf3pp32A9d1OSHt+WNovxc6VuP9NeP+9r2OsI+fS25VZX94KYdKYFUEQAlf2MPCvWEnSn4
rAVNG4usD3HqmsoCUTXlqKLLtBuK2g06PL+K1OthZ+Sxa5aRXxmgk5BfLEwiTe+o7B/ltS9W+imD
gij8cXhvYAcEHbQzxZbE83CeANVfXG7Q1xPrUsG9nwXsDkNr4DbquLwoCr00psb9d4B2bPtN6SDH
BSgTmLBoE4GZxpeSq2zgXcFeFONgFZDsaUj8O7EZk2NKftKAp3hmRM8r3b7IxNoEaI1gYjsvR5fY
JUAVEdR3eytZQJjFfb5aoUgaqW+dQqovpDA6KZICxonmBFk7c76YWdF2JYXC+cAglqItdH1WnBJo
IJHlnNa4Bx2mp72rZNlVDnEw+ryhnSS5fvIhkdLMhR/AfUNHBdvo6FuCI8QVxd/9kU9Ck5KGXPvb
MIQpaWl2nRHXhJDmxZ+F2K6tm1PgbcF5te1ZdcmRJ2hAZcIY3V0eEay2kIsljuRMCpioiE3pE4GZ
dRqGyO/C7gLvbjemYZxnrfW41RBHAos+rKRf3pjsJ6SsriJDWpYyy/4JuQcZ6KgsRQBvAMidiZPN
GPDUw3RKUvb5UMaQ3RTIz45BhjmVVGAvDCVERSTa/1lvN3+Tk6DAmUmxsNnRm5Bva5xIcmkjAc0w
ooF7BA6hRr0qdHegbQZ0t47pvdN7IusITjhVLarVQReBIdgsgAOJGst2hR1G6mW3+A7t8b5kPSp4
KIjWlsy395oA4t2pgkf7AhZ2aCgsjhSzsjNj+GkvrMj0hrV1vgMapjGMiyGM5QOaN2N3qG8g+wf+
OptAeLBbH/NYNfy5hdL8LJYX+FJoJKCxlDcTiyHYCX+p0AmVwaSI4vxUnkHlJv9+wa+laF8oi9Lg
sYvXE+kdyXhXelmN9m0ZGsV7SQ9kq/aYPwNOnlqRo3ZHmEsi3YjTp7lyp87PfoCYW1giWfIi2+q5
awluY51Rqi4UpX8R4qmcWaF5CU0TxInKGiNg0vK5NEJAL1gDy7bTjQ5eArYLRFPX1usBly7shJgz
Jbl8VLsI0SQ22OaTnCZtsGxkUcMD4a0zzhPJws/zv68YcTzxxsa1v3a2nyzUlxOQw9QvY+MmO6Ni
Saj9UCpfWLvK+jIkA2o/fxOOa6q48pcp5nKeXhsrbyS4w2NwhHgwatoVs8sVoH0HqJ9liH3Un8xE
ZXk7koLEACqYVjFshx4rK3YdbSkBMCKovGRrAB20QPWyCoYxVPGj4Sgq3s5fpBN2mZ7A+xerNglA
3YhsnPt4g+1ruAKvV/psVY4HwINTzzVcb2+Brfsho2N0qZOCy1Eji7LxiqpXgEBNOiPKndeN+qD3
2580u0yHDrdEbdNLA//RWzIqdyFFW8Qcw+lfitzz7cBt1zaATBFvRNQQzJH8OYYxBD+JQ/ng5mbH
PT50KPBlEQodJ6hncWEv4sBzp4y2P1B6bixTxI9J8CiLPED5mZ8IyZqOqwZCTgF0Ax0UCHFEQsrx
opw0Cwu5CrUidsTsPzQz2MePla4v0PbMLCx5eHTeVXQK4gcwoR1xXYbBn3Xla9gDmvPQnC/BZo5E
cd//LtpnijgOHMMC5mDUb1DIt8iCeoYZ9VzrgWj1o8gYYdzkuKkLVDNOV+Zem8+Y6pcGXB0O2p73
i/61YYDerqfugcjiLWn+dNqnbEHsBmI5g7wSGpj5UyBnfVSeKysMAg8UaH8ezIYWUrNWZmpc54eC
Vqc0QIo+veH/3WObfO02IlR9XoJve/BqWx8cRss9XJA5ztiUk0ZBnEZO0ElhOpvodhuTLVU9i/DK
jOG8htTx3UgTpVM3/98nhNWbgJA71r9nhkJPCjYtA7PTyOftowk1ugsKOKS0yetn+avpcC3kJNjO
gayqErCIhL13fzJ+xU32LR4zulfBHzuCQ4sYl/ZQrkuynAo6+h9onehk36nysVgy0MUS9SIkQ5d/
qsJJHon3JbfM/fiUsxf+k0V+T3n9PWM4cY8SKr6RMF4Nmbx/uu7zPhP8fnCIUR2712zZaPt5ZThR
coZRWRRp+yz3MRp8jCv/uSJg30DH1IArSwBVk22BVBr2Qa3m8eIcsnBJEqcuICfShxyPWRTiHysv
qc1clRaj/EDAnYAlS+fpvloBZfpVhYu4JsdKoItn41PgxjcHdqu8jqRU/D6vQWzg/Rzv//Zxjo+E
lz2oOHmEXY1izCxZp7Ccwj/AEEKnFUqA8eNgX06mu3PiJcbkd72jfuoHb+drLdM8utC2tH87EvSh
FDlZ6KvqaPhqNbXMYqfe4oPQsIgBlItn0WFUvfBb/HfPThOwgG14KfqTYOROdE1rvK45mOpPLsbt
/IU9MitjLA3LZwXqeq8v1X5cZzo1clikk7fqESlRfiDUK3+gvuYwhvMmJiNWLLmupWb+Q+tkWMhU
KRC8cFxiDvTcUcYpNDKQdsDrHPNIKiCG5JQbtB9cqhooc/YBnWW/VKN2exqliIbl6z+lJeFWFFaq
BZ4Y1j+81hfyheqzX5BK5bDm3kmJTwQ+pZhuHrGk2kQmaYSDirvqDFJGCTg+J9bcF+rLSbkCcxYC
vNDNEa9WJsjGc5/BIkRacsrTciB7gzfv1wCAJzR5/IhY0s6cWFUOERdYzrAlADupgHHdYYIKy239
TwM3YQHJmOcB7kikqI7j7gzXdgZ1PiTkPrgtAcoT9NMM5uTB+INhviS+9+WqsI6CsmajY/6aikAw
jw4s8VAGL9gyP9EC+AE95EyFdy3lrrLyqnidpd9PYPZ93W7RG6ZOdPVbKpOTTfu7vDQLXXs3VqpK
QqpTfi4bYAiXVd6T/IPkXk2mStq2bRfTxWOQ6iFjgF5wWRxjpUJgEVLxBvx1/73C83OcYMdzIzhX
GNb3P30DgGVlfhOelezZr8vuEo+0l9r911NZ0MhvqovqatplICaQPYVpoGJvZ99QYjlJyF2tJ3ol
9PZ+GUDxEGCspYwOvLarewtFcWFe0FpMb345VBJlNaT55xGhk1id1p48ssKoGG7QB9QSANxqosZL
G22/QcxmDuQ/sheQuw2b1vvtEPnQSKxKUVUKzY+//pOA2BoUx2eCxqlMMh97D1Vce04eHZGjDSwc
aF1mmwuNoH4BJEMaAAsDxmtZj/49kcM1qo0iWtLNpGyXNSHhNw8VEfHF2bqfsKIq/ar/uUMT8uZU
ZxyL41qlB7eiVkH4G/KsXDS50EGZZUBmuKhkUtd8+lsLmx3CCVFH+CHQa6N+JaxagHXfawZn8mMk
lvmzf2uvBcV/xF+QG2l5imCcaXQRD3GJzQCwHYR41Gu1uThjQRLqLR4f2g9Uin9hN1mOSo2LGmic
WtIbdoCT6BTkv8BCyIqhRpqwnCO5KYwQaJOpFRCek5BBaKJJDJbH7/PL2/El3rInlvnCSD13eR8v
GsuiucM0O3cTnYsWPlzIHlQRH+GMsblipSvIThXQlSbxTwOQ1PO9sEmuMP/W3QwAqjsHhfz4iQYF
4QeNPYX42UGsm7UMEOF607Fo0UxoQJ8crw2I5xXinbK+rjKkd1NMissx5JPw1sndUE6USReOzU7e
8IDZPRSWRZKaWPVVhOQ5VkdtHITivfNqM18NH13TXsjO7Emdu/mm7VBNXOqjukKg6d7W1NyEn67M
vDQ3+LvVvEY7VF/ojYDONnxUgifulA0zTWOfwi7FkxApjyek28DxaVxEYZftyoMz7ka0kXEJ91VD
LQEbrrnsxIkDKovO7zCxJYD8QErUPFNr8/ReXA/odqBIBI71zffLtLhV28AV4sV2nTHu2Ae3vlK6
lYu6Aw63vetnP77pSwE+NQ4SFEUiclhR4lmTWc1LwZ2rvtjqs7reY72QTxb6/qO7CmjMUpnjUqrj
KLQXufO7zUXC4rHG9KD1XafVwcDoCJDPcS2H68hy0V/DfZ4YJ7lYA6/MKE6Qa1Y5X+jfrUs3Qukx
9yjO62yg2AVdfEUayGqPUMvAI8Cyo/YZTEyGCLyHjO8bPNraOb6zsSl4MeecfbWOScDvfl7uxxaf
6amWoiQmKXb2+eQBZkkztUY7Jw+VEDlaPfsBhQh+xFlOnkx+hM82V960cDzM1gFCfZCFoYAzb+nb
+CNaMIepsHvAGox2P3aCJnhZeA5LePjGPMlhswk1x8XnjLhRtWKireQ531Xbbb9CRNABBBoTlEpv
Y4ZW4Xu8JSRAHvc8j+myzl/37pX/+Tygtreh1fLiY6KQK/Xeye83eq6PpKZaxhkvMjWwYClMDdjc
LqbYfrVrQQa9XNKCQjE5V2mPy174P/Mnvg6r5eVwb5fKaB153U/nE+xZhNNPfkXby4+W1W4THX6+
Oq5DJGMLut9eyWOunYUdlOzSoli7Fh9oqFRRgFqC4VBvSpMCEcgNzHq7OZWx1CNwU6gxI6RjPFQW
NLsArgccQL2w5vDom28zyzd89GmkyMoC2fLn8/D+GmQ5ojquohL5u9IXKQz96YxQtA5f7f2464Gj
PJNo82Dte+5W0uguCg63hoZF0/wZjOuHwW8dfJ/3Tj2E1jgeyqqdaOUDYDCx1ORz34XZcEsl7dFs
Ot1mC5FukfgT41/86MC48eRSMFHyusJv+VhVTNzJH4B+4R/KjzAINboFmZRe5OW5o2rMsbW3a7ks
YRT+JadcHUlQf9vgwnyFJC0Mmxy+H13lNAY3SjX3CALFSqIfoJF9XxO+MBPz9DMIVJV1W0yLaLwf
sVUDSG3kAt+U+vim7SVXrU2YJ6v6Y8X5oXNZkP5EQiwdGVF7xAbNTU2m9vyGoIM8gatzP2YIGNVy
mb4YK2Szet1ycXBZOLLYcF9zZDkjVt5LYxyD7EtVBDvVSsxYWcwv0VnLuVxV84zyowkLwtPn1f2T
SwEqoSjqfsGLU51CNHPgz8PPLecZ8ZM9P4PmcwzVMJefIu87RO9jGmeXzVIzJMobsr+mSwEgCdOV
VFtnOerId0jNG+WSnWxZdK2T2CJh+xNBw18lxsSQCNYZWWzYlzggfP40l+fFOuUlTrrjeLjgv25L
n0G9lxQjqzQqqRq27BZ8zdEfBgE/2cIidijdlP4mMgX35BLIby6g7QY2vKhjCz7x9x6fE5InoSZw
zuBeZhjSWtp3nY/xX/2ffwxHnx6TuNzWuF8OGROw4TQxoAgCChXkgn6WzUWE+Bx5+ZoKdmQ/Tyk0
IeqvUBUUOr5klyVBpCqGahd0fodco7WC9SbcDRxEivxMLopSY2v/RtSex/HmMEVpSC/kY60EDZgn
3zBwdxvr6CZoE8T4UL+Ja0UU1fbmO/Y8YQXc4kQQuKYZC8b3sZ6AFH93dH2n9R9SiDb53mN7dAje
Py1DebAxPZtBY2xMUcAZHNPBoNgyqE8twYUWoU9eL9FwRFHwFEoKdENs0DCGjeFibRgi4yR1HwWq
m18RD1LapmzaoziQrAkLu96F4yn7riOsueZT0SgacbdGw15e5uLMeIxFRQKBFjG6styfo9o85wzc
ZPgropFk/jdPFXbvriT3SUt792sZZUaoTS4qLa9LV1wYBd1gRKtRUKF3x8c5WcZmnQWLhqHve+v0
qiGke51/0Ww7ppfLrQzstnUA6KrEz/6r9UKrS1c+cGSYlUWS5fxS9QZ+PkLqR9mDWu9y3pIKh9ev
WXesc4/0JiCyReqHXRvDtMdSVu+8oYJ45qFxtOsxfMcf+i5hfWOvnnYjh+bqr3QwgxFk68rF7YCi
mlLtgMfxqBDAW0mHoEOecUfkCXXBWgAn9pidXSfHzakWjsCioH7J3NGWZVOwyXx2v1XF4jlaQFCL
zGGIDM7m5qGjrZ42Ffxv8XtnOTjaZshTvUuHFWNKa/KPGqxN1KrhQBS+0zLh0ZJcNkdY49pUryO7
1NJ3z/xMpE0nb1OQUAKnj3uNQpSu+wUjvHsnWtlcZKVfNUGtyTfKdAYVH5XTWOvvqi0G6ys5HbOb
7I9wF2HUQHEHch94Tlknbz1BMgSQuetMS2XfgiMSkjohdEAcBVz/6p9wJUxXzU7XfhEyFYonpQyq
F+bZWwJbs44XiHULbtGWAAOAs+WhVVKOKR/791dUpEYMtDMgzia3SsyjNX4sZiEh4KZt3TATEfk+
5jap7zDi353CEdIEtU3KS/3YUlEaFUgmMS09AeoO/ROdMhojk1sfsvS2ojGOItH8FmknAlyeOgrm
53AoFGsfKaiRD6m0r0WqLJKidfTIk7blzZfGo5KpfV6vm4fluU6TOPl3lxatRaZvBVgWiO81kJ9Y
LOCx1H+4jRRmMRK9zWsxLpqGx9rK6iBu9YetB4oHCaGr3wnOCYlhjWgBk6SKCPNnNMnkUqrEodkb
oWMWLsjhwUCxKROXDnKtW2XPJM8xGLOuW2zanwM/VabS7YcQZisxnABNTZis40BszOGBe6HIggRN
aFb8aHo4I1ZZ1XcfYBbucfQdEfVltsLiuptJu8lwd5g4ktaTvFLibboABaxWQkDHsNKbitVxqsIq
qxW1q4lo5+JqNmM4c+pNVDHePtNUoRvV+zUFVpyp5Sxt7wHGKXfjXlgTaTnWjPg6V0GYu8MfcQu7
5+5+O/04WQaQLWb/8tF3LLBNoJB4USzpsYcurWjs1CXGaAQ9UASc2MH/p65ElAkmcvZvYcpbBU5H
RkWXmS6ZfO2mdzdDE/c55Po7sbxokCF+tkxWcgqVxTjdK3iQVMjYku7UMCzCFM3DKCU7V/2/VVcf
2AuVcAHmxkZFa6DDfxQBAZlcc7iBo3wGtMcOsshMzeUuhbEhgkiw6KA4FLRzzIMML83R03IRs5uV
TqMbqIFeHV3btKw5zNsKb3YQrzKsoBTkxSMsYJwksK2KCRHDsA4yXX15YpqVx/FtABfw8Ys2YR8/
m4RI9yz8gKzSAE+wDl0y+pygZGyprvytW9ZMtpQekm3AzO8baXPVb6rpZ10zMikQcr0d4NlyDGmH
s0ksJn5S5J0vcHAr/sUD29G3PgkAwEGMAyVSkBeCeggsVKcGZ8VZsPBrYRdqUKAcG92bMGDeTiXp
ip396GQ9eMBRE1Ohzr8m+Lilt8zxBgbLPh/mPqVR3pFAKRk3V+jJbhcwaK6keR3kUdLXVniOhl6A
qA2HXAsZ9/jk+d1Ce4FOJx1Qnf8rdm5bAYC6fFjyiWvCtymLLW/azwxkiN8tqeGuoDlTH2/Cnl6i
VDWiEX4W3LqFrXm/Pd+95LDBJTPREYaB8DpQfEcfUFityQHdlmT8o+tx9A8zP4ZQIKcnGT5DIUhV
ZwVXQ4+jwCOGN9EYiPIj/53kMzbTvFVhDFVE4NPzP/irJfuwJ1ilUx4X4gmaDzv+IWshXtt2a+t5
7ykCBhrdVbE7DxFcLiMmHG7OgUtyj06Vs0ekqDZDTvYkYVlAM7N/PCWYbRJzk2T+12hQlAWywaU4
Xd2tO+Ed5Ma9Zag71J45sWy3nqV22DIvHfvOVyMwrpmXEqq114U0lnv+T+g2jHzyYzDhL2XWRsU/
e4b6Gle76GNwtRpd3YNvpzLRfuPGOUPeNhHSIoY0G3CHFtqL1nVS23Q4fSiqmxXCUSpakQ1RKfpq
ic0L2rmqFqt7NA6GoViggsuNJ+BJC8iHQh4rRHlMnmnqCNETtbrh07gTqjxRGc6k1+1em8ASuvrX
2Ce/vsBYww/Hac/OfuIXL5U+81PRdacqucProQc13SorH0T21ktkXtozh1VjVoQdIAvAYQx0GDob
2uH40DGzmd2UoDlNzgjhls90hiDYKz9Gw9Rp/9tK5BlwmNrhFI43/eleJaGUdCUNZ5l62F8EvD7Y
ckdwDQqJ4keKFPmE0jFP7q7ZhIqDOv46eEz0IN0wDYOMEV+MC0nuutFVC78izGv9aDGzcdGgzubY
6KLFNB0k8n7wMx7oWNUmpFe/9D0wwUa5ubH8q13QeKlEYG8FCVFnBtOLesJBQBdilhahN5nhAIKZ
x2V6QrAem1uFHKAmwsa+kJHsoyVV3S9ff/x847R5uThI2AKV4bt83RdsVda6rKsMpYXUDZdenS51
X3o1g2RfOT+4kggft1AlZ+D5og34nwUwEmTZUCsryyaZpAgNx71auYplbkxJ70up99tJRFTyx8jz
ewaFDE2yi3OBp+XbcVpdFK5J5pO4R7eUrXLDipUvrXcfFn1frvLDdpCgp1MDEwIS5LW1omuzPdqC
ZVN6pCxJI3EWE5lCb9Eeh2qMLYUdfeGCU4/kIAeNthz3CpJtoO6jaJEqUsyOdEnqNLAts6um7n1b
1YTxSOhKKbqI2VSlnHCG/DB6gjhGy+vMc/mzJe1drz4afZCND8AoD10ZBPo2Bi4rJDG3+EsqGKSB
899xah2xR59b3rJ83o/sCsn8gGJ/QKm8H0oyoBPJLLrBMA1MStDhLEDvcYaCVwobBLLOCLq0F3mT
CaIAPgdXYSEbcDqRIKwPOzQsQT+dmnloOIY4D0D7qO1cLCuVSc96RL6gVXgFbm39JPvaIYcdFOhH
cLCoY28Y9hqr8PFR5Xyzf18c1OTaq+zJq2GMHz8cRVVuF6GlO0SoGBwUlOq4wK2St1fMVW5Wj3LG
cU8UzNEItcV7j1atbDqO4HZ7TYOyACiCfS6PtJibUf4bSF6YVkr1M7UqBx7vUIlgteVEiXCtymh1
5cK/0g/9QLd9l3Ul7dAcv9/X8Xe6mcGi4rhVhK826A/NVfirWBK1s8WpLkJs7qf6bYiuFt9C3pcF
yxaPz96mcAA9xP0gGpFBFPArW06lh+hyW2WbcWtSonEuFtRgN1eOz94euwt7ZjvSIO5HPIAlq+Ph
LMuZjzKo6TwYLq5c/RbQrXj58eCsKHUfB+fRFJj4Mu+XEQb6EfP5mr68txLrdPq1SoAWed4ctKSg
y3n2qW47yNero56bvgEHbGmGpaw9x8uG8e2EgYh5nJwRlS431YRJohI7tSRMmXHznCYP34zadw2c
tvdp7FB04mfmeEgIWaFOIE1Iy1yyBehxdIau9VN55J//oeosVE/wNqpypGvwmtMOHXOgnyh1gRyr
0vjXEJoYHg7vHH4A3n9bcSnFff48zJrTYKJunmGi7tBIcPtAOqBrcesm+dYtS+6UcZRbbn19W8J+
CkRE6ZP5rR9rRJHaPKsY/5/ePsZSreiQH0bi5WstMZTo7R5hKa6I0PRZXBc29WuMudyXEpt8Ke16
E2QGzNukGJmkevxpS6omYDRn1IOvay30MrXKKbFuPSooOWUT8VoPtWTyT3TIsorQ1Ru0357j/hYm
aNf6+29v82rm8PySfDLZgI+WDho/GD+1HVkzxd9NAP+Fb1a1PGHAAgYNnCTu9H1ZQ3IUWErFVNSs
hVgsuYaSXWN4TEQOOgIyLAD5wJaIhkHidfN0hZRN02pZrQmJYyXphJNJ5x2nyJZgKPgAG90bPlrM
VsHB8y3cS0Boo8SdM7AKICIxrDCiTykZKKOSkzOkO/7BVrm29kusyPAxh4FssCSuZstJR25U7g4j
oM6GHQ9MrVloV1tFIE1Hw+5gucGykzhB6GH19fB0aCFXyIlcwm4LX0LXX5qovDrzdbkzCFZhz3x3
ODRVkTGTKMLDcekPUvOUrIZeFpBISQuqCgmp4o+41wFHKBnSl1QGp4hZpDuESQLfCYwAgj3UTa6d
kxQS1wCXyqlrI0IUdMbugjj+bafB+aHwsDF30FOyNEybebNilSqSqsfuB8QG5eYkNsESHPOGhoyk
iFImDZYLAyiIHXgyvz1pPH+MW+Jtxw5Z6iZOqZx4FcEsuonK0lwul/9573Mpa5g5AhNqgiSj1FI2
mfSyX2Qml3sQrCd+aX5j2mpdMmYqD2a/+o0KQkFPAYtbIUyYIlTFPm92NLsE9gspFQ+efhOtTC4x
M7bBtjA5Doh2dLfrdKQk+BhskwkXs3qXdmDERirvihnerUyqNbiB2If+tpGKW7hKQHAocJPn0cWV
zg/PZ76O5DmPR1GMiaDUf1aELdxaiZgeEWj8w+du61dHYwRaTybMU0cHaGULs+bzLvpBpivgqrt1
VcJkGgEPeFs8UhLB36sBGY62GAfWeTYEAOJD77SeyXZQ+Ii4iZ8Irfs3jtsLnrfzqPQ97gkQZceC
bEEreeQDm9vNnGVkFkN5kuGN3iHMRx4hwmDZpqyBiux8KIV37MU+w2f8rnQIggsDo6v+MuRH6zKf
PVtBmzvqhicGRUSnAK5BR8JDkkzqtAhqkfujZDblcby8Oz2xON72Bx3us5hpRgNdNy+iv0ltgGYI
U9pi5066MakK8Z1WgUaAVZtN9qqlv8Wz2J/+4EUfOYzhMcLFYo4mpBSBAmXDWiHffB9VH4CBLLCY
HjAepF0Hzr8iTneCuAch6//nAGhfSdIlfIXWCqxvf/oGk73x5u6T/xGHljeOwvDrOrBxZw5Wiwk3
q5P+etuF0YrLrPwZIKDR41iEd8KXm5a3mgrtImdelsEGssvRauK68oBlH3VpEkubAHG1mu24eBdb
wdj9K+v7rA4QZ6+RWrQVql3BByOIVSH8FmzYB+Ia4VYCSGgX4Rg/ph9wlMNOuh4p+6+yDc9xBdgj
kKTX+ME5w7XNZa5TWTRtMnYARcK7n3/iJDAl2grGGL3cd1nl57oOBhFwOFWd1mGHp4b8ja+8XYZt
3Dw8gEORYOjH/8bXU2BkOxizbGy68AlKuT+BP41UVZxvgD5s8Dc1T3FYNr/N6KPCdr65XbFDmDQ4
BZlIcFw+HusngjxFby8kkxLRRtS85HYVW8y4Gq1bgjPvTAaYjit/xSj1dXnEgoMz5k7D6x1pqvjT
1mQVQ5emtrKx97T0m137mfsxQburb75Mqh/MPeSpHhro4SDjFwHE8gWl2e/pFPcPt3UZXEP6tMuR
xqeER+23HznltJwwBxFDQmZm+f7g1x4bqag3GV2vPLR99HuFTh6ppgwnDMKCNA75mkp5oHwZoRdn
08DUfMhl1BXnTj4UPNzjKbuHSmtq2z00kvpM7nWEQrlBwOSxDfFIqAbE8oX/GOowe6k7cIWTwtDL
hOBuvqsqsiUmj6wSrORd4o+9pQ8D9+jsoeEq1ku907SOup7HkUpZresvbbLIU+L7nP1MnawthXIk
GnA31ZqIsiPuDRWlCLLEa/M+r/sU5AnUwpxC1by5UGeRMoiItmMNtNIaZ8xOze2XB0fny/JgchKf
hzqvC696Z1WSp9bf9XUGhxUd58FHivrL0W4e8N2eHmvl4pQNXsuYchVFPsXjI8L0wXrXgr2lkl1l
HtxBV0Qsfn6TMktP0FMfB0YMuqod4UnjAR6yn0NRffqyo5I5QXg49uXBkCTTUJlCF9sYIamN8ZcC
7IHg0Zyjr6e8VpiMPJXS99WtB+JQv2KCbkT1BZNu2OTqDJCeAw4pNvPIC3HDncJAiSUN6enWS/BO
A0BCdHy1p8Sl9cLrcwTMVeW1PHe4XCe/h9+TopYDlLJTAej4rBTdg6mSdhAMK5+Yn5IxPf3XnuEi
WX0GQLUgMWEA8gIuD+RmEOnwsaNl01/Sdj56IoUJqsJGJFUFru20/wMj3o+laKrJirofNy2XOJsd
32Z3gPqxxh5GkOomO2d5fxqmMRFw2P7Q3XMrvU4AfyldfF5IDyd9Y95l2AvMtKBheh7UElfVjPKd
F7E4vrT4p6o++xvoOJ3gZdbo+i/qfHwMNo3/aMxbUEabyv7TwWvLP5/dd62t2/FNt/kzOJemem+3
NVcFxcn2qyv5FU9YSiEjRdFtbFhqj+DSaBOhUfoS5D/jRdnDJ88OJXn92CSfum/IbKsOiTTKXqEV
svMgBF4jG6pGVztSS1rQ77fqpVcQUl5HZ1U6fFy9u76B/BDBuX+nbjytUu2/7CAKSX/+wPWwGsHs
e4O1jyYjVmHpbmHcCcdiQ250xx3sLvO1YjE6EaVo6278Dqnmu7zfjTvUh9Q1oIWtpMV8oJVGy4fn
mejBRYhFiE+CMlvKC1cZn8J9n2eqmBU/UDT93c6nv/7boanovkqVKOo4jf7VvU8nkZjFh1W9p8Q+
H10W+xsAExoMYlIlND94XGQWDq/zFfupVdbHKXjRSqKtR6y2tmsA50l2p9tu4DxOnImHW7hBxM7x
/BTnIWCMolA/pWta7YKY37gZZtDbyxagq10Y6VvkqOXDAPwA+Y0WU/Iy+ZgDvf3yw/eFMqxIjGW+
U2s8+LtpZK45Nom/rh8BowvgyVPAbSdfWmcerkDyAaAY2Vt8/zdiY2fFffD5zCJiT1YdBfy/OSZm
mpw+yQk1OQmv3F+Ufkr36LYlADSuE0jKN2nMDyRQDonRwlnFchbSZRPlD3k0l8zwU8GN45II/4aU
GEmPEhXhTFXrkDnwmEkDTFYb8YDAalLiojD3j4Zw8dKNlEHu8/vENsbFFagFxEw1t/k4JC8AFnXi
H9SQxoq9yD8E9cryDV1NVu537IeoL1/U+gNNioVNgl6goz7VWjvj6pWTVFRYTkZ3uga+RJkLJecJ
PdZQ/7iQcLgxyDrC0IKID77Cd0ZAXiSZ+UmQUsbrrgfH6b5PFuU/YdMaAhsT+jzhkjRuukSYL+Xw
Qs+U2LIjblh40CFE66rEJtwfZFWV1v/lDewGFtzZ/pY2GPb1hRUPio1DCt1HQBV1iW9Wz4LaN6hA
ysRo7K7JGQF0g19mL1ROawjL69hTMt8yMXdRo2+FNADKl/o0fW/umc4mDcUS0PH/Aji+Nd5KnQNs
gB5sa9DOLMbwDku5/2A1C18hNpcXkAPatXxov1sDZ2FjIMx3hSbQqRKclZJl/I2qMobIB1t3z5sQ
52uBHOVPuXPBWZqTxb4hQ6ILPUrsr6ZnbqlKM77GtoRmzKw6HdjkPRFllSPSEY/WGXXoPGTgIcM8
+uakeO3apYiBh10p8tC0x5zaap92i0HGb5WaCB4iVbGmvt7i09DB7t3rqGRCdzkGO/+3epvP7C0f
S1KeztJp1hwdBlYP0oHHw5A/YKNajRYAt1mUzjnoj5xb2zCtjVP+bdtvVyspvCKpALk2K5VSE2T1
T11rk/yevvtdsEJKbmVvRGq9rYNAxe2Fxhb14m68fZq2uls3xdWUNgZRR/S/P7loMCvpyK5BUxZA
6/Y9tHIIzu1ct5mS+ZKzubmWl4eKgFfs7gBpNCtY7l2P9wI2VzESvFx9jsUuwxcYRifpfe7HeJz6
u7PZN7n7NK3Q96j6QBP0UWWcVFiAJeTnPxqkJd7cnAvACZQGERyYRwg0haod+EGLJiIllu/21F7d
xc05vrEjJdXJYxscVaSybuLFWKNf4ZZFZ/nuXa84xs0Iwj3fhzU3L67PLgdvzyRO8gS85ReBnH4R
fjt04lbucAp8ltxXwb7GcxlIkWqdN2GoFljB66R1jJgPBj4+zxtneNaqnIO8v+/hs0TaQcFj9C5Q
rWOPNZ+j7qdaa7qU9XxVXJmzmYaS13lxOpLtoshrSBnnQGyk7mtsKhCptwknx5hTo3FjJi822nQo
b+sRw+NvRiTwlo+2GXfMvUcdaH1Rxd4L6JgKrFcH4/EmOC6i315UJF4flM5kq65nEa0cJQZgHFha
/ISulu63L/fjIgdMbsFMy9R6uNpHc6x80FUwLVzwpGbQKWjB4f9MA6Vv120mdQTYykXfDgwKOxwN
ZwOjYAi5eQNJXUJ23n5VYu3hyJo2TMT809Dj0Ez/ed5Iw7lzNpNfe+QG/cnXrPVqdGIVkwwD32I5
+Sjz+frsSpDB3pRlBt+3YdQlz64P8/F+qAWvFjpVIekDJlKdWc+i1MwejjAtwbkWwLC0ULjBkDuw
4AxqAiZCwQ2hVoknvjtjYdKKuu9qQX15bghtZEw0LA4a7hn0+f9uJyghrFLj8dydagoMcjskBz6Q
kIhYA1Pkcz9RMXkX+lcCpIyw0T05Nh4FB4Eifdd65cBA16QZ5OeLwAI1NlGwmpxBX9pGCIuIvLhE
SsAzngHuqS7A7CQ6tXnYeor1bklNWJErV30b5bQzQPdEqm+/4/EgDfhXMLvgRN8LyUsOT9zx0esv
qE0AAiQm4dqq3pHI6/obZI12kSsUfYXDwNwgn/ulTL6OtrZhqwP9TkcI/LvP34Lw4JV9qorpWxsM
8OVMkdt4YQxf8ONjYOCJzix6oinP+Vwn8IJYcgIoa9L53wPXJk2QYIdKMDDnYntSAI0uZARLDSmH
P2XXYanys+n3ZhfiyuOtWZgV8jgXBMOZvissIOpijWsuXWx3HYZ73s5zcCHZZ1M+ngc8axIrcYr/
WEhGvbBRFgwSuUbFGpLyEFuVTHfGp1N7n2jM8B6vl05WCOf0c+ywT3ynUsdnJ8Al39wG94GDdKPb
KbdA6i6bED6tGaOaQ1YmmRsAfh6nY0Hj3JHcMkWIW7aQX9vOEeaojxrJx+QemHUL///rFIejXSQI
IPFQLqVK80kQz+qyw4Xq5YRJq1Zv/GtKCd8GuVfg5Jl86ags1NH1vjqQ6clkEfxe31iOgq+GK2Dn
kHXGbBVggVDdoR2+x2aA6jCmRHQoCF8u9YMNqHl8YkQ1aPW5fm6PCT0btwlZ6D+fN+unCTEi2hK/
2r28wItiqj86TGL5ZGGAuBv0Eex+O1x4Lvf5Bh6w7rgNFRNgsGFBCJ55rWi18cXbcZRezTW4SzD9
TbpVCfdw22JvKZNBnpVQZMtzi1waPAJliC7ZJLk78MW91UPQQ432qmqwciBGfmc+J2fQf1NBWXGx
BJEnLAxbOkBkHKcCwxJZnUmdZngjsAkwFqVmvM3GKnMEGG4ftYh+5DKMOoXd+cgyFTXrA1QIrDT8
zD77P3CC0ITEazZCuAQ1mEbwIdz1gw9rOm+Ce4A4E2EVHmkcKQBUpIujxenNJR1pXIiubzZ8KISF
gf5tGVWJU8Aq0Q/522BMsT0uGkI3SSbSAiXwOLa8ZDYfveQNP3RxgmMY3wZXQ+hKy91leXPYl6BG
mI07gpyCCQOBwGmDG3czk1EfGC+75DRbJTpgda6T1gZoFy9MTHsZvZ0uzVr+EbaUZPF0pCXxAGou
T1DRh/lv4LVjVJlpkouoYtujABSCivLBoWijlZsXYQJt0z8o00huyv18uGnkB5XftHA9Qkj47ORj
wUyHHMsYkzHNQq9EyCC4Qqa8VMM1lXpSxnFZ4KvrBZ1ocrqHpZPTFoPcpkwHrZsnLYvCMwBy15Hc
e050gyhGCCpcMDu6ZZVIvMG6HatwKodsnx2IrdBA4BPwCbK4BHXcLsJLeH5rJfhiWInoXBzRtfSi
PKkfEfPPinyHL6ZPI7+UnBBZ03aWiw/cHjeKJECBionF/4yHzcu0tXlGm/DISDRcq0zdbqSvwpOM
OGB4oEQFH9keBg4h4CmQwypjcF9ppduu0IVxFbCcuuHKpCqmJxSa31QHl+KM1F0z3SoGqi9Yy1bJ
T2xnn3SwpflEvLHI1mKd5J4J44xKwuaq1IgXaIzEZjnYw2BScy5OHxev2bLOfCTo9bUJ+RQd8FzF
OU7RMJJNndq/u2mUE5VxMQNQ4RYohwsKw8tbAzlTPHQaND/Hb2lbWGtT72sksxln4rb6LMdjq9C4
Wn28EHuCXSaCvcVnhquFbAqlOas7t7nSjojlBUmpCDrSPZe2WJmvWBFzUBWvD2SneJC2rt38yw1U
hEcOLYpGAqQcoupkZFoiJOmxW3GIvIUv1vUCdt9p1+fGXA+LLr3hR462TpLTqkeXbInv+HOzl8Wf
I0ONFw1R9mV3eiaA+kjLfCaZHLTdI4KpqVLf6dxqrpaBEzJcLT29vqqM1z5tvzRa3MDHbL7FVGlS
Vpp2whj30HRn4x7gZsCjbaKR6rxH7h4VE3w7i33Nl3ykYw8fKsQdLVO98cvwF/wSasl0xgKETrce
oojTw1a6NODhHKXpAcJkiXSuxshPhCqQZ2oFYF5MbMYuOKAnUFMn4lpzKdt2f3BEJtsdpg3GCurF
gKFMg3IZcnPht9VibPyFa7PC6zRPC9NCOrQaxOcZ5CFultN3Cvq56uEodVvkoQT5nkf+ddjoFqBZ
fjOWkhHhsIwSJWU77ErIiPH6WCOvZPwi2VTq2x5dJQdfcp0YbPy1sbdLG5CStLQTMom/cPgN8EuH
ASIptMPPu7ZvipmV6IlMyWKLO1AZHNoZdmGDx9zABlJaZe7f/RDmI1jGclVvAXl74HbycOpduAs2
nHTA6vK3e/1SD5pib2AcEYdXbsCOvrIZIky/5Q4bXP1mEkeBLEI+ow32J/NpyFUALXFP/cIm5btD
yhp3QqDd/FEO974KZV64xK97ZpS1Amf52lYO+YaibC5tF5UdEYR7fd2SaqTzRpUljTtsLsjbbg4e
pfRVcSFSM0oM118Zhvw9VO4P5aV/dJii2P+i7k/8K46eGkBC4K70cddjEUEzsF79YY1jqQtPMyT8
4yNpIR7VOpcYDWCpEBN2Z6Z6cn3HbfM3HOGHnwNrUb+DxZkw7GeTmN86YXOsfwEmiGFq8hVrqQBo
i/dFTwhpHOaquAH3OszjErWVh99Nr+B4MhlVBe8RI8vXCRgde1NspatZ+9g5DTynACd5ul272wHI
/G8yF6ML7+Ug6OM9o51JVoQ6fdD9T1kaAD2jmU7uA7/NT3eSoWHCpLJ1nNyqf7h6sAVIn87hUVhu
bvgDF+5JOAO83wxEmGT6dQPtH9KGAOM8+4z9scRkZB6tzdzBh1kTFDhluQHhv4UK3rzxLNUOeRYF
z1vG02xNhs0HNWfTgNLDip8eFOnFhmg0qFJqP/FzuYdkXXWmsKSiZwq77yTAJzQO19/3IiaYuftT
XNDwwMFuyV08+CvApvWR154gLjnHClhCqLddn72xctvJTM29bQJfTdLAA6T3VBUH7xTYiTXUZYoa
Qoe2KRJ02Q62+67huKYrQGeORNSzNcQA05HXgPctRgzp19a0heyaJF/H6wgz4Fp8oNZFO1g18OxA
dRGxwZpqRvwijPEFt4xzn4HRUUwom/yw6Uwog41V0mfl4UEoKY5X59T1D0Bxs67uYjk07Yn/ssfc
bv3d2IrCY1dxBUbOi2qsg9uLt6iJJQFX0mPfoPcO5Mz3BlovtFxC0F60FUqNTik0iXSeBu9pFugi
9HXX5i3xHpd3ZSEUSz/+7Bc1FQKrRRlPsLtGmLAmtW1Rz2DBmcmkrTF0q1jnExOViyj5FoGnwI/O
ZXbTHpmkSkEMghhVz7DoNIMXj1GgHNuoGjWB6JLlSq677WK5e/AETTgfDamoivRDKvnVN3l+5jpd
AlRN1ZsUyZvPhO1jO+STRGLRszsCXB/rCS274MHv6j80dcY5RWPmYpjXmnEs0lSh5mUFdtLpURuA
CWXydRi2E/WXMrXlAcK9vnBOV26c3bPNIVmJrUeVw6+viaZhyEZuRRzALfwTiQbUXYPLD8NnpMJ6
Uy8aqS6RaZVflQJ+VfFpWckmwLpxwtpPUNkwF7dI8lAFERjKYDW6KKtaU3D2RPus4nv6QqNhK5xW
dS+ecJ1r25T7fHL60DwlfJsTdPYyTRP0qwv0jk13OF2qT6LBvaaCz+BiWPrc/0JSrUDKqLET9ySI
tbp/89wv8SpMZTlfdHCdzK/oX5ZtrInA23aF9Xg2RpkfenmzP1UlsEJhyChY30poJq9Uq2FeHzbr
Os0ELA4qQcGy5QYBnCgeHYtU1R59LEE+0eM2P3AyBxNZDgWOtS7rLHbv7rjphDbfUzqobw5jlZxB
o/fe7GhMv3WBmDc3mW/oF/foD0NLQ/k4yc+ikgh2HDZjXAePfJIMFYuCZLibO2TzoFdeHsfI6vZP
8HinTN+5ghLeNQpy4PhnfZQwCAMQTGjv787buGYgfanvZJSzbxJlUTIUd/0tqOubnUkgzhOd9H8q
z5ZKnh8j/Epjm6R3eJVmOpC3Z1mm/MKULrHVo9VlxggUuK1HqnwKuMFYLMJ4dwXhhtxE05/czu2x
9eEMOAI0h/M3icn+pyI34Ggb4/xVYpVe3duz1QomTWWDBbsJyvUmBaOgQT2Tyc7B4ibFnDIAyA7M
eVrf7iovUZOyYQetgKre5S11sK+GZOekJReSMVzwME5lKcgvqssXwaK8YUDLxWCulmW/dEA48fvh
W7FsIKEPkjDPsCmmzrxODn5dYAjQPxSMsHwmmcjg+j+JwlRbsss0NKakb22wx6d9qjoYcBXH4vhy
EtSIhOtFt+JGluLyyYz4Se6TsJ63l9NGOoCivuL44gMyhetG+K3UQffEbvExtSMLDmRxSlypudXz
GZKYNFcaY1WaUzPb4sp3GdpxPz+EeCjgxk2b+Mr6NJ4+sQ4B1gw5buN56A27cDU4zPPMEEIiANMj
qNc74Pehv10TC8h9kl9XwCtFTi2e0cKMbCygdUdVkdV6Q2xQk/mnC1svedfWW+21c1axfYl4suYg
XGQb6NLtWQyG9chPfJJE8nuwl+acZywfVg1MwFbRqMt3slO6YUvoE7N9+/KvHlMm0kOfb+R1YWg1
KBlOhz6EBCKaWfZ5JwlvvqZLdsnXdFl2znTvy5vva7OR3elv496w5//aufgqMS3bFDHq5AkuoTqI
WyiJ91oK7B5FsCNa00A88UzYVzljKx9YV5352CPhk8JVqVwPq7m4PGYJW/ILJ0ZRceyc1BCrLM2n
+LfQGAzKI2HczcEIOSxG79HYUwtov/yT6OFpPMSGbWhC6FDrnPtsFr5EdUXcphr8HV1q8paTlRb6
iwe3yfF9Yq7ohqvNDPeRM9ox+z98gCCEicDnQvry7I8EcRRtCSfagDRXU247r0mTrGz+Z1eMyjJF
DSnQ9d0bve+AN0UxGPtpkPs+9meMVwIMg//4As1YT2RyJpUS3iEJfdeeoUOEapxYaMUojLjvcGdh
Q2Dv4HF50cldCEx6nvkKmMeLzZ3clsI08XJ47wcX8mzbnbB9jMzuw4TmaX4Gd6BvmqVTozwmFAdA
eKaJPZwKBHkEyyj1F3kuKRVwW73EXIe7gzSJbpFdZ1MAMaB7jyR52i8Gzft8MhgXHPk8dqn282x4
5rtMLtXh9gfDa8Sl2ElxOg6SlGeOIjoJoXfDHtpZSyZIBM4zOENR0Fsc2flslpvTEIUlf8vqoRag
LW3SMjf3BMe/OPR4PGLR813P16l7def7DmXGXgf1Idb8994IsTbS5s0gZ9n5WI5yJEpEi2N4K1jm
7ZhRjbpxVfzrrzsgD2ppoJmcqhMB4jh7jJ9nhi3jDowNCQQ2aJHbYP5qIYbcb3kmbjUBDAYQXjZf
wSW543FEbIlBun0LoUAHQTOUcVt6DAkCRDV/Bw/clydAva73gmOmeqLGn7NBpCkJGDScUS1RRNj5
A4xMPonjd0Ki8/yeDEabC3uKGWRStkHoMwfnaITVgjM3Hbsd/14bM7LpjLz4McjMifJHOCod4Vri
u0k/BXHw9LK5tbtszEK02sIgO8g/k5E7+fcIoiZfCbrWdSgTKZKhaPvRGa2AufJNzYrkJdMBSrRe
XLCVenfDeOANnzEb6zCiZlcZBfw6F1TC1ai0NwlXzf86mGDtDiy5Shv9N5A+Jlf4rKJr+NUGg4WT
iZn/XqPyjvxZybBRomvZfoMUZPG10Tc3Wm8o0ufMljj+NvV9a1Z6AKfJ6NhHBOkrzh0LsSo6HVlD
vHsb17VXT2KS7R7AQQt2tZIIk9R6C5vE2lc367CiOqhqLdzJO5j4eGyGuYDSJ0ox4NtDck+iNriX
SOY3DfYAc/huMg4Xy8Pflpk4acLmggJ06LkvDGheQlls0Gxqi1ZkGfB4VEQ41HM5P70u6/GbqoiT
cmv4/Bskzfy8OBoYHiQ0zyVqANVwMg/FuJhAlzUDi3Du9MOxMfQSJyioppbvcgDlsOkKmhyngugB
2LtuTICQr9cvF58k/shFYS+7zu+0JEmu2fgqsTxlkIkEBJdJXrSmyiQhRBi281ndkTJnxTE+0FMB
I3q/XJITodE5yS2vgc8eJkwuOnwckRCao4bh9hqNtBek0xTlgyO9ZZm6E4SUad5JyGxhZBjdsDbn
9jowf2g705nx5TbB/2Vnm13aVRoxSEyaiGCrumNCVviAT5d76Orq/NbE64mVVqLyMrpGoiYLtd1x
Nib/P8oRPXtcRY9Jma95QcqjBRR94B9aziD2lOXs9dBcaenYciwRXNUJsE4JD+e9rQLdggIGS4bB
bOjjQ7mZUB708tiWCSyaX8DmDg9iurLN93kmQeTF4Go1mUz+DUipZacd3nJrzwg8dDc9bYlgv05p
gQUoNHmcscSA2RbQifCGtHobAq9IbImTJfIfkV/PP2WqqW3YRPXmuDDUw0xQf0GSbkhocRp/B3dZ
k+GG/0Wzndg2YN25ce9T/e/Qs6IIlNAW9wuags8Ed5kP0gmF5pbKuMS9B+OVQNBROVHIFwwmTwCx
b/YmEOuvcmbuIAlorbwKN5tK5Epy5aSfkg6dfSXBTudybXIQaU4jMf271W4HeFqZeDB4BQa9xRIf
f/r9s1zrYVNUUZp+eJeac9FNkTbL4TP5+3e/pupWFEvFFGYx/bSy9rn7Uxz48fg/m1N+XCqetyiT
xqEotgfS4y9pYXJQkTduIPDx45ka22s6aAoXFds80c7kzQONM11PJHg/ifKw31EaQYZowwpOyDQL
ub8zuThTPxgD8X3Yg8VwapFrb5Sy3V47SiHQJ0yiZS+uXKPqw0nWKRmgQV+D6R4sGuCqiZo+U3IA
Og7mLcgnFu1RxjXBweHICbUzWdUi40kaptFPeeiqz1W9GNq2XcJkbD4YSf9q61fXAZkPvtWrWrVI
0k7IavVDqwcKKVoQK+DWOazqfP741zqnwRVVSGnGwpNa2ph+F8QyTsQY/2wErFmm4MSFvjlfCz12
sYZuTG7dkb6Czciy6Uxp93naPfVCmsDRxMwbZY0xHbOecY1e7m3izRe2i+vGbT/H5BC9LKMdUjBG
7TdFEHdBGSH/KqU45Eud6fR7oJ0t1ejBNiuOhmMIAkqnV7dOJsEy/JVwbkgaVKdpT/t2+CVivwkm
vL69NrPY7qEkqMoLcvD7/eGdbxvBt6lnNdVg8Kvgx74ajf2kFcZBvvDwsVCwPCOMt+0pvLsZsy44
+vHcrBikgpvKb9V+EMiR5V5NZhGlU7BOoy3VwvbQMDhI+ooglClRIcYEU/873UlmQwNzjO5a1M/M
MJB3dBvhkXQVocPnVxIR+SB+DOAYpfdJRcp5o5boL8V4SZU4fJ2AwWug4Kfej68yCG6lFsgU1C8W
Svi23GTtMpRbzG1BSjUyfG99oS0sXfNEDhavy/UIFx73/YgjvbugV3rrDWKMBqSU/WhflG8XBNY6
Ed5G/ZrtkH+oWsIVqwqRbPn1YFzkv/BuqkQ1skPgtSmQnwxeLuGe+Id3xABVgyulca0X+i5PQQi8
Pq54X+cdVGA7YxtQ0EwiVQ8bWvTtRx/2+VkxqEbxLTfKUMuUEXCrAkwcsIRi1EyDXK9waXq52aL4
c+Y+t1U3cbmZZpCXldq44K1NfJC3eTSAFEOHe98i5CxKC01PTBZFtNWlB/lRCJx7fYmb1an2e85I
vBDepMdU4z4gTDTcS202K2jnHA3jX/O7dTyPGC7lvEp9ZYWEtoTFJJMqmVxNflWY5RHZ6Ne5ZNyO
e/CpI2NY6XQ8OC/no3kXjR26m/B35mUR1wxxYnuzwf0dwZRaeoU79WqGOAD2WvWLt7CYwVt+DQgk
kjp5PiNDhjuiQlVA5rZDcLfaBcjYoA3vmYw0CiXdqkL3J2YNOcOv8RwJwf1SqISUUYA0G4jbYvkw
WhznAYuhvVQEJrs/H/buSJBlqkSeiRDvzkE4DA2iNGrZjq3QialVxWvRdQkExjtAimkXG2YA38vj
0jqejOFblPrsR4vX+oso1BT7r7+Xd63iANrW2+k11GkoUCJsJ+m9CRhtjaj5dG33dIoHS0bIL8I+
BKpruT7NS/ikocR7Ml0+dPU2rJi6eQLrv+AVSglUtkZn3IyzzI4lY/XbbsBYtJe1uYim4isJe2BD
fL9gPEHwWiYsjYzp9+p1ZpMtjMxBBXhwaYMtPoiQnrZtr29NIXM91PlFkOVbc3BfmdCVjecdFTW6
fqUEggQxmDkt4QMKJXosbYytKZtE48RIoHL0tRIQ2gAKHCkbLHpwEcMf3cdZ4Zi73QhFn9V0wpWu
2ubTF1HtdHh0+2GEkpFpwdQx/ekpBRw9JKwGoKvMYS9aOlz/ffRn21sPeygp0hh7OHY8zKBQvCmL
WTdp4dv9UrBUDm+6CgNDN1bGj4FaVqVsqrn7YeLjNExf7USHYhy9Ath1cbsMmqBCjfEbjAa1f1nv
0otIIGN69/NiGbx82ZJHSLaI+xpVRgdEp59k9krn8XoqiJZCAnkGraYsTRzNMr8o76y1JYP+eO/6
EH0xIvaf2uNveuRAnax2xptjm7iZlpSseKiYUwrPKx61pKhWWLsHDq2C8/LBqb+3sr7dUOYHAvFQ
c26R27YD4WNu+/pkerSp1HSRtdIc/2W7uizwMYHLSlicL7zL2Hzkhu83Yn8tve+zjNqyeLqDP3+k
WvpXorr0SD8qOdXFLN7l9/k7Ly0REq+47mLYoreyJ7LwxzkNALAxHg+5PXxuDpt5G+ZKBatXDH+b
BnzJBf18Dnk8lmOALjxc6JgLz8nkjLNmSYZIBETxGjHEgAUMWm5h0tz46b7Uk5Irv9pWaf57NdOu
9GKsFwL9sAGqxAjdTzie2cHzJMB8ryr4RIn5pE/DEsHPeug0/LVOvLXoAEmmAeKhM3AQZxBpEf+1
TW0hyUizqWq/l9C4OQU0rO4VBGOH1K/OVv4Ru8Djekzhy3c5BYIv+LlhUZWTvIoVUy3tZCV0+VMb
7LiFU3CbFYRXkWzW3fywa5xl0TBq3Iiq+upyDZ14XD7gvdYHONxrnd9nseXb5FxHjJPYd53WOKVf
rY05AHdrO26WofYBwLC22o1eDODAIPpW0focln4E9uILseoEyWA122ryfM6mRY94x4XLhkeKtX05
zUl1n1is84ZCQQGANGzo7iOgHTAJ/WTxy8pI1UxZ38s3RKKESmAUGbNesqkQM2K3AJC/IS1gIRfa
0IUU54X6BYgVyvH9RDu1dlaMfn26tjCembbqDNQlMOkpo3DA5S0xH8EDfM2QHt0MNDlVzNduDKdc
NEehoQreAAD0EnuWaOB6k+pU+/rYabM9InYXhasYWFTrCiBZpIOkqkwCHcVRvca+2McPSEnoJfub
ny/y1pCDa7akXLCOgJm4XItHXzhY8kC0XISDKABEMli5AxKQy+eiJzBT4JGp3yIW8vJjaRLNk2Ee
PjGzt91iHcLyLN0lgP5PqGaFvf7lvqNx172rcKZnyHDwarDF/xv8eZ4Bm0gqzauHSX4hWddk9JZc
CY6FM2DeOxHqWcrm7fjwI5eB/mdXU8khvd54FLtYh4pmqkcc7tW9v3cbvOaGO+Cw72hcBjDVHLMV
Z62XcW6POIOouofZD4GWLhbE5i+jvaX7rZgemqVX8fZ2bHVoZWpdQZWx518WZ1hEBovip7d3q52a
cLbBAEVKF9Ohw82VYIdT/6RVvOzPVMw3i4K02KXjhoSpf9ChcQZF1YJF0nZyFuf/S6m6VAOvv0bJ
HtCBzbNShbB8QJLYPy/lp+oYgle1T9EfGxniqSeDYj2KFULzK+Q8EbgUB94m9DpHYXL3iuC5lzje
U5BPJXNqusJ1N9U4UwuowZX5gNikFQsXhb2ZSloElQx/O5B23OXi8omgeLIPeDxyGm8iZNRK6pbx
rmCeT09WNfjzHxTAtGUSq/TS0k807vOMqZaDoTNTXl6s62grkHXf/boPyn1iqbqcYponmHLDiMkY
l1XxRpL9rB+iizXrpEoW9oFsl3fPNWwy6Jg5rIHKQpmkuh9PbyTARYmTDVZ7s1XRwfPUXAunFGSi
BjjbNSnE/iC5RhenIoYrc3HDUCHNB+DqtIep+ISMZC2VmW/3cmDNqxrbigpb/21vOcXZXfWFSNsQ
4rQwZimrDn/VMvb7c8L9giMgN7EFV4gex4T8ZpRtlOlIR2BtnZShWLmSuc8WD74BuCoK6lq+jf10
SF8ei1ukPC0dzaLSYI2Tnc+rdjM21uz+75TatW+byWZLKqBtsnSCaOQKmkXblkcPeiHeSFjFc3ba
6PGbNdxxfTjxOkfQG64NSzAMzBD8oVkVfoQSdBXiJYgv+Qx9CyGW5YoFmNwGnkgC1U21fzo52vhc
fpv0KzJdPmGWVsxIFiBxEYwNiQMPxGZHOnA/LJK5MFt+ef4/v6/E6hNzoonAtOS6Kzj5P6ap/KtG
83VnKbLJ57FvcAaXaIFFmiMVf1CJmDQdfiBzhy1BYHtD8OHdmZjL8JeOK9X3m9rstshA1TgleGra
kAZ3p8Y3B42GWfr5J5sxKxJNGwTB2k/+cFoJTNIh55RYWBYjPS9so+4uYZ69UNQDHTpb8aALLPyM
GLWyFESlZtd0Y7TRH9Sel/S9f/IVucJ1RC/i0B7SlX71leOTdVfQSiMW2rt5F+W+DDHIphc4rA4G
wKNN6L5OvBlQ1iiCVqZ7glFc2Ik7QxCixrOHtnRlvPdsdw9fZrkGvprrPO5g/qW3u3frRJOVTKeU
+pUrnwBuyzVaaUZIYxNQCCtxp8fGRPAakw2hQ0PI7Uqr9exUACW48zF89gx0BzAIuyOV+xz7IG/r
8K0eMIQm8K8B7rBJ+skcePQ/V03P4o4h9mn1NFzdVd7pFi8EDUQ0r5xO6NUF0rd4AYAZMovtH+Ly
5hbkAlkOmBSDkrLtX8Z8u/pe3JNKLEnbuvDgDpYsXefb4SiZezebCEQVUWeIexEchNI7H81srLY/
5+JcueZbmOUg8nandNY0oG74jlMWjrB2TS3tBFelvGsq0ndVJIGN9+1ASJ2DxD7GlS+G8sYEltdR
FUL3CeDLesMSfRIP36Dafh14PQdpuE9IbIe6aek8nypg630kxhB5TB02O7HRemC5ayvpCwYhtEJw
vE8JwyLK8akOXEIaGPffmMJc/dnPchuIkXX38FO9T5IbnoTqBPcG8ODCbvlGQww8jXpVVxwqJ9VX
hEYQyzqC3fC7LO6N9q4tQ9lj44I+WsHxzm06t2s0FEtCl/rUU6y+40ZrYAkgDMA/kDDEIwtd1U63
bCQCvTgAaQA/P3JbIsIGYwTPTr/VmfAgpi9Cv7VdJ2/JClzqzvPoUrzYTETBGN4XXv8SyI5UhlRW
/MuHiakdmh4OIdHGmX9rPcgulCDl4zyDpRvRL3n79GspWquuTXP9fbHOygMAK944OrS2gmCr+LBr
cEx3/cOoQ75oJRyh+lnyYo37y8L3fFQpRpSTgDzYxop8dgIo5UCwZHAVzIOtSKDG0bOdZFESRtGy
YHWXySs/OsTQ+XwRPBZJ4ZzrGML18TwVWiQnh1ocVVVgTbzFxgRnw+wC/PxWXKhRUyni27JXPNrj
vj9FamkR8lu/El4c+SahLWPCXf18niCy6zzXfNWCXjYD8smAZ9F+VxsdYDUjh3FaejfYBIzQq0uf
ffPd50Hoz7Iz8fSK/S8jZe2x11sSX8FEnVxM+6j8i+lw6qUH24BOo990qUQ+Wcjt/5U3s2iVidGe
KNywjVAbFn924FHtu0k5pNFPhcc0PKDXc90NvCpVEGPgK7su3IvDW+MCbuP44L2yv8Y/TSj/1RsS
BoOrQ7+7tPWf9Q7q7QnBM/WJXxbjsWgIAZGh1R1BjBDP3rJAQDWb0sOdmoXu/wbbhuFQbPDo+WjR
aKBFL0D8ufUq0s5Zd3iWGW39nukUswaLHkOYD28RUt1Zb1M/7HD2RK1X6fGvoEW3q2TAHqE7UDBq
FXJwK+ZwvfGZBKLFtRoR4oZeO89N8jdyp6w6KUGnYdPv3/OnYtwKjHrQPgDIhAqzZFOpMa45VxO2
edLv++E8PLGjUhb4FuvoBlj9UXbyeePGLvp+LEKNiq2djiizm+xHyuqU0WClJJOCl4CT3xvrO7bY
+XTlZBw5k0TbdZJR5zeJWer00VG49E/v/fN5p6DRjOHCrcAVQsXPYukQ2aQJ3dR5rUXfT1AxZxTw
HiVBPmUN6NmqR1FA4UwUxsd0CicbMVYiuiWIYnIp9YTDVR/mOQrtD6/IFry6UkqUJo01/OS5GTx2
Q8EnPyo8Y7HgPxL8hdzVhOlr2Tnt9AOy0DA/NmDxErxQr6uaeaa1DhR+8pYyCo3dMSaAejCOSpFr
rqlgEsoGOiU1UgAZsahoNPhvCbzo9n3mlfxjAM4kx/OEqAie+HorXyg2QG3ecNM1toXUAWcL8r7s
9cP7ncqmcs7pPT6q66kKpNPN1CwyqKwcTRELkAuqVnHGhOLKvvWPnCMGHvdVzZ9cInW6REE0S0OL
hkfYv8EsuAv3uAhRAoZk6o1AdkXJNAGQdYmidSXevJsSg82ht0GWR6Ckqn6k8DpBvRe3FZPzDUn1
rG2RIFkZkJBXjQDYI5mJ2hUevs7Z2yqZfr1JwU6dpIW8P8DNXghF+nOwISnVNzkRVBTxQpg73R3S
sUciDy281jeus9hUwBLPb4Tg5g8E7fnUUqO8WiOU6igBGY9a57p3CubV/oGSt4WJjYYw/84TtjI4
D+bbbqxZ83fI4N1zecozV1uvJT2j0CaoK9wigh0DJ7rbDbnCQCY8zhbim7oIpwO1EWEQhV7NoyXh
DA6QIMGeosdZgQlfG9loi+Xu0B0aUBq4A0IdRyTvkg8y61OAH1rq0I56MWW0mWAo4IadWL7Zzrxk
TUP3T8PbZ3L1OXvggrowa8pbu6sZXJN70gf2NfW/MPD3u59A8fVLUcGXEFEP1ZXaT3UVXrTa7qLD
wqXIs2nuHYZNTu88UJNryonNUuk1k3WlfaMrdCUXuAIJ8bUmZ8dqnZlPc5zWMBMbG4t6o5SbLEJO
IF+8a2Fh71UAyfuX2WOHfG3kxj95IqoLliNySQu4t1dOzS/hKi+E1dEF/lT6nmzflqJoZE7h42cn
yzT7+iV4mzRVxTaFhtRc3aqnszsZD2sY+Tcb4VyeeL26ZFiKgNxyNX4FXSaI060F5xP0Fk5ypMf4
R2UMC7fIOvl6rtP8j5MWgInwMdUJtwQ0YJPoWn468CyrD2fzGgC66+/NWlAWLXsasNdzwcfghqWR
tyOi5S+lp7b5eQ4mLpq1M/146fkCEImRjm0MNVllvSgO6dvTMjnYKqGPaVW0sjtyufz4zIT4AZOU
o5eaAjmh+WrAgcRHKjBzmOhqk51cgwrS9bSF1E/dpYBgYjKn31++LyN8oeERe8CUIQbrabEqwnPB
AGQipJ8c+qelmfmbNtjBagh/SzuooawYkJEBbXXCVXWmXpXiGt5gCSwr/ZoSAc5a7oTPidhyToSr
M5NuL8s6+7btXmnUusX9QgRYnHZUwQPTglRdjQrPFV0weX87NX6lIGNnPEfOIXjiZ+8xPqX9Cp2M
eWwp6fcK+SbSgoyeXDyUNrL7x/t91xFH0oS43OaFGrwW/m5ps5mSqaSeHvZwXAgZVq0AVbr1a8sX
50+44YEspByIw1+w7sKlbMxDNvoiE1gUU00zvdwzOzn4wD7FoVT99aBNK+ueefzCi6eCit1VNQn1
jWteo0dyx0zot1j1mjNgcn24tE8wfsMh5eYOyy/lI48je03KFUl2OpOPJPsCcUGD2Qp4NdFMsjlw
Fq+Vkh3bP3EX+QoocXe1ESKdbbACZPC5VlCgIsfBFBPoQSJWFr4Ku8kz7x1PoiNW99Zjtrlp6o6I
kxxTeHJBJiR+Hxao2k7ocBiMqd24nJ24Ow5hAQnIuKHDOtFXcbCERL2W+TJknqYq69CAWEGV1Lg9
Mcdg919Jyy3b49oZQEnsTnYK6TX2rXxROEzbMkW4z3D6+04BPP3s20cNe0r2Fx38lwWS5OBf30pm
JmXbOm3FUO/HO5MZp4OD3TCyn3xGNmvbbY2X3GJF7CzTMdIaG/dZchzaaDHAnMxUOEieXS4+J7+A
WmS/TiIohQm3BFJyj0494IOGLll+gl99Sn9Nt4Is+krjHaSy6NW/g0CG2BnmLODBRuKC/gL+lgQ/
6XUewVFjX8TlDcU27WUzu72ivYwf03NZz9NwCUu0ftq3sltcPll9Lcq/XvQJe303RZlGsJTHc+Bd
aApq4dGFiU2Ykn551af3sKVGP0X6oBvmcunhZWmv50VHDXeEaS7MaWwTf4mtC7doSdrIpNFzFBmL
uaJBPvhnkmLQzRjUB4VGbOtGQNo+7xrPC1+abFQw5FauOLS/e3BjLcCaaD2PAxD887DSaQiVc4/7
bAgp1F5EsNI23UTlWB5LvpZUr9yjAvXwGzF7bkWX28CJjFPscea9hPUbaCaJp4zw7g11bBOEKTaG
HakjkaC3Bo/xV7ArPkrlixDjiMbIfF3dju6jWMELJSIw6uh1nQPmcip4FxPNPp5Ykys12t72ac4F
BupebY6aGTlqwWR29R5U1PbtBB0cpQ9jWAx7GnGU55KmZWL0JkpPFNfbFqkECxCyTxvSrfkKbhY3
VwD/2aPWJeifV4TLw4oLa9/NzUR6+V2Ao26XlZJ5Ei2PzUGnYqURylFFkyf2DlMuFjeXkyM4QW4U
8q8mDQj2WE9WotgOC7NUKi667nTuXjEqKM2FP++HUeqnhdRnB9iS3thNiqmU3qf55XutRK0awguk
7ysiZvf00I1C2jVWmEoPuitOOPjZn1qsqBwcbR30HLS6Q4iSadSZPxE5HiJdHoCU/CqEc6JynXmo
yjAAw+eJV/6FhASqqePdTBm4gvYsaQ+zMD25A6IZOa1sDcWVCpmb1pw2w+08OkrGWMuosWkJXQvU
clHzNM5WTTY3fqnOZS8ABH0yL5m+p7Hmsp9mMfdK49dhtXrGe4/82MpNtwQZ5VCnRq0q/GqRlTag
x368T+k209BFo8HcpOHxbyG6IVABF48xhNv0FNyOhzA1YhpuhxXol+kRgzBfzpec9nET2SMcILve
ipEZas4wda6bEO9Iru5v2dNC8+LCurXYgEBJkcKCMgndmQ4dXiTMZmBVfZh4lRuWDUKOVAP6IhPK
5NZn3iGiLb7evYvFr0chuXcYAkQbJJBR7tf0iO+ImGwxd1BUGcdARBORDdNdgNlyDQe/9mqljCWV
tDkdZIIUbzvSPFmnWSRUEZVHw1P5cduBrMudiOBk7jyz2RkKa5FQPPj5jslrN+bisk4h2y1dQBl6
5khIBmWIo+6EC1vnKhWDVSZV/09CbRi3oSKYavrJsK1W6HioDkxkwwMxKscLM9mvEJyEUzZAJZm9
3ELqV5EN6SLadYR7lrspNIfDcMofKT7MHA3RWLg9540Yra5rR/LDhVMxW6xJ1G+R2RD2eUa0GbKv
y9pxoWjbS3OkLRRVXpGSZrloB2CXAnnBAgBKWk1c7NBP0SjwQace9XucXMs3biTN5xbGMUyaJ95T
f1Mfngn7IBPl4hu69cKd5CzsVAs7JlQPCip+HI5WRx6HTmVfTyBcnS3nKQuUX09Pnldh/7RSH+Fj
s2og59xzVQ+dbfRNcCqracT7f9SYVCTVtyEBrfEYxI5TipPX9LqOjyrZv03lEmdRgs+YYcI6l3dr
zTbyrPx3/9Qrx+b2faVaKGEDSS+TBwgnIJSnSYp709j1m9nHQIu3xzp7MYazgE5nahRCISrWMNam
PkhHQaXUR2A3iQUE7sF/N26OLDimq2rSgA0aj1g2QTC6jZNj3Qx3kLYY5qSQcRB7d3mlIm7Ym/+8
Qc82QVkSLtZMaKv/Myt7/b9aWqrWGSca43ynxHvsQcfOmjraMRvhc6TsUL3W1IlHylJcjN6jve9r
/ixepDt8eG59lF5qNrUVa/FhFw33O/U3bzKPcq8iGD3EKgqfuwffvMQjIht7ncrB6W5WOXQaBQeS
3GjVLBbEcnXbPBK1DMd9VgHv2ycaplt0ErFPKD4UtdCPHeYwBOVCBWVAnsCyYpckXUmhHcCLk9sL
u7rigNJ+vk2JA1Wi5lelQ60aw5a+3yoL7pJxrI+IzaYzI9Lcm/ZaEbLmScUVg4tecRVBnEksHRdF
elDoh/ojVz/DS201kIFlX1yeBk2/GC6GCgvsWkLTowV0C0e9JFX9eyzsUygKOfJyUC4HTzIhbZwu
GarVJEXaq4p/MEzEkpbyS9Chpvwo3G1ZDmvrAI5wjmG0SrbgTpWx1yNkVo6N4LPF4dzzDPtjKA58
GPiviPG4uO37w6Kxo3ejtRXmdzvnLWBFkxT1P2HeCHlxVTxw/Vy9eAYsZHMExcgfyUTImtTh+Hde
OcXWtJxni5gE7VeDPJ+aLdG86szDz4nt+o6dXBPg81HFPHVEU5WtrrjRYGDtZRUsSdRkftM1tvoZ
aYv8F79w7nQzEc80F5AnhGR7qsRAfOb3VYh7ft1745lRJ2vUyILlYjBkmq2/BqAgthZx795GMFN9
QQIbeDg0TKhWqVWKKEma+0XNobLveX695r/Qo2v4LwJKrf+tW3Tn4LvB+tB6ttXO0HNggRrEZ1qF
ale5j9shAHfZZjcatRvEn/4ocofeNuLe+gGz4iVPrfB4myq8gJ1yxiQPEnmijrY2w25gdYSn/hu2
CMSFOV6mv7uXs2D9ySB09H3hWuLyW5s7Oz+BKzplf71GbAU38ovYpVyuG6QYt38exthjhxZQdOY1
o2TcsTt62u6R/32JMV7UexF9yxhfs1RyQl6VsatmBSJcM2JSDw/BDhoAuj8iq1JAiaoXvtzeYR/5
FxRyJo5006UTP0XSnPtKEgKUlyk9VG3oopXRxFzKbbvXHcQb0sCOpMWrBULv/TSA1E0fJ8Gebbkq
/KaSMN9l/zxb5DtDGY69CUjbGI6rTaVPm2YZQPaJhgGnq1gXUU/Gr+2BvxXgfNre9ASiBEqE+Oue
jvScpqsyiD/oXKatyseoWXzPLCVsv8fWo2kuz1rduR2jIEJDdZGcHyBzDJiGO6Xw0diPJqUGomBi
RhZ2tjH/GzEoJKDhZ5cBHNGroHWo28a1k5ENl8i/4lPuVjt+VqTV9iwcIST3wnL3PgAll3Rnf/J7
Nvt/Ia9aGS7EE+3Qy+mg2D3RAkBGXXueRXLMbvN+1WNfLOMNuZk6M0QisYL+/Vgh9BehkXjMNbXS
AeahVMivo8unjoULOutKQR0lHsWYY66yXh/IGYdIVDV1fp3i/oDK8ZDi5+QZzKSgH3nYgr9spajR
867MWRkRwhcPOHv7kIoO/GMb6CG0N6YZswLqQ3hQf4mKpvtNIm5JD2QE0mB1cxaQzwjB6HXN5VSn
/P5Bweo+7zo5ti+1LOKm/Ey0fLmOKSYxuvbMJIAoojCwt6f0W2crKDw+ENJC9NrqtM2dVZyugtT9
u+gvTmkSLP8OEzQHxTY3ucoQGsd3fWPhRrdqQ3q0Qc0V3YSl0eHfHzcyRsPIUwVjcoWjCwMCGGRd
tQimnAvivIrvAr7U5KqCo6kNR30zYYsTvZ4Zc56pCVLWsFFbmTV6eikjw7wonA5PYR9ih771PRin
TqoZYEf9lB8oecAMQ115xZiiL8tpv6VT8sXJ/DBTGU5zuR5P/rjNvRxyK+qqHKXroa47mwFx1Snr
2dS5wqc+XLBIQ8kte5q26Owv14LMVYKMJF56Ui9N0QxeI64LBAXfuvDj4LvCi0YtCfTF4VOCR/qf
xjrfpvqiu5uRUA4MgEObNeklZlYE7PCf2Q1N4NUQJqpKBG9TzOA6ev5TZIW9y6MGFQb4BSR88C1c
Bt1R5kBHPHdH6zOzleVue9v8at1dFwwtS4qRuLs00/AMacIngTr97X1+FK/3Wed2ck8I1fg0HpV8
1Bj7yJ99Wgi88GCJLHq4AfpldPlxfHjCQ0ievUZF7C0PYkUtjhtjFV2rhKaCygjpHKBUL99+Lrnt
h0ANOiMekYyNTCIBB+UdY85gBfASmfhIq03G6NVT1iKrYW+oMMLAvvcEGvWPOmHNlcN3hTCKM+1G
lL9ybQS0jgLz4XLC/pQyob/GQDMG5A1oh9wT20wSvcwe+U37D+e8rY7OEshqQKHTKQ0NMC1nWRwM
Yi+nMaHEbJrUU8oSTU4FMFYeUHJDPkRhlQ1x/mMzlh7tBbgHxUlEjeYnkGtMFmbR959XyDlB2tA6
LqmfYIb7/NL+TaB7oy1fO/2RivxxlIprscCHAy3s/ibApHFzgD4Za2bpZF4tDWgOtgUJaiw90gvZ
rD07nzQklPei3Z+c4XKXn1MFxTagx7xzbUX65e2OxH8B2thcNtQ0NpEE/jCNgGW8M2aCkZ+O28rE
BSvuJLYQiCO7YeYgxbO1jdfmjo+ukGA20Crc2V6NM5GGM5Y2YdCbULUabOppsw/AfnDOzEoJIu3N
SZDjhy1ML2GJm20/eokH6mIPTmCU0dWgQ1mM8BE2JVv3R01HI0SLpdtE6m73c7Zi+h045YHk0GpA
xdvbWqPmNii60SAS1bhp3ozKgZHpqa9IaVplUJnA6xJUkLM2pi1sHnGwKA5nqvkKs0z56+MjfEsm
v76do0DTO8SDEM5ICzDhJT+wf0XOh4VB8qlsSKN8melfSojE3vP6OurzPUFpEW30EpWu8HbDKy6d
Ar1UBC/JsL3Jncc7l4iEiG9ti1nyphrFKwKR0IqzbgnN+eKso0e/hnlAJyb08V5lHuJh3h1fYUf1
H4oe2y/kR/3LJ4kaPkObHM4P6a1DisY5RFRSi8QU1kdiJRTpYSnHIvJjXAR/AdQGjWwkRb0nNCtc
66wKEt7iXpS927s2QiG96BexumDECoG+dLuvu979cLHh0OGwSiel4UfwG/C/SNOT0jUmLhBIinMd
Y6EnPN9d5ByGN4LtrUMHHsJ+ifQ6Iap2wo6ZvjaDY0Oc4UIZuAaVCjxnCkRgScQZUDEQFvGA8Hsp
pO+vsK9f8m/ktKTos0DtSfbBGyoLw/B0GmfN50cG2yzvCR8z+EcgHZ61GbxUZtkMkpQSJFJY/tYN
dZWnN3GkvZNAh/IzB016PMe7Yk7NSeE6/z3Cu5KWlA28uL8EnzovzO1NdG7tSZIZTdXuYlycbilT
ZGq7DioCEv5+I0xG6CnSr/XkEqxeqO0LcUKyBeeGF2L6fRMTHRjGPa47I/+646nvsZixvXl8izJE
a4xHU8L5ZXZbJ0OLzOwIgOmfrMftA36v3OP30ubW8V8cdjRTUFVHhuJasFNTSLCjUtj1+/bjX+g8
uAod/0CddK89vAsVGAQEd0ftHJlO9mHBHXpcg4Vg36t1Ud0Lh1Zugy9aElUY2mH3Js+T/g8PiWyU
dNQOl8DPOiCWEaeGS5fsV0+UYC9+9EnIFY6z9kbY7fw/AJxpfTNJ42B+EUutS7ULBYkHTP0MYE1b
1HTRjcE18y14DdSgEKrPIf3/VZIR7HTPkM4y/LjpUajnY20CV3PZJpogQSK8OuP4dXnM7ks2muNp
9pEb+iSxPiSK7NkyS/cv0vZAAMQC0CdYTwBZUCwQbeQ++OLbysmLlAQkNO8yiDkj4RP+X+7Qwwup
kYERZCcZ7Y83PCWmD0ao1XKKPN0OhUVHA2BQCaW8Rrff3VGG0aKqtSeuGONV7u9wWBl/GPwFx8oe
CF1UD/YcRB+9kKJFDNDt0GQGOvow2k11ULxJn8A1pg0eDlcR5LYbso3UWxQ63ZC0MnIx0W5eguJw
pajHk+5AR1ZCtQvCH/f8jOaqChJGOhs5A3aaG4n4Bf6vB5nOtOOyUPaJ9fupxy60ROSvbcZ/zP1d
qZI6EJmWXPe9b0824q0+PVS2HLEKGPh8e6Vv87VfArjJEsNykucdjtbXw2dhuMcEEsjIMgdMon3v
fgSk82toLaT7xv/NbrNkgHZDEGsAluMjhoDDJ/IidxjFQsLmnzxaq12BZcb6HdH+fKnBlKgnjLWn
4E4nQpLd3XzSWVuNfpkfU+FS6w6CYpdQnJSUXxaj9KDQmZt9yKYJ25VHSDIM/fipYSjGM5PXJRYl
9nSLrV86SJIhyzCB8+fWwHn9u617ze9mfy5EZEdR1NG0M6hNzUpX2kx8dUBZ+yvNhx8alkTLdgk5
+f76oZRySYkJPbfLDi3Dl6S/xBau+XbMIdYsKFQNu3SLval/IgLBc+JOdBbCyd6McJy6XZC2aX1L
JoZIjy1KPKqCwzihL1qASnwc4MMvzhBtrQ+IBBIGncFgrowCyFDfCm2NVELrlhpkk7Xu6iNOvRPk
rgvw7Ms5AkpcO/JuOSt+OKmqlY+9yPWtGbtdCotSV1Ij9uJwbcoHZeBUU2qqO0cKCneJi5CIN2FS
gjIXyvPhUqYjvqwFOx/KLuLBx21BjAmGb+8lKCKG5TUmWzVevSXfCZSTmq1jCWEolxFzFoLccq7X
gXUu3SMDWk7lfY/fYxv0OxMMR4qoqAGu8VwwGwEHrj+0bRNlbcFoNkmNTbDfJ5PbRAcqkLMs7g6v
l6Y9a2MTyZh8mvz+i++2rbmuyb7257NbgyX2lSrNHqYP8r3d5lPCfk3dMib+fkM4o0xwdADeflun
u0Pk7PHg+ndUzOumIHsOuXLQmp7nhhFitsInjHWtsnSX6Ct29VMMTAIUbjQCjCKWgB6tZwAoaqjW
D/SIvoOK+avtrCfm6kg65JoctgLTju41lPbgInBZtgkqUmJPb702EN2pu1hVitI5hm7etIckb3Ad
7N3ccnfLXPBRbJ8LqsDtvvE4+9VYVvEStL2GdEzFL8+WItmBYDnadn7N12b6BEOg82cA02iLhC7E
ewFQwNdkSx7HBuV0VyzUc7rOV7OxVtCV3Ndoucr1ifXLT3YParykYJer5PyilaVMbuzCyF6Zl46k
qP63CRzD7ZtmwHj8HLU2e03qWS/WckxzA6R2qV8oRY29/+KhyYTNhx8LsEFVw4Q8wjg/q0IRePH5
lY8ee6fHCgpuW9qIOTFc3Qss6cJTRflcx/cTvZYgpy75/YIcHRD9Baq5DK/xX79Mea9zD/+NuAGa
3iJSR1xvHlYADwk4u/XxK0DJLGqFUUZQaoZo0VYwkijxmSkZ4t5BB/29ZKpCmoRzfzsnG4iyDFho
QM/fd1tEWtkgBUBNT1UliLUh1rw813NDEclFOlW+SCizU81nTlaOOKGS0Crf60d1I7V8EG/VtVEC
nUh507zMKdm6vuZ0YdQuTqgknMgYsL535rZJFf8szx1t80bkTq+lr3AJVluqrg/TD6lT3c7fXCLq
7xFGr3tpQU3gwyegW5Ctu9oBqNRKgJshEEvFvDJTV1SUP21iY3gVBI84QS+IGval7xSiifgQX7Qy
z2u3y+wah+Aeicu/4CriRe4Z4naOOEd+UV16hDDA97DeJto0DygGywCHP7PBFLGHiHBwZ/O7DOpP
7iJkEysZoBaqmBP+fwic8i7kn36QchUMDp4Gls6Ref5/ryLNoA37SB3/oC0yY/Xxq6859x+aGNBG
+CP/1L1rkd9NOqXXlPUhkdbysJl7IHhTt5XSVnIBG3ZJAqQKbI9Vni5ifE1BiRTM5HX9xQu+UlBk
0OPC6CmmjET1KTVXjF3C6PorBTziJJj04OH+sMRFf8mbOE1bNtu/mne0s+afXudfByOWHmeT+aWt
oHZrpYa6tFqQFzPwei7VCz+LORhRjeHLAz2YVGv6L6EuuPI4CaKRNallokJ5aQpwydaKmaD9dCLW
cP8DCnkelYJ5/47XGxoVaDutIaTG0Rpd5Ajj1L4uq4yBg3eq8kEViXdNuxYZXsPlw1JKDwsvFU+y
G44O9jZNLXk3vheqrYa30xnOwtGJEeyCAGqMzObiJs/Ezo1UyD3KW9eVBwFywTnfha0/7uwmLfIW
frPYK7nQV4KgePXxXdijs5NTEbH26lSoYXxneHax4GUbOsC0Lr4ltGuCvDiCWqjGekjhoaj1q7GI
uOOnGCYv8IATtaAjNFbdknTXnmk9mMEXnW9z1r5lE2cVhNa4nSCAhLs89OvlWxCnC6Nwwca4iHrt
C5hplPpQC+b8c01GWYgM7WFY3tEpIPeVfz6QOMhgXqjXO9RUw9Mo8aFNErYmYgvSzItmYsLiasq7
vlxaNT49KpluPUEM4gNrL2kKrypS6UY8LLLhsPDRbglHcleFqSEBZQXp0k59fN44BaecvlSTB+jE
QMVYF4VTymzP5FdmJOvymjJ+OLr41zojLe2lvmg32aQ0uzbBK05VlDv+kBDk5/x0Z+RHAUPjZJBO
HzcRJeRLltPGcAmk88Cx9PymUzwKJY9rgwAvISG9XZacz3tSfm67KQLIQLeBZsg5IyA7MFQU72EJ
vt8GDuHL+AajnsLWOyE2YBxBpqF102eL8gnBCilS3NUx1ictAjdmzudlaaRACc9IYOMozyhk23io
9isVYQkeUIGxW/Lzn+mN+8phFUH3xkZ7sCepgr8aQdil7bsG9rCoytziysx735+Ry5VMJKxlEIW0
sh75rJOqdG3lUsguRM3GYyqWghDKyTQBHh9iZWBzCgUqgpKQkwOR9fvki173EMMFuvjkVVfKZfWQ
zzzqAqWLdh9AVKvQkPhkNiwsixGEzyGmbY2Kaor4yzy/RokujMf/FYFKLUT1xWIaXYJZ8YTWUwEH
jUgaQqRg981BHjqiTyTGz0VEy8el4cRcUmU/Quxbi1hX2QNCNMFHjtWtpg2682uRkQrotzxCIBLJ
vtrFSdrfxynA/5idekiNjw9V14uS9k5ZFtUALi7R6Z42DFlqLxoe3cuOB/wS4LM3rlHTvIl4N5Hn
2ZevqESybkPY0u335brD9mhs0TUSBnM/nsavKQ25J18gbH0DaraslDTJZMvBY9vh0TF7WEbsIZOQ
rZgIjl7xtzId1iS74EcVvLP3QkZ9pBLSSfn1FrXmvLpMAz7062KYLD1YyuoAFsI6Xf2alIyR7Mk4
yul8GP6pB59bHTTSmO+GvBsuaiu8SizbezD29t8B/Kv/YGMh3/qkJVEH/p+/zzt51bKADdriYTSn
Wan79T/N2zqK8aQfFBO7GfuAXIPHmlRIw4DnpNzFqN5yAHDuLgkwPr1LR+PaSKDj1ffLFJuw5cTK
p5AoVi38KGnUPPilV4BMSN03e5TN9fSVBqO2+uzuVASB7+zeAOXxzNBfMssnI9tsPmkwr3lZPmyl
YvMriUaArB0A3MwwGCmVmLo09tp72NG9w3JxtHLqe+5W4wlfkWIUMrwrxdq17lbbzbSZeVp2d/DI
dLorIgBCaE+/ZD4Y28HQ3IgjJZbHx5aEeVnOMpeeqw6FCK7C28/6ERqwuX6NV8CDyRj2EO9zmVlj
dS8M2X9f7w+GRxi5vnm4ye+HtaCnOMyH+j28Yuq0gR57l2tlC04yg8tLZoVeWwNVhm7MFNdmC34/
oZHtIuh78FSvzDlWLoFBhpsW5o1YOZjoSr0W5zeFzDgGeYsNNNP/SisxtA9bZ9gbKEchnT3Yssk9
1m0UBJ4HM2Vthrp2mduWL65+mdo294g9Ozd5v77RMSSOn2BVRcQypu/LIt5kpmQLCqhuYknnJEyW
jT4CKSypKLWa28VIItZIRae0I1NjN+nJyqtvlEpSv1aDtf6H2pwPmZzdaM45dVE0K0s3cCDVgQuZ
QhWuPR2bySHxfVtx1xP/69++Icfaku3tes1h/jbnFOchM9YOY8Ia3BzZOQ+MHNgoTsbkaanEsHWm
2aAjT1M02rZZ9UL9/KQS3acxigeezCFHLmvC7+2AFhKXLQnm351NPnN4gg4r8rgH7n5hl/BktMp3
2JkM7t0acH72KQ7nEPsGcsHel0l6t6n799rVZfSxJHCMXXlJpyYKXBenq0txPyd5cTdBu3cyCxUt
Lwnhzp9apyN+aFBA4L6yssy6CYzRN/ObIZq6GqCRIbDLL9vLPKOwJM6j4+0nEu07oaJCTn5nT/3a
bIfNcb3ThBqIvOLoGbIKO8Y3R7ChWoDxRZaRun2iaNKY5hwDkihNqxu4GbM5HCjOQv7QPhf8IDxs
If9nDGsFN3HNpfR8P69VMCd54/49lrHlNcxBOXo8sbjBTyGUZCkrt1HtKvPvkpG12xsfkAAUakA1
bouUF4cO1Y4Pnbf9lDSNWYuahF6Kd+T9hPTByOHeiuGhDeOIyNGUAgMObtVMGB1tSypMSYF2kBNS
jrYcxRU3yrUEvAOW1ZR8Xa4rGyFjd+xwrR5R0UD/PJKhshO5u7ojfB2IsgGqLDrs9bdZYdeU4dIC
B8nIs+tUiDSfleTn39uh5NOVLOI3YlXtevGoidT2mnfZQw6DE/1VmOma9ZVUT6V4dqCKPmDET2pF
3aozuV8pSl8cSe81P3Eelu0pIZrCy2NY2QIrHevGFyWSvFo3DgONWg7gyn7umI5m1DjrCSd0oCuq
7//OYaYdJ01UGRQ54x1UylHeW8U+7et6/2u4emCy2R5XGXypLm4/g19RkZjOmUJf+2fDtMqkTxR6
FvKpMepCvjqFu4gKWIi6WGFJKdSiitH11W/mn9JJN0W73DOLhy08uaGUqcMC/yuvH5Y4HPZiKkDi
xnNeAI5t9djYUGG0MXjEdrdapYVaJXl76ghiSPejcnQnBCs5Qxk4gN/Ht6F1sv+1181GrV4FRRED
h+yVsIdxwBRmuVe8oCOoUOQE4YQFjT4LN5AWodAgZOLOOh2K/32dZnaGNr6DGbRBO0dF+04r0RaX
zJ+lkQQQKs9fLXTB8OyzKB6hbyjglLgyIlOSf2uXBSpC2/3KHJhIq0tZnt/9gUc+Z6Om2l8itelJ
P57tF5Z1YAPLDz2wGvC0LGtAl8mtwdrYz3n9YgaDIZtf2mEaRDpF9QZgwxcxwMZm/dDVrOh1iqKU
tuPTwFLxuOVsui0lDXJ7CGrtwNpVacId7MFe2A3NZ9ABd/GzzpSHWUi6c8waTEc37EqZ9biNKwY1
qsCLFKmgVo7h98+Nciwzq9igrBbZEocoyA187Z4zHKHzPAN1Gb7Llj5CkpJEie10MBLF2O3MgCNu
IQoOVEQLGX3R1qT0lQnk86ueOn66xcKI5130yVAu1kDDxPPIFxlSt6QasoK0Hdb0QbYne5S/5a8f
lrIWshOaq2c4J/4jtT2hB3jH74YKS8pKuhpjoSEui9SAtXEzZ8ol6VtY97GVzTbrN9MBB7X04g87
qh9dTdtqprsFISpz90ORXbqKiw8gDnAwZogYy12Moytf4d3MlKfhSZl4jnGpCVGhMg3Zg3ehpADf
3JtTGU+hbbX6OUOq5TfGteSCwXmPT/sXomuBzVLw+qUAH/GQ8L/UZjcBFxCggK24ut/wXWMmgJPw
JmmORMyE4zaDe3OvG1HNTTiw7ILBynGD8jIrHactm6A9XlFQI0VSy57Qc9jZEUjVUfvfxmcTFiE6
7rJxD1kmCF90IkKrSYjwAzBBF1MDapikAHHSyEZ//CFALYHdFFa95rIsyQViVN7Ww453V42yEUyP
8O06xoGE5iTSNknWA7KCP05kFodVGDdqrMCTZQP+Z/pDxf0Cjzp4RiWUfC6p5KJ4jIc7MgAXRemS
hqBT4ym8azb3B5Hs8Kts6ozT8/M3Z5tNlb/eXAnlZY7V/ZbLMOt5fCzKXKGiHlK++m7Unp60hPgR
K1dk9YmmNnB0tawYAQWxugtiRUsvyMDKxE5+dpeO4q1pVr5j9p4ydZfS18iPH8TnFAwz5/oCCFfL
F/mQQhDsZc2VXuJDRGcsfkMvx3bJHFqv1CEzqwQGUfCJ/FXmMCLihOMdKD0DCvc9kirEfzRlDT36
NG5X64PbTDfhQ2yzKyi3VRuAHfqfk63cXVtM0GTzD3lNLXtIpXXZQ2eCU+3wwBBcVICq/+V83xKy
gI09efpfL7m5FHaLQly89XhsVhLoycygPaaqU/q+mMM/HtZJ63TYh7O5f0T+HJyxxyZoP6TX6ZTG
Z0nrg8nbf5Ip7s15dDYxIMkQWB9kOex9h/kqiO50DQS2BFm7w+qqESX1XYX8dY6gGcgq/DEJa15P
3XOwrQYAzNjFLgzRwDCGlA69v9HlRCvp6TkCwxWpl5vC5Ug5H7RuMJ2DRUMNgF9bfC8nykUgNRWY
Zzd48AlU9Q4zK+jlEXgg8frIFEPlKEJlQgR2Rusbik2UimPs/P6fX4GUldMGoRVWRoFbCqPQ3MAh
pkiCnER9KQa88T8BSeeJc0fXundVLrFGF33zEF+PFae9B4IhpLtgMtajp3LnszIXHL+YfHTD9gJK
+StlsT6V6Zpb7SOtM9hxLwgeDg6T9c7Nh169VHBNDxT7fSqUNhvMm8SVi47wGQMth+3IFhzUh55q
JOsuCPkd6X20jx/jqxs6fzbRr8qBwOGcCxxjrZSmq66VWbVAe98Hj0Fm1uddSFY9xk2JBbezYeyW
1hXxESM15Ir+Qh31OdpT+Bb5qqKUkOji2rGhh8l+jbBG3PwZKb8q+BYzPgzQMEduGYHlXKUOer9r
0kNtvJFTXbrwEg3gwSQK2Ek8Jm6gF19DB6ZkwYI84Z6pyrxHNhdBQsaTXX6g0Tw5zYsT9FV2QD6w
t8oAm+Q8KgsEHRnlHZrO78RaXRBeAvSU7MT6LGeAbpwUrafBE6qyqLEAJQByepdGiZlfImdDkZp8
D3SOLAAT8kJq1ODh+Br5hmgR3AzG4uNe4oyD+xBi/VXKcI1btWlGB9Tp5eeZQT9/My32pnXKl50v
q6O/iR1XB6e1egd4DnP6TWgISztGQ8WIEFqEbKk3UQf8JdiZ1aanSaihJ4ltALL/3BCKwMLXkhHV
QxfZKzWEJkTCCmx47g5p6cgh6YpHDLPeQMkfB7BqXxut5QsaFBH5rKQsFRItqbXe6BBcZ/tYYup1
ikvTPUC58vB87GNVFNE9Rbgt6fh1B9taBvFrQnDTn7AawlJ0M1mH2Be6+bJDjvc1ExmWH37wqKnq
u4sN9UQNQ5Gyk9GOLlGY+Cc8PLGhq6+tTLW2gkSeg/VCiHpzqZkcpGhyIE9kaQl4J01CXZjgRTvW
7KMeamiGDSIhyYO8NfeRmuF0uepAoDbaNKd6AWRwEKB8AG/aVSK/Sk2RLpa9OA7ASlcEJ3c+lu12
SQs/JRiYMKCobWafYMfTZZjkgluJ0lqB6jlxxEOi/ddIC6DgA6UoKNQcehjRc3r3CGo/lUe6KmoJ
THUMaNA50eZxn+LsCB48J6IFXu+nhz0tGQbrRNRWA/vgqLaZG+090quU0JFBEmXsErJ+36Cfyw4m
tZb6bPtksP5E9S72s3dn8CMeVDOJg5iAfspEDWTQVb2Sxj5OgspNN2vI+v8ChA2h0YLTzxRaHrnm
/0g+Rkd/XFy8O0cUNN1Xd+aOxKyfzluifWrSErLYECmGeqFmHUSeJScLlay8sUg6IyVZ+W1iQPz/
FeS74iEU3jInstCzV0EX3tjVWRllrW6FvFqn+cUVON2ISx0YtoyhEZbWaMKlEua4UVeiS46VNo86
1tFLrBpuxTI5XuHnGZalvI2CBcPLpdXgotrc2LlN7ULNUgvKuBNThW4hHn05VMANMp0Rv/ir+TDk
EJt8Hpir95eUZHHJr0rN2iAkiw/JTqpM1Ows9p01tMZYNFrU2FaornczcRTgBqwyHpNOjO4RFMhp
1ZqvnwRBjlMSCmUh57AQu+GSXlR2G23DC5zc1NUaD3TAjsSewSTS9IbGf3i0PWI28KZfR3lnLEgc
vQxF8o3tDz6lNpdbRnAYgyYW0ZVk1v0kxy2Uo+jfI9CgDH5iELCHO8OAgbWWH9xKkd8rdwzoPtIr
BZNhBqF2ONX9y/L+zm0uuhrEBVScQlIHrSzskbHSoZVJ+5Fe+cBK3ysZtNWsQw6QiL+/YryS5lx3
49Rzm0lzjPLEeLqzgzJOEeS5ZB+Ii9nd+RkIgNrEYW12qfV48aabDG3LYTMXflL7bC/tHDQva+2v
YfKymru57ke8SxfWqG6N1GeEzbqqBh7mo9ZS+05uWmDGuSTORgbymc4DvQHKAWpuT4S9r1bzRVDN
CJk9FWwFsIbmFxr8T5HJ7t++rBPNySn+lU2qk8hJ+Hl+yVO/u3arecqYQ2ksPsbFnRNPCV/9Q5b2
pPAdsTZ5B3ay1Vk9phoazkFKPXiBLC8BexTkUIFfxauBmMPLKU2zg39Vs8Q1iw15fCBNJ5tfiMXO
+DpihLc42ZBZ6kDBAOiDyfUdd6WMWwBiw9YDKoC3JgTipgf1gOS5ORwjRDBT7cLTqwlpomnHnCT1
50mQk4/j6zCrB91nozD6Pf3injllJNuCLjkkKCuE+jah88fYe+OLp2TogTLU4ekXu+KxoImJsFee
QRLD/6RyThv6XIKihe2Zk0EJa+9CfXrPcuJj0KR/a1uou9KSMSaiJr8AEZK3r0di/bpTvcUMZihz
yDODRfqsMhk4v1T8sjd6M7FAKqChWLF0ewMsoSvH1Gw12ZWFG/iHhdbWGhHj3BoZaFTPs+XrzBRv
wHv6LC0o/j/ssgvDHbB41919R4gSRIyEHJVTyu4IGuDpo7OaSZua2h0jTnngznRhaUhIkPnunH+M
NVtSvPDpNPLSQYh7c6C5+1pxqG5/MsAssE7zF9EVkEHNn7dY0HiAm+WfHa6Y+/Aj9vWrLYtTvJFn
eedqgZrbHeuSuQ64zGKNCK/QuMW4ql8The+XQOXMWAiRs06vWwOfLC9REr683qXAZqwKmZyLtDf0
lafdexPVAChTJpHe4p5WmbpL0ByzHQzNNlpzPV4TzSvGMUysGdmefqDoiq7jqa3E/eta/a9gEYu5
lAFkKB73RScmnknKYVAys2NEzj38WQgKR+Ryg72bVB2mI2NTh3N6u8uKLKfNxKf2hKPmmS9Yb/lc
7Rw7PBSX6UKfONPgaDWIkRtP90vbuUNggAKOEQI27Gs3SAThTqLlsAXzhCOvrf+qMA4kG9EHEhGb
qg5iDrInwRaBHN0jmTvAUGeehzaRFXldO7Eb/douhzSf6ewQcKBPIeVWghHqklkNlmibLZvuV0Eb
TA1D6q6uAvtJM9tYUFCYZooZvkN5E991T5N740zxx+SBOoV6fVNNLeMuAO+xiKZxVxTkeaNsjt/Y
vE3wQHyT0bJMMdhZGWFRilBJYvqLxXNJBiQUAYZSuxLe7o7MUJPUAQk5D3ADoMfIwZvX9R83pM03
sU8LfbfU2jUdCekRYrnh0cF3mc0rjaY5sLZ4JAqF6hAk9KYbdIIAESsOPBb7LUogx8HvZiH3df0/
KWoYDP4k0ZQ1xX6y6V/DYjN3Go07Z0PdLCP2tkaPndz1ozFiT0CjPLbjcYxzEr5AWLjz0rHb3MDo
/6PNKaWwhRnjuZEcys1PLfBhczGDbSqPftbXESB1i5/PJjMGpo0H8+gJkjSSZgRtkN1Dws+1O010
Jfa0Lx3JK5lKFpmAZhPvnKOclFxRw/7H30F0swA2hDJa+AA2QFv9ywQivv5QvhIa+tjJox1M7fvB
it+LqVgvLn4ve21QHThpeuLhKZ3photVRh9xtWMmSKvHMyER0jMHNV+RDEYXn3g4EbtTRZSDtQrt
w4oHu81z+dsLkrW96EInoiiZOokoqt8+mV+SyfOoTX1xY6ijneIJJ7C/a21+P/c+m3sHEJCUXaR6
MkfmYzGME1TQdiWyXAeWSiAjIiIRCw+8te48iDPzj1h4xdYH7Q8B/nDKKPz4+EmetRXToG2c7KbG
XJ257W39XD7mRchQkmGCwvH1TS3oNUkBDF9WbmSqM/IXqJlHy+xjrKzDpY0kXjTkNS9szAzI9bE3
Zqeq8ctbUetcD/zR7S1mRtYlAP/ynlixH/OyZweq8f26ANzI3/xZlUblrbly8uHZjiT5MJz8gx60
hXiHO0VjOVhgMDLK5KHKwKKnanRr+HrGM3bd/k5YQgVODdHipQnpX5dmykPmAc3NgeXmxvZAlzXq
dG7LoMz3DDLa9RQlXfW1a5lIcy3AOJmYaNwl5sm1PhRgfxn/Rs+mabWxW9nO6ZleWB40tO/nuURn
m60YMSQjHZtZ/lae9PyJb8I9RejjB2RrIlo8ynx18WSsoS4JldcA07Kwf0G0lLuq3qUyADnKpUHt
+5AjmYk8UB541bveA/PYnJW5G47WSYn75YMt4mintyEfNkrLC877ozAw4Dkd73k5YEyJzffqrmmV
Ks/0yqc+dsRGu/dk442v4SlEEQo3GiMVjqMx4RrG+xbJN8DDkSuDzp3U0tSDOHMXPsJbduqD6PQu
n9oSzNd3f8AdB+pG38uBnpD6NyB8SuUt6SPbu2MU2dERmNmLRTdkpRcFuLtlqWsk3mSAPct6YDEb
5XkQDnL0VikFq9DY45yYVuoYg7QtVIjBXwTUn0U3cvmxAqoma5ggYSYQmYLfYBw6jY6RQYyI/gae
Fk4pngN+b1CPAi1loGnxpJxbIizYIpMkWIHZXMbJRgsMX59aN44Jn9WaaQ6VTN4k8NvtGCQ4Ej8k
L75OJwNPkTiavAwwWIhfB6vdzK+T7MNW8aZATfuNQuIuKwmWKEf4efaGtrdMVvUOCmlIPwQ8DmuZ
s8z6N6gPahFgHsMYIprgDLT22w0AtG9Zjjx1zm3555X/qimpyHk54QE99shEi9mpU2oaWdzTbwTa
V0dfCFaDp68b0rJgkmM5pHSs47zxOrJD1I+cXm+HCxkP0DfwPOF+X1+ppeU51wY9wUOYk/1ZpjU4
qIovNubVhCZKR4fAxW+TIZjGlGu1sXFzYoolKnca6UEAByHENpOxLMLCym4nwFx9X4L+WhT+QzIz
H/aoRj6QnilUTAICcK0hKhlOrBluAJJNJM6xZWDBa80FSLIz/SPgnX6IRQJW3lfwcgCSemCQA3JQ
kukslD9g27YtCOFZzKrLkGcaK0E4DxcD6xd38Ja63QiGGr9h6BKoSqzRQz/g3rWV+K5JzaRm64wC
KvX2k4Zieb/UmknFkbKcCouBeF6Xeva7yyEsYBdhfHrh9uGX4gru56Y/gcFuru9effgYfaU4xO1K
TwIl8Cl5dCtZqCTp+9l8cxcRGuMJWSx8/O1mG3hdx29m4jSWGqQSztVp8yqIZcuKkN8IJ/Fxp30j
XATz/UDjzb342zjwKyqDIQUBJtVs3xn6x0v+nAVsWCQl5zXUAf5CHfklJnjIUMaq+Fqk6EFbm03f
J7Yx3+u2LDfepNZCauGsyrhZk/5gaelA/uZGyoflnyfY+Qn33w6LqrjYYv6ioWKea+qGypuAFH65
hbB9ULmuATC3rVKps75ZB5cG/APMoZGa5F7ecOMcjUAqpHeM9lbQjQC/+6z2ydHRvkov+F4/Y5ZV
GexwFaGlWJcZWzss+tfGmrpDk8RXv/t5KHkfUo3snVEvNxUcq3kqrR5hfwIOZ3DCunTFoSnBc7z7
Q3vycMCYx4fT8AOIf1gflgcQeQJgGN+rWH3gtTK5T9JCqtvUnm7Kq1JnH6fmuH1ry61v3ijto2Lv
8knpLv+/nsDnODkSjtKnV3XPFMFSPdi9yJr4R40snVhIYzHR60qWIF/bM0uZoUPtzyCb7zjRQJD9
1wX+1MPhCG3wUpX74nepZM0dbQq8fzOxIMdlNLL1r/xtnzMZftcGbrCIi6bNmSj3sbcsknIS2LSm
Z2lkns0tGNuBnsdpMsJnff6Yx6r4+Z2bQ+OLAfOZENRuWrPRt6yd8m9fZj2ACZyn7QOiWN9ofYT0
9LLS38hkdZYGYbYRLe0JtjJJrLwO397bU+8zZzsPMAao1b0BgF5dHgLHoivQC4xm3OxgqdUnsoRi
9M/iMzvC83qEAd2daQEb+IQeku47lxRnKr6xP22FIveqfThe4iyQz0Csnu51YkRj9dhjn9SC5xBg
hd2ZQPy90EdRhC7yWJ/Xh1jdjtOr4A76a2qf6DWJAnngGuxkWOdr1EZT+gizJQcEubZn2nu8uRXx
AZDdvdY8g72N1J9ksSjTnFR334zgGWrKtbtV2U00qeerSif+KcTq7f5uTUYbW3syz2YyXeqvgD1V
wY+uzEWJkUcIVD9E1RmDWmoBlu1jhZaPNErcL7512wMrgDV+i+XK7mbt0ghum55wToGNWUQaioBm
YIqbAkVYrzAGGx3Z6Y3QxbPvIufTdLZj3e+YK35uFqn4faLlEPwkj3rKfQcaTWx7pYrOWTqQUJxI
Nn4jL1pe7/LSfs0bw9OifAabeeli+4tPX6IH49j0AgXWY2ATSIB/4PS2EgrsPi1cqYM2o6G0oGVP
bEagbZj2By0p6gz/vwKBInwLfHTcakGdstd6b96zUnUDU48GIMwhXhPZf8gB2XHb2oShEiPXLgjw
8bX5/XH3F++k6BZXU3O3NKXxl4tIjJlWa1Hb7VTjZMDp0Ql8xYqZ2eBbbnkGNRn/IiOe1w/8D83a
2RXJGLuS60mWnQ8YsOWn80fkaHBTcAN2Nx1BaffOSmQzJp86r/Wdnn+YFSoaqG1oGrhy9AAkLPgf
LgB/YdLnivcxfd+i9WiKLyphQUuy5zDZIQDlZ7p7hX8vcKQKJlB7CznRXfWjAvV2dtoWr2GtnZhi
trE5N9h6sB6HIRmlrHC00Bwj1Sj8WxAbzNLFkvo1xquWBUYc/6ZV++zYbC80JsMZ/TpvHzsTZMwH
8cH10yq+EUAVtrPDxFtR1xIJ9TJ8pm+TNqymjKEPQiIYqCMRhlAV/eYQMjY+m/yitogfm5kId8Vh
TxxcHFZvJvQworT5QzLQpJY5SohlyXsHVlDLVFeKPmXyBRIFoXnCsCuE4dCfTfWKpcfPwm6hcvzv
ja7EbuKfrHwDjN2ZZLth4aRbmn0MCjZG5J1XFQXA7xvJbzyO72jHJgSaJRHfhr1Bj05cVW3T6t67
uZXaLtpSt8hO1lGudzoeO8VWrKvpr5VdSasq08Mf9lDUSA5WkeMc0sYqzNO74AhWy52PNTJjksOC
27HGfIa8uZPXOV8BEKTT6FQNNsOcoPQhfWccPaZbOeSzRJmwf5LumuVqOurP+ytX1Vqd5Cm9wVfW
h/Z/KsmhlcUdNDmReV//KLoAzU3CA+tZ90/a+CEpLszFMIITPRMcOfjtRwxW4CGxQfMZjV8p/VZl
eDNPq27XeBCPt69ChQi9ofNu0foJ+G99SlaCqLLuLN7yq2TuONN737WrrtxaALht8gnUz2CPMgj7
bUHCSpVKV9E5XtjJMoRVQJ52Wt6EFOOCpLW2ZcpKlIDhFGTHFZcNT6YKWLtIbEJ39PxPZ0A1vhSR
+eSL0wlaubDD43zhMkxvhXr0if12lx3CiZ5sbfZ4vBkjJAYwc6SzwkXp7TDT1ud5o3hdWsA0Q1i1
SkEXY2Uw0DURissSUEp6eFYCFq6EtiPO16+uUeJ6DdFB6undVhZMWGZnfgT0hv6xJ8v87CSYUr8d
3mfKVF4sIbew08dEogyh34nkdhsmLsPHls4eRbNyxfXvqSfZ0uTqzwIPo8d/u5bI20Ro1yx8NpW8
Z/AlKEg/D8qYjlsIaG25pINuG3D1jWQXgIEsNNA/kHFvNUTGkZsTTreRLW5PcgFQwiTvEEiFOJ6Z
fEXg7stgdZcx+K7Lr2dZMgNSaFU3jJ7C3RNLPXI6f1ZwIUAATr6WJ9wzFK5TOTJmrHPjBefJozJ2
zSDG1eEO0cR57aplAzvOBLeFEP9qqtIai+UhaWDjkZSbdz30jkfCxumF+QcTdPgsWoZlZHSAwH2o
K113F18Too6OchMfZESwepW0K2wD6+MRZkUtHD2j1FxQR2BuX3mTAZ8mEx7Af6LqEolrzyv/wqhE
MDI3ygYSbnvrFwOwNyfNvjRaQV4aHFe1xrPivhmqjCcrmQ0MdBKPQRSi+KIEqqF1YZoMf7XOOcEV
4gsiEhgisyFGoj+rd+tSEAuhwUn28wclZGSmJ5kyzJQ+g/Rh7ZYhvhqlgAMvvvnbqvziiIo/o1lD
IJO2UJIo5zCcuwFx5EeidqhT6InFfpPWoEaZBCQZIloV3ba0g+CiHqXBuDhzESP9sQTKfPr7tTB4
t+c+uKtliV6lD7UVlXhlj6MLlza84TJuOKPgNX9BC4DA4data1B87OEqNH/tCam9pCVfoPbTIRXK
weqgrOkm61/0B/F++kRE0OEbJKcPlSU4ULyGAOw3KP/kkiVuUpKwVY27iPeojgzuRvHufH3FaiHd
4kP/1DGOLM7H3/sU4c2Nsh7YLDacyHaYPcMjlXnjvUhdlX2ukkmZeuEa5Xr4b8JxYTB4BnotM4q6
nOoEUrweHZFOcsLxOiOHb7hdCcDNnS5qXdU+UgNzZ5mFbff0V/IbLgmq6v5IfaVSQS+8vxMOitf5
KoP+jHmO87dJ1PP7sTU/DbJoROUf48lDkL7WtE2Rl9YdlCgFvMFPQ3v1tCOuLH4ehrDkvF7q+nqI
zON7P3LGggnUCV7GR9ipxd5htb2LJkUvpMo7HZynfTReLcs30srAwMttnq3qCH9wUtVMnEceuvaZ
SA3Xue4Go6Ep0CsrvzPo4Qv3a5o/88fRRx1w3D+Ynik0rtTGN6nb4oCKCpWMegNQimClXfQVTBrg
KyVGpO13IRg5lJcLexXE40O4SqaL7MCMs6G59C11uA1TuDmZa+EumNmL6hJt2JOBdRmeIHEUJixg
w4dAfhfknlDpUgw/KPpo5ALd9Qeyc/FiQ58FnOai8KRNHFp8RMBPiBNAM9tbOCoNP27GlMD2mG2t
AZoNvVehKdPca1yxeoryY8E/IVTbHPdU2hQE9e9pI8qyb6d6IIbzi83I3TzRzKN94J3obvA3+Tbp
pfzuvlIUNX6bfEOYELDUBsD0TT89PL9IVZ9AtloO8cV8OyI37/4ojxoBaWaLjGfRfP8FS4XmW+qn
cixF4bXc1g0lGQBSmGVtdNNR8rvdkAb3Qs2I/FfbEbXZ96y5O89AxF9w+9NbHX0Cawf0oKSk+8BU
YevQxDYUfZ/H9YE+N9oT1NeK/QtXX09QBNgm+VzwUoz8MyVQt8W5w5yolW+bn33boUawcBpgHjvQ
oZZTm7NaMNdUSM52rRO6ILK0lj4naJqfTpQzSz6iPOU/Uq54EJhuNMIRx+IR8XjQYo43hIRzrmZf
ARp/b3joQVcDesLrfbaWAuNObaw+prizMe+G78pFiX5Nxa0wOxeafEo7VAkPuv2+ZOAXJBH583Od
08pP/sDPeV8Mfl0EzXtGo6YZ5DMRmpmj5rMDhxiYMeF14a9SO0ADKeJjVL0s5Ygr5xravhXnPixt
Tf66NipXWPup9fxFv/MDelbXv2Crd8sy++Cwz418uqP6QDy3UhcvqKpGVF9Ca0dtecL/znaIY4dW
fwFFjMmRCFEzePWbOscOO3RG+6rI4bqRzorQhCREYlhW34l1Z63nS8eM4GuHnExRcl8/ceCxdbvJ
vWZghwaePBLMS0b0T+F5sg4QdIZ0qp+yxOZao2+QS2GESbMScMwI/McXCEBA6WT4oQS4LDkcfMbI
epN7YOTbw2PbeaZNrAwSo5kYqht8hFtJ/N79y+gtel94wza6uCJtdZBaP08nDJE9JiwjfkRrW/gQ
wZ1EKMKefoP4SknLOP17jroT9G6/BKD0BNZXiYTraR4SAcR+hLQK/63kCtr2PTVvUYoTDquYBORG
EAO5+8GjOUEEDYeEQH7XP3jpK7WibKMmOY71TCsTN7GMFDmYHABV17B2c03A26NiMGu6OfnminEm
UqqpQalzP4B2eybMZkrTirDBVWiaLzPQVQMWsQhbBg4+dqGyMTDQQLCrMj7/Ykos/66VuNuPgdeg
ghOlkGeetZNBDXwblwpuP+lIvUbghmgFGKJ1hzMc56pqAtp6IMDo41e7kgwTyEb9rYu/r8UlHsG3
j+lvDWtxhYApw3H/yBvtFUf/U0aKUN+NZUVaur9ebx0obd48P3j2rSwnFjb4gkKJ6o1Swx3CReKk
u/0+gE4izX6Mn2bSJkqHvuDXDjKKAN8qvK+rdgoA3m6xiW71lBqAaL9AyC7l/f8JL8ckvFOQQ2dI
QCv5AL21gux9GONzP5+RK6wCjzYV9mHlnfVkZDm+lpl2PsautrexrRwgco0Y/S1foGdmka7i42d6
kEk+oxvcEHCPY8DaPu2Q0/UT7yWjCbP6r/GS64/z2YPZST5uttCScDLzJFDlcI/KUoQqfZxsmqLV
KOCY0vW1ImaNmpa56TnToJfrxs/ONJh3nu0/gbqhmN9h0QJ2PH0HKyRXlLIZb0M40cUa39ICMBDl
LkCVdtCNIg2pszw5xpS9hpR0ctyON8TDFJnvwtHHha3+aIXZgjXGNTAKFl4RveJsGNVfh4QIaC7J
PZqX84/Kg7c/gNZUR38/pFgWQ2nbNuRr1GL+xX47KiuV2ayy+5Kl4a3t/0QiziGZ1G+Q7xJbXEVQ
WQaKWtlBQ+dc1W/jZJYteOFnf0Agsj/ah2i+Y/BqS9dNqpMSsAG2QgKphPvcpZQeVWBPLMTcnOqC
G4nG3DP2YnFOYC+QrQmwGAfSOEZcdXGzvFaogFcs5kZfF61TGD0f8WtmbXp5gpOjrAVY473QgYGf
JlT/CURkPrSgtCDLi7//fVcKUwTC6OxGRUZ7FkTjSEYPhpJHu2+bu84iCh7DUsQohY8XB7gWCH8A
M/Z5u88TcJjZsN6EjSaDFmFDv1XvD1q5sNqAPfM+UVwHpGut37ycVbwXO+MnOihPxJYLXXNA3dyy
5UDcI2CS+CdB0PcXyQRF8Bdo/oxm7yb9618Q5xxMqnSaPL/93FRPQnqOX5hqsAMu5ilsQ6r1qmfe
q78fqjnxgLAPD74woal9N6WDrKTA6Iw5rhXvowCm32bqQEJXx13y5G6dMY3Iw8XNOCQBt+peJ3zQ
idkM1jfrNlvDKkUB4ERjdI2cjlz72DJyKMQBjX6quI2CjT2kuFLRBewmqntyNcAgCSfd4PFRLrE/
HXqwbhenvnf5hQ/SAxAhlQHbeleiocNutdDRdtPobmfJp+z5iEXNO9Y6eI/sTCpZ3u49mWFRRy1Z
Vg71SEZURIOhq9GNfYPGr8ixgDNy/YF7kRY4kf/1ZmyORbPjW2EATCeTR/glAvzReM+CnQQ2waRr
DF3HN78R+fWZO2pDeaZv6geZi6JXThVPlbWcD/lokqD7MZHDYDMpFHaDwA39cniAmVPcUu/rv9mK
ixLlUhwRCoG8rgSnqW6jUuu45W0W+MyOO8U6UJc3pMFKlXJ3kb0YrZ74h2J8rMOl3jFcnYKdC2AI
UUMQqGUm9y5F1vO/a2pK88GCoruskrLy+DN0pbQkKSoCQOSoaZ0zMOgJFekxcxJFA3weC7BtsF1v
58xWIPLO/UHIa64/D437fZd/YhhZt8G/HTZ2X8DtnTPT4x+LpeAF0jWBSecul6A/134IVng97GSv
pUqyQdBRF4jYP8SbvnZWmM8kB3XKJBnDwRA8cIMOiEy47mAaNkxY8AEFvqGtXLFtKq/rd/WPE4nX
8wFj5JqdBfu8bhypbjYPbZF8wipakWECbu8bkHQPHLYE+p+ggR8MOFcDJRpJhSXz3sp/Fs4p4s9c
L6F90ZNhzqAI8R2CkLIVOj3/TVyOC6eexpjG0PfJeDrmgdGJAuyxHSunfrl4sKc3odKbtrBb0J+7
NrfLn9XaMrGgHtIuWwCeDQdISQKlnBkW2uxfvrUFncd/ifWk7B/KNK96ivWbYvKmsou/+PDnwW6V
CjyblkOfJ4yHOVRThwy+U6ujCUejFh2a1JFluJ97qQ2xn8f3Yci3AVUt960pflVsvEGIO34CtQoh
3V/cJA7tHqt77EDql027twVp8ewh/yHDyeKH+tkYUXxN/13IbaOZtbagCuujV2PpndxSLJThL9rF
r/mfyDe9gs2aHtZCCwMAQJ/CWipZ9tXkDzk5eBlmEPyqYvBFZoVLpcG9EyLEOXoru81PD9a4GdEa
rFZYF2KzD+YbC5zZz0fgCmk/w8jSwDyjY9gLzUvFj56kxwlt7Vy7SN7FP3IxhmjGvWRAN5art5F5
W9jdL1uLHlgqnix854JPINQLu5T8C20mf20VbwCUi6A2Bj9w7pC87AgQToYlJiXgZWMDWhbMx3H9
7ugRQf66zUjd4a+03hT+qyayBSGdw7j6Px1X4v/ZPGaPg1eK0PlJEOCGPdeK9tgPDCnV05yawSLC
YLHTv96AUe3wa5KurKPNH1zoEOFjWo3MGlKvQ/kWJ90CPtY7gJOUlEWVKEGzDVO0CpHjs2DnQS7w
o/k2woXa0aM4mdfPzEZqEUSnCF45UYeSxBWPNi0QQLNA2ZB1z1L+qYos/5BXuakAJYs1jNY9zOzV
PE/r0tD9YCI1FkoT3b8C7foYM8ddmEf+39erplV02kZz33+zttOTJLGZsckedsVzMNqpDOdE2/KQ
LA64zms753VTIJefKulW59IyiZGV3WkS9qJKgeANX8ncFB+NQIb11Nl1H5Eg9NBI8Alq6DPSubiB
eZ6jjkmySQXudSlXUhQFD9CsWF58iFE9mALDLZ0WWql+035BPdRrtHLH+K6qmQSV8Xxj2u2rxCOh
nEIfUyCr0DkpeA2vMzEkB76PdJCo7DzOvVuJveAN22365YB/6u38kp+kr/NJ3tpog2miBMB/gNZU
FS+me59xXT/BJ1mu+bf5iNQnq+/QBCffg2h/NgXhCdcvjKsdATVS7jp6D8YkkNlRQeWzTssbj70H
YCa7CUKZtox8PvoVZs54wF5LcvuMn1L2MOJ5TsX8o8nY7T6X/IbgF/DHn1SqFFNUWS8yzxJEiMmr
iX/NhexlkmctlQIIWpbpdw+kOnACayjGvaLqhvf0LgcRJIxv/wI8NOY5re0FF4NEV3wf5Vj9SsH3
vuGqa0DOKE9mvNZndKCQXCDLjwr9dT5mkTXtNTTtYT/xQ9vdyIoCDzlTHGaNwqlC6c1yt8iPhpL2
/g13q136Njoro0VUKH3QDT1cdRtdWMsQwNEiOEtHk0Th6dWVDm6hgoEOQdBxUT4IDrLZAY7AenaQ
DhpgBT/8tw6BepTBxZ02Jd6X3e+8XRzAjCSLhyW57J9ciWzmc1Cd4XKp7jLCifO4zMsRnbDGDG44
j5D3NksrAYHR6+OnIjUvAt676Z1iwbz5/3peeC4Qv9vcdbQ9kn8QUMNVCcztUmt3buZEXbwmVpQF
Xf1V3e+frACvFUAu9nqq6qchB9xy9e9cE4Cew5vXhonqLhfJGPWi7BJJLAwsmQrmG7lhNwVGxwc4
gsfziBucoVZRdd3ybBBTPLRk5pEHxgDmnepY4xBqvIBNwSEebGCr89rCXtT/+y3uNj8nGsGQnMe8
bhjAo4e76i6JG6VBdvt/oDJoNW5igr+HdnW0h6LwHv9aI2ambAlwkHATRmib1gxWrKqHX9xdVvLa
5rsDXFhzn+W5ijnVKqGPgC35hFH7znjXmn+EofMFtU95H+Ue/fho/D0z+xZCf/amn1LJ/uizcjit
w4CwgVTH1xc8uE9CVO/4S+IE11QGr6ILpgYo6ExWarbsOdUalUxIMFS/LL4SYdY5Kh9Q8DIMYXOD
gveuBw9ZEbOF1V72l/li6jfu0GqiG8AptIIsfRtL9sVj3B9B1oAtAp4sX0lth++ihXH2g5F/PjD7
n0zChXpUhs8Qc3ucQGYDKGfRnzwpdrG0UxB3VTLHukThgdldUrn3Oy7mdwV6O9mqN7men/f4va72
yU8iE/XqOlZefc1X6hxjodWtkUTBFFhOUBHLNWMCgQtO2h/gWlt07U9m0OJy0lsceFOhxghEZmh/
XCi8ZhZl5S3jNVPo4EGzHbFNGi2seP0bkv+rUfQDevVj3uSSI4u4OyW0KVoMydFxQrIq0cSBn4si
I/7EsL4Na3eLreq59mRVT/6dAtFpMq3ry0QnXcKNFBrF4RNGCpSK9waizgEIoyfhlzbJXAKi6/Ow
Yuk3kvpKLe7NVHbcwhtLK7lIz+0zQo4/9nqhLwAiV0StbkOJ38rIUGcWYOHWFPGswrJFbvphb9ED
aqFColWVqZBe0JPvXkSKpnIzOoKSlmScXu3At/2hXHDloQV8n/9GWSY5V7+AzUIwZ2vMNkw2KB/Y
wqI3egnzh5xLJqrlVTXPEX9y+hZ8KkxygIyOwDZirDWPmusFczch23cIqgS3wabl7U3RFeq5anAZ
ZC6KtsFIvO7QYGnnM4gnpD2a4lafb59SKTMCBwns+MZoTR4U5wR8ALdsGhO7xiY8H9WgZLXGlKJ5
P3sBqBSko53UOFK9t61q6WEN2Mk07ttREwNNM27dIeKdpTjyPAqIi2lheTLaGFnGCVCNI9AK+jeu
lPuSjJipn9v3t/KTwvPpTveYBfRM79+ulyo9CltCMY6I7b0Ek8MOBDhsprhsFFjLPBSg0cY6aHa1
v3JbNBVuxTEw/nmrx9rRNgAFM2rlsxX2TvbljP4Oz9i28Z/L4V1oUm4ER85g81jDplbdhdfyYs+7
A4wAmunEvf+/S2Dn1I3RGj50c/w7T2i5hm/YtzaJuwJ5/i3sgobvR9DV2lfUKghM1bstp3aXkCO6
MXxKz3bCoAyiqTVuZrLhZwYXS8F4OMrh7iO9lUXb3Cf4TT52h10fwXPLHfp5fadz7eDbwWMjJu+C
lUHjVofgHncPr1s8YS2txdNVqJTOCLrPpyRXs0amjBNkWC26XW1+/RpORYHe1DVcP3jTVSF82DmJ
M+K93ERnLw5vS0m9CL6d2PMcTCGarNMJctt3pdjJrGjnxFYzIS5uZniV13VrzRwOUzcEMWVKIiKk
hIcUKXeqE4yfOzwgCnj1LHj+pKpzFzm6WN5+D9EIe3reUOPQYWfiCe+oHWpqpfki+UfGbqWYMqZo
ELoVPA/7eiMHo/jp5ntLVbIuqV+WJwrlPfKgec2TbiSUOGglFTlRoWF0rT9vdEYQHDyX5PPQhni0
TraHzPf3UeWtWAJFUF6HWyCT/2yl7L+/666Ru+wE4DuM2RSLgFL6fmV/A1rbSsPGoT0I3AVn1rL2
Dwa6nJAVMmv+2fG+K02OzvxTu7UCErxCnZkC0dUqPf9HidmnfnJVetujt13hRhYcIzJXJtIVREMC
APXx6JK3Pqyj3wtumcG2ra3i7fAWRNwyZRJ6lxane+oaNYfK5qAaciaKvwvsLpzJuUEyLJwOgFOv
x5rWjxikrKb2KTG8yFyiwjTGMlbiTvkx3UYinyLb5znDvRUJjB73HmmNtLvip9JdjvBTNDgPsvOM
u1804UyjXYqOpLfS/JVmcU7LvJ8HeymNcdIC0bECpyCTkH4BxgU+jqYKbzo2Tufzi8uY2COkvzZ1
4nkXmKA3B8L1SMTZ2ufjAHOQXfWiWyaDkhCxsuZMNTFSRtGljLdCZE9hNFu5V0wp3di8Qw3DxGOp
WMNB3KUDGl+HeK/IxCya29HcD86Qb7c3WBYZPxr94+7KXucr54b3H/8WqzjCqTPa5WZGhGqGoPU/
tKTXgGgb+gWRAA6gm3C99sHZeeF+3SsOwMZPxYEF9pfOe9j7krXigMQAk7xelxiwrIlpiijBr5ic
Dve7g775NzZe6zzz1leqMiWyjYr9koUvGUebhTlXtHmQaIuzdQ32x6ie0t/cHbCmU9/jnqbG89uF
dE5AuX/Lnb9E80x8DZ2fIFBdA/a8E738strOrUSShSfT1C/+mAbBSgrZ3uiO22A5IUlyxXYRkuJl
UfjSH7F7hMVaEC97sK5mHD0eC+CVxNIrXeVPN7161IbhhJ/bVqco10k6m+IqBVndb1NQMTE788Jg
NtqWLnrtlpw6XYyF89SkHmwqLm7pAy+gwb3hrHYZ0Wj1b4kZ5ccOe46nDjl23d2yUM4rYA5f/+Jn
fE1nEt+CHliLHFgYIPhS1qD1NqCjQ9fRLMLpAlbpx25rpeSeKKr54oD3+QfQTxbM/OX73pZBvdQX
yaQKW1NFDCgbk6MQA5Yep2LyClGfjhySpuqSMbV1If85SOafoIQLFhkv8Ixvnet0kknMZgnaINSl
yoAQ4GnKNRHoEOny+aYxCZCesQMaC/i+H5xn7arVP/jJOco+oQiwkZTWOIoBRMigjI90HMf4F2Ld
qyoWoseesyzDd/S/7S9aeG2Cc66zn/fbgm3LbHFfDzwSwyR59Fx61AYeHDyRQbyC5lpAjAA7z2ve
9OiQ8UjEesFCHzTIAen92w/ViQfCXVFli9cRHyBQT06EUQWedERckAtpGLYNH+mf3W7HGrz85y/3
biK39CrE2aSdJRB/210wdZCHBYFmPCFNpPCJcLDeugcedtOd31/V1RKT/7uR7Jdu0X2hmeJo3noO
kQ+7Ck8JyhGpO87gwQCTgnLtna+OdNSrfxUWGQMdCyGrhri85iQGpz603qTAdChjWdvu03tVeJF4
iKsGbcU81Ix+KbIW7zflRwcKO5975T3dqYYSDkPx3poN/CS1hmh4HHD6rvDwAIIEVNLMPWNCqDAx
FzgKR2obp5EgHNw/pBZ12zi31xcwVXl5MZ3Dn5kaoRMzwLdWxH+9E3F4Cdfc27p3ICGxl/y7v4p8
VvVzltezCIUeld6VQ7q8V55wR0Jg4vWHic7x4Fb+/EsEyVL3FlCcaocNgR7YJ3IM1LTm0rU32BFg
dnoY9WIlIkAyhy8UDCPGOLaC3xy7M37OWQMUbf/O9t59KGvCC99/RRc1ezJf8scPzqPm+Y5f68S/
Ha5xcSQgE+IeX6kuQ3Ir8MWT4O+3SiD+T5IIhBh4ievG8DwJcRpOJVx2OvU7kfaRXBgAs7N/iKYp
Kx1rhB/Hfi6otkb2jhi3IU/d4DyOxpsIkSThNMD2BnvMLraTu2Yx/BcDumZ11IbQk2gdhhAnRWEE
5RqzCl7u60Qa6ihY9Bu9JL6hLc0kCMKcpSMkI+TJj2wXkJxBvPmLUdcCjDxaa2nW1pzXD0lbVKSa
ub+4sE1qyWycEPboI6A25VId3KPuP/ye9b64JjWjfB2J6us3RvcBdzJByXKU4x93/XljwiUaWNJE
LHXAMBPRKrACRdsRz9BVGKFDttumdqPUELopUbWEBE1vvWzpk6ynO7HTigIUZCZ/6HLg4SH59wDY
CBuY7Df2SDvZSK6CvjEdpd+2FQ2AkQWRBt41UwcgkiTCQT/k7nIEkGeflEvjn52A1ZE6mZZZCef9
+f+R20yU1mrRklT70PT9Aq5KcZPuxYt3qr1JhT0EyKscjtmdF00xEsHogNgEB1ncclWD3t+xWkim
X/Ky54nePDGw8b4CGOvB/Kz6lDgA06vv1zEd3F2X0E9Y7G9bgrg+wnW4xMV1Ffz4pDZGhkIVnpIW
iEbfkjAyWSJDLjzvJ6WDhAV30xwUdYXl3OUNTm+0I0TFCTfldkGxSS6CF8BdqzINJQr1UmG3bKzp
McMIcWOXxSvELkY5fbAIMxeBHvKO71H1fy5Fqhica5qqe1ZLWeuHa2uJ8Oj2P00z1aiFcIWkZgk/
/WYZEcz3J2Dn34lAzGrq0BJhuWVF2dz3xIZ+Ezpa9ncTRZhLIS33HUq7BgkFXDKPK/rlc0URQONb
Ut6KJiYuJ1/7ZZ21f6wt3F4+XVofC8cz5u8lP3KHhU2PNlJzOiWbmDiOMxE4LEGFzJqx/ovAY3jy
Ey/M15W3lxsHOHJi61rmXoEtQvVig0YRcegkjbkNBW/961Dkak6zZJvDd89m+mEJfnUroPqKrMoP
56IEXe01V4+ItgGzxM04VVILvJjd7ajdva5FEjjImmxnbHvZqRHvUK4qmcfVwrEC0vaBmuRcQq6n
V/OopBGEAAiQgLVY/B+4iyhTyahSUNaUbKzaqUjvwIsmxnkVKe2TEG2XE1V34tVrLAPj9y6uYVSp
0TpcHzvMk5Us16ErT/c/TXigWedMpp/77lEYKeZPieCpQGQpRi4xLWrId8Ty2fyXhVN9lV5J4NTY
fam/Zp5N6Mgsf6jBpWr6XURm2GbE75T1ag+ZOZu/v3F4zQ0TRWqLd2VGyEqJ+mdgNzU0XG2IxTaT
DUBSH37Q90JebKVKOuPX8otaykzar1/e/0iBO5BWbUW/0IHA51BODo45Y+p/3KeWrWDTc9UvZUQD
J08ZQNcO78OcFQQWCcJldBT5NMenk4wfoQVsRM+ox+htQ05l0IhNGSjTWAXq+oTj0ByAy2Zka8Wm
x8RusEdshYjEmruZGIrrlwjqUHF8Cfp3pnL0BgwbXpGpGjx4K8q6EpRYQRxso8OAqzsQXhUz1AXL
OTHeBEVDd8WLLuW69PMcNG+Xd4VCSCFBcEkubaDeG5fh3hFuxsIPTTRyiHamiCry2fqoO81rrfcl
3GNmHlqgsgL5D60I0dwo4jDzc19MYr5w8ftdVzLWdLmdBTreVXstZEPH1ETss+NP1vCNzSiwELD1
r0e/ENgKP2DwCfqgmoDD7IpXwYteWmtJS8mSsWKSCELobKW9/f/5UeH8yZGvXbVrH9e41hp8rf6G
OXIGvldJVyq1PODDeSzgsb+uAUVmjX37AcMPU5L1/Kil6R/C8TpvN25KugOZbwpgGophtHB1Quzq
ayRKUUI1MZt4n/re8WSAc/JNN02Mupkusi11lTrV7tgXO8qNcTTKA1OCz7i9LxVoL5bgQlhamdEN
PhRarvKiZatQesadj3AaRezzqK8lAgGGuM5hp3nfcgrT0LAr8/ASWwlOZI//F44rCELl7W+gsyul
aYnvdqAxLH6CrJGqx6FfkIOnAucOpMWuXONu5gNyKkuX5bwH4AL8zGMPMY64P/TIy8Akusu5Wmbz
ZA9VDb5vC1SuoBrv8+mE64puLB00pJODRlpIeqAguMxbb70LRfFjP6QNUg4A4FORJ8TboBJrS8x5
QxvCdquQ4c3P4Xvgr35bGQ8nWcGwhbmt9sQRBx/E/XzKzlJ2xkquedcMo1Acpqh3btdsddLJgGvr
ex7imdALY5hlnGT+Ho/pHpUpcKiJPanBXR96gNjEZiaktEg0ada2CHpJ1dL53+bbbndwFDlyNQ9o
tNufSWEuluVsHdcRI2JiCsfLrZLQrCi2lH6P4WIq62t0K/qfFxMXn/mFnfeaOjjv6NGhwx3cxS3d
/mqSlxGIkAIL7WI6X+CK2mcPIHNmFM9V6e5FsXCNina+y3dwGfKCQ0FRJ293RYIC1qQ9RpogE5WO
CupafLwPHjUtmglB7gjGjlmaGudwTGm5kzflqQ3iXo7PgdvK4IuHG8gqoMXEqIUrdGyit2OYAuKD
lHBzP3MRNrx5+hE6GKbPFcf23Zedkhi03qr1WIwxc39YPd2gm/rtIslx+BkchsFkHUGDOC2iZuEn
cLhYFE+/TQE+2nCPGUD9VSHmoyljrB3+hRKg1nbYj4fF3Q0EqrvKITgoo24XhtyWrzmxCd4bfKvp
jhkg5b3Ww3VM2vrhCC/cXURUAPHtHE/VCz8dzYnx04YALwlHH77mAqdN2uLXGPKCkHUiPatMfuLl
2nwijJ/Pop1gtPe/gwpApK2PxrnluTnsSh7brm0zngXSginvE/VRwVtvjOAjShu7apfhGAb1TMsY
ZCx9oU8NGZQh6ih7uGTyONtgiU2AX0RJRbRzfNZ3/tA/eaf17FcCAqYAnznt5NQIeKVNMTykjG5U
wjnH5HLm86WQcmglyYCJao2dG3m2XZyAm3SuEVltePOqDAsSVc91a4Ij5A13syEbaLMBHzoeiupe
+X+YAqTN1EQ7I74fBGMQ3CeH0zDsTrhW8LqjUOOhfL2p+etu1RZu/5EZjgzIEIowKUOCR7wZq+28
lbJ99wkKI+jqzhAGXFO9h/RX8pparUfW96qPVj0RnqmxXIDZEsjjnw3IezDDTsYCcHQCNLf7P8qL
r4XBidRUa2OW4pWnyRvNRm1CnGDU735li+98vFXo4drY1gSFRnopPGFEVXuBXd7Lx8+tppD2+HNP
2M2mzxfqULwHmuX1UMqngMid74jY/y/tIqhfW3HjK1XYtAUVUev96dR0n5JCGtPmCltsbQzlAJpu
6NThmYSiovKjRXO6Tftf/BfTb8P8RPyZN8uxdM+GLeJoIkjZqlpLx45W/u884UtLVbzdt6V/02IF
FfIkyv2bebDJSoHEFauvJKaLXTvtAm682vy0KXlte7zSGkS1onDxKA3ufyaEPOqAisQanmx+lfbd
8as/7hxwtmb+vDgVH8ASnSaYkuu8NcaCLrXItPNIKTwyi4uleWu0qe3xpHElOLYkqE2+6BRxjapH
glMs2nKo7Z7xMfZiIJdEPplNdaCbngfdZESaKDsNhbtKo/C1whaSG94cz3FjjPexLYZJlMzQa2Oq
SKB9b1+MvH5hLpTWUgEX4q0Sk3qib8m/NxoqfM1ovrjClHJx9m02ziRj+Mg0deUYnG3TTVReOo8w
UStMqmQTKYyHnR1Uf6DT8udwfy18JfQzfy7kqhRCJDrbmNAvCD09OZbCF2sKhYeiyvsBhcqm5hxG
NCWi6txu0RCO5llF51ZWroesyuDZnXv521HF/szkIr3k+zLgcGvRfd6Mhd39MXtGvTgPwKh5pgVH
jSUs+54OZaCecZLE5KFh7+cNECRl7wgZMKAt5H2/oBiv5rO/62yGfzQxK2BFCsMlS/1hIA64xQMc
a1e3TuyKWFUuSbhHDYvygTUzl5qiSKsMbAM29xwY/mLwbnPbgj1jLXZRe732L0Uv1aEOM0UAMZKk
5O9gwxqENtx95lIK6VPeYmHuEmZhLRE+lhqPxTxVF4PMU5z6vqESXw2GuPtrK1W5dpDxIEug6IaW
N+JMXTJvlYVUTUQ+97ORe0js+9oe7ZnLXuJYgeBACzxlYxaZ/5dlqFe6/WCW0nFtE7+4coL13mPF
C9vvwQaeUgzQ3pgkKlB+jgf2D+mOZsZ0fvttvajmiYJMnjEqOtw7TGIRBp2blYh8tha4Llj90eDC
uSJHP0FpBftnSZItDyIAdrN7x9O+t5OenXDKC0FHuryBQo9c5xLJ3Gr5kp7IyLtmrHdN77yUmOLa
hEfCDGHFUnD1BFwj49fEkaolnQK8xTm7jGogWreAzQmj6F3mRcnSn009PMiu+RqztYBqiyPLqijl
jkurZ0OA3rcYbguM2H1qSzLrkN5r4gJkYYHlYTCheB+TWpiQM8ZoJ4w6vlclcBGH1cru1lRJerOH
5pF89t5fbkKWGqHja4KFD86X1FB1UB+I+jTmFx5aR2BPA4ps91kN5xFubajoX3QTYo7/7AFithNo
+ieSHsfB3RynuTV7BcS1WhfUQCzTLKIFRpI4f01M59dPPm+ye68CjFbVtJ7JqTPzOuV6PPryTOTB
qOxfAg0fAIvzC3P16Xwsm55x+Tx7Ggc+illjwDwl0TNA1Veo+np6A/WOFe5RYZWKz/prJfGyThpP
F+o8Lpa3PyR6g0b9icL7Abqn10knh2GvTmttkEOg736OxnrJ/pahU6ejb2hGYX7nsO7oqF7NqT6K
j2iPyqr6slCI0VpMtiZ6fIkD0raeM2eK2fCod9w+kr6fh1EXMrL52fktInR9G+U8LDvGec8qM3Ym
eSTvhwyHJ036KDFc8fdw0rrCiQVaVTM2/YqfJCkoefivQ/QY0T851Zt9IeAPt1MVNpEaN2DquIgo
VjfJC3SMoXFiEy3Xv49B5zHLtl4c6c2oF2ib48J27V5kloZaeRB0dvPk+KhE06vtEyi2uhP2DW4n
1t4lDaTVpRIkY3/qi2xmWRIOvczPa9JRL7o+UEkw1foTUsuuDFLP1kOqB9hR5P4wWzk/2VOqAAen
vVeDnxac0ANq2CcxXk5UFr8AFFfhRaCu8EQ1epMHbMhFxhkIX/sN9SJdc/ln5A0HzwGo3aUpC7Pu
3PViwrdxxxjY6bXAiM2iwGrC+H7uTiIyUuhqdZ/Kx2Y1E3DlkTWZUokRgPMRb5qCbPvll4cp6yuz
XBUKrU1A5h66pyJRWrFUazUetAkPDr8layPgqt5TUSPASDOxFvQb/pI7thahncZdZmMwme9zaE3s
w8p9J6/+o+mVFxqngpIHwnSmRb/zJSbvUBbUA5/s30yKUiN7c0eX/hy/87OCiMfTwSxe1l0NgdU5
GjmhHN80NpDDDR/E/irRqxh30kgRzdsxVmcL3LIiN/YjEkC0rD2xTNaqMzc4XFQi8ehpzu8/N0CZ
8Uylqzt/67k8Jn5q/qXRO2vsJf8PMWFsnKnQZp00RMgvNA+Q8DInr3wHv4GYqfelA96YO8YOl2PN
jjvfXbsvE0q1rVahI1ZO2S7Fmb8lubN/E7sop/LGZKIm2F5arNKdXJrPyfxtw0AZ/ab3sOJfXF8x
VV7LQye9NRgFrXmBNQaWCkhxFyN64SHFb6Dy3pv3qxJpGFgcgrrOeOIAC61dWiP9Y7VSM3yIiwl8
cUYXTs25rEGazMjRnR8eWvhpUZZO0Ow2e31cYtzwsS0chcHogaXPnk6ha5o+DJBr5HR+pW0APUu6
10BaH0Zh7UYYUYIRfCM1RUU7jMj5IvHoSkwH/7C4fahPB1z4qDk18dDMXmgK5N1O0j8QKW7BXn+s
mJ2EDkmliXlmWGmqNLjjYi6y6WktdgOPRhNY1+coG9U4+k+a5YMCDvNTHwYnnpF63+nb8r8jx99F
bFCka9aDrOrZyf2qE/skklbJeJCBqLd3JWKkZaVMZQxvab3wEJ6HY7UnpmfgG5yQMiyFOtrEnIQ8
9FCXyrl/JQH7/38QCSuOVgbm5MuHZAEX8rH7+hnL0z+JtR1cIrhXI7XFNTvTfZr2zhcdV19e5LMh
iu+/SZHXkXeONRfisxuBJ7GHealbXHwOp+EhLdUTbVIqYNRpzpWaYO27Dnk04oBRPumOfdGlKPJM
EaKje4eTRQ2qc+5i/V3SNTxQhNpAWjAh4+S4Lr/UjRhSq55d5XsP3hsRY/SDlg/lg6R50g8oDLnH
fB6GZ/BnhZtPtDjZIXpG0vmLRhvaopvrYRbIJ/Z4MUpXKRFR7DYlfH26qaOHJLVryIi8un90bS02
6+BXoxOKOvBDdCDv8R8qgOTcqAnR5VutD7uypbjQ7vZMPxLTlHARUx3pGaU531grSjHfGeviOI88
ndj9LDX8gZu14NoLKAIjjXO3sJ7Oyo5UQHHeXhzlRh4CJsZ/UCmnXOeY53qDg2831jvD1BZdJbRC
1aD7Fj+oGyTxgRxkCaxuEct77xDJ2Kd4+PfaM994+TnwiYfg69K2NpVsEVSwUMXByFeWRGNeSRYT
Xmy7c/uQLsKnNiTOexfrWWeXPD00u6cDbac3XGlkSDbQppvarVIuq8Bbk6FINeFMWmB7q6fcGwGO
73VLrWcEyWBlyPSApg0qxyr87dp14IgeOingxoX9ifFkgQfSVWuT3iRU/ZZIRg+kJcT5MR58ghdK
Wyr2VQPfFnTFhGcbp5CzfZ/L331R76gD6qOOio+Un8pjFYGYbDINWJvqxbIwjFb09DuIRPO1NOoF
bSEIeDJQgXjLht3MYaH71KJInsfi59X0Vw/bUJ5vASShzZ9KBKWJKl4cr0FvKsOKITPjZJIT9tHX
YG28hVJs/9xlczvqnFD9205n73yCeLuq/FjYgFkjGEQQVb5cvqDoEnmJvMdJcz6pfYzguU7pRDAb
INk2OX/75pjZ3ELKcBQZNHXZpese7U8N+lNtY9yF85Gf23RPN89qQFs+a9D8alwpI+dR+nTw2/5Z
CtUnCBgnJhpYjF9jsSNwnNW6F4YRd4QwDTtHDGzRq1z1MEEFYi5RTs9S3lPsJurnhU1Wfx6cloa+
bU9bVAu9I6OQMvQBd3c+wEkO9GgtBOf+xb0xFhKtdI0gFyMW5BMnI1Q3XdWaDjHRuxZVIt9UpZM+
K+MvEZJGkaXuY/Tr5WVu+OVZgJ8EwBR1Y/DZwS9nYdGOhE5mLOQ5ok/J33XeQ+l7ORTHbWb6NqNY
gqRKKJBN+lBm6zA/dsUz0NJ7J9IoK9kA6LIBop6rDhxAr3q5vf584V5qctm5/LB4fN6wlmNNgrML
ifFIcv8l+6JC33Qzb9Le2l4QxcCgx++48RYVUkbg79zt5vrLz4KTYc52Aei8sGRzq64iXkM3QYVe
KUNt4NKKGwQZXY/R2i0sWW2mIkGeIfZch8tZavobX331ucKVjM539hjBRCm6vXBJGwEx18zzfBD8
owoBhpuEEggRAHxyll5KbUZDYz/3kP5kaPR7WKfQ7VtXhdBuurkE03823zz0TQ1ZgUVWssTCnUDm
vUnGjYaTOtpjBzFEZ/gvCLZc0KWiRVcwZr9q44yWRQGP433LM/IyCvMO6XNhoY4tG0ZxD6YQFBGc
SO7JP71Hyy6PSl4hSmtYhZwy19vIi8//Gl9Cfx7qIKwC+rEPX/zfDBxTGo/yMv6JkcJLaw2e031w
Nuua/Tao5uJBpSD/NSRvf/SS/QQ9t3BkvhtPsVYWqPDsox6iHFBJGD9Z1b5jZwZFwFPDs+kYfdCk
BzCU4l7B78Lvaohij3WsAP+U+CsElIwRohqb4vsGU0M1CD9U0e4/PjQMOhquh/7gg1lOII3Z2kAZ
ocZHwtE9fPgasAdy+JT+xSdnPnpYGyK+nC83N138rJoqao/S0H1grlGyueGVBxIPlKGEnBOTV4oY
jRP25A8PamDoSqFXgckvvQN5wcxhfVWjA7QQa2dVMR0GXjBpNHS5zUVubwf09++TgaAzODlfuSML
jCLcwW9ZgR+sBPM87MJO1WEl3ErvaPlpE5CxQCm6EaLHWVcZ/Pc0Nb506uGpofphJPWa/CWHnvms
tL0uvoQxrrkquuuecZ8QBeNAtc/3PuyCFk9AQNguCd4+8tDcLE/GwTe6ewqsXMiHcoeQ9bf6Q1eU
Q9YT8blLaNl71nJUV1efw8cXfWVhFyxUcnGjU5SqhOhCm9H0Hxw+PSElGTM/QszyRJl89fzHacY7
hdalS9fzkeUT12nTuOPL6kCYB09ggUdEpcj7QDlZ/F5uQIJ+++RxgExJrCyl7Jxp2CMk3fMxizYs
QMYEUl21dY2DFTjrYNbxKtrKEaQHX1ZrMZkSHp+364H3WBpqsYtWHqUwEKTA10OuFlJqAkNyWwU0
58EJapZQlnoRRGUtS6MUHK+ztDDQmJpxu4qCLcyIfogBITtkDzzs88e86ELaOngdx9DoO/EirTW6
+Hll4UvrF5ZgmeRnDgm0m848ymbxnC+JADzffTfPwp9dpUsVcGiZFqL3wWqeQKArHXMEl84o1Ohg
rZ3ae+oxnLQuRZIw1K6wjQ0Y6WFJh0vCayg5xY2Pfs/r1w0KX6LcRtNsPQ5pWDcsta1lE3d8RVmW
mQpOED8EAzvAke9PyPzlSkR3ezG+xWAXBK0qO2pK1TbehOO2F/xi60BUV6nxNOoWmAiACtn5hlhV
i0L6xmaTm7mXNWjFZc1LlydFSBNNbIiX0+BZocgIuCwXydhlSXo9/T2K0l6ArJaqJ/FtpEBzjKK+
0RdbdsJNfO0VLxr3HMe3ktO9SbXfCybtY2ftTKkYRwYRASoeAVF+Q22Zj0RYV872rMVju3BLzlDz
ReLoX0LeN9PPMcHlTQX+qHvu6NYCL/f+o3J4BTX9pyfMl2kWqZ4TjMaA/8KS2+TRaQ40i1o70Rdw
2qx7BkrAydFRMiYlviNUatDsVF3kkunCToHoVD4jR/EVmqC1rbnK2n4X6XKTwmmTcu5tEkZb2eTq
yRbgjX2O+TnIn0rNaQNAoVfCk22LBhIsh5YZXzS6u6rEff5Wd6M/xQzYD1qnoBz522uLPA7NDtZX
MFnc7x3kvXN5IZ5n3qyhCL7vq1Ft+UCpz6/aFTwayuHPLb7LX5h5HRqRZZWfkdYP+wpmVq80XlCs
MQ8lNmcEwWHrmU32+jbTc5T72bY2n5/pQUqoqmEuh09GbiH26mTtorRgxUJ7WcNjUpC7MJthe/P1
dCDIsMfwSc7HivwNdczlvrjH+svdZfDrMRf0oH5yZ6sAmzoC+7b+mpPVGFJDmFQ0IJPk6eY7kBc2
eFo8QLE8VPre3YdO6AXoStWyEBRMVfEjdSsxqLfTL8jxgc+AwId45gqPfb49s4AD9IbNC0dOLsB0
k6bL+MpcdI53PWI85wVoR2G9QWJrYOzt7cz0GGi0YhamuanhvVYg5bRjX7R8NwHbqt4PqFkcnxbE
fU7Zhi6rZFrNgq7WInXaq9nCd/c5jKCtajmR/pOBgrdlTzF8zaj9oPV7cWR+oQpbzY+IEMWLq9YP
5uutoMlXCB9Sv4JyG1Kt2TPrHnLio4xwTIBqKTHWaSmn1cC2BXOlfujvDu2MO5B8uhfs3Vdf6WUT
JB2upxQqZLmtvBteTmkMz735WvGOZ6Q4f9i5WxzFNAAN9gPV2skjYoRsRgfn3aaoVkPxLqWUxvwC
yW7qYxe7VxU8S2NZKpzhZdOSPctM0MHvBVTq2wpYUeXdBd1Cxmf7JCYcNCbS4zokI7NhGN9vx0nQ
q6L2EllkIULa3hwOX9GA7jliJGPcdPoSirWgrjDpoq2oupTWqZDHchOnpM5j9+UbYXefk40V8c/K
Z5auBT4+PYHs4U2TIXrRUi+mwq/9YEoGKDu+6AgXZuB0vBrk8Hd4Hne8fNPkJM6PL4YxTf4oUWM1
SRIIXLE5wuzw9HOozTTFSZz35UgWQTS6mLHEy/g/t97ZmzXxg5YIBU9EwW93VGN571NZpyjho9xV
hThIdiXMiCftohKdrJfpTxQ6zmTpiz1WSAucdBupaNojfmkmCr5ZO2gACwZAh5b3s/1fmk2ByMA4
IXpg9khfGWRknBeBXAyqofexc/5ipDBXgW7W+bdUgoPqzLAd8i23W3kLnXGe1tUzSZSWg3k0wT5+
yGPt0AsitavdeOh4sx2spe/vILOQKbROqEsfnyAdOPaiuCRtkKUdc8Il+zsqICoDptDddq4qGmx2
JVdFf1ElIcAaULTUOmIg8gaX3GlqnQyTYtdE2LZHSD8LQZLWjYdRTyU6Bowsl9wI/xRIppE2DL+c
oQILu7PSnrCnkhztl1Ea5facbUijatOJ1Y1MsIeSvff3JfFgcwhKJuV4uMIaDE3Fh0wtzNxC3GBm
v8h3hRUuOv/wDx4MFC28DghzRGZ3/SHIowIgPxy2GH7CxB8ztpTPkaSaj+d23kc1a9HUesxvk2D/
Zr45Jy+QArzPAgEZEZVkZiXEr6/x1DWTAnHtsJqrHY8zCEWUjs3JvD1/nKytyZeldrs5gqMKU+xZ
X3n9Od3I6eVW9pMBII1fpLLN+QAeJiXTso0IMzXru/Oe3Xl/SvEp7oEeWiF1aZ3YEK9Csy6N4Er8
NZ/8v9CNZ1GY9tU+zFuMQGBZPYKeUG4DOrst9/RoS1+te0F36UC9icI3NOmp42bu4LPXO6uqWT1n
ydSJ11+r/PiKU5R0aABx6V05MoyKCri+eEx14Xp/RKbgpogg7UIFLl/NAkiZNXiQHHnEUVOLjB4H
fIJBv88tuqYRttEH01TdedbUIeZnliWUbwEfgK+xydJ1+FBgONeAT18hRiN6o4u++ovbPIom80DT
XxZzQ5gfeL8P9UYc3qyEANRRpo7slRCZR2yKwJ6o0AdHtXrr54BPt4UeGRFe5CovesBPvLwqU2jo
Wq19Ur3pgg29XUXTyTdC1k9kMI22jJuD0IW+uxFJNGbttT2jmi9LVfgU1Q5512J++xHnbuIW8WNC
mPNaYwlAVWQPWCM+tn3ZDNUqV0PvpRI3d7rQvGSsINo8tjsoXFc2dpG9fIaJfWJ+pHcrzJef4X6F
SQWmDJjbNqmsCsv/Wtybzg9V6Ha4Hd5IRv7K62/GN1u3yOuHBZ2dkUqD2nXwo4z/Vd5tD8mJRwIm
Hu+r9pp5pyCd+btGm2YVj7gmGRnGUeDCFgBPS81LUTeMOt6UbO1cMjcAsWgrJQziO8yGTAUMJ28e
Xx0RH2gbUF8/sfazBoR1Y+AHVxMdS1YaFOH3LBjyMU/iO6XO3nyS3cc+0QSet5T4XQCH/7hyL+LQ
PTcD3MS9ld7chESrZc6dYN+Pg31wPvR1yowTkpgCK0k0TR5ebD538xzKlnAE+P2GPESx+9LQttWu
3JyiodALwoaBDmFUdd8ujDMTQRLlmAnoOYTk0uELQlaCiTdJfr77x6ieI5CtSL/O4lRgS+bZn+JQ
YS7Sw968ePofuLE7FZzRCmxHRoqmNTE0v8khxAop+fCBgXhFfG9PiFEiM5KLCfzviMbc8gEnp+Rv
Wp06IfRRby1EtpOXAksqxWIvNYNihtuOs3MVFxLiEFsrxBbVHrl9VOaAZKQBW3cC+g9L3fdRXIQw
ml+Rz1tAPv02HsOF+RnvFtMms3Y+WhiZebTw29EfWHuoB5wl3jKU3OiYE8SQYC5ieOLY1cIAKXaL
kb8MYt5fR9UEhUh6gnnAEfdtRRsP6bmxyNgBB7oN07gcaG8BjvILMBVi7aAewCzlFmqDpdKM/9l/
eVjaTzI92b6J7lVnBeL3k+pjH2I/TIzndt43zZAX9rmN0vbuvGZbCK2Rv2kwsFOfUdL3c9d1xMUR
4DWQLwT5D4gW17ZfS/I7WZYnfRDdKDqf/afXf7Bv51VjhrXUEe3xOM96FNb708R6KYk6UBUjhrr9
IEFQLz9ZIOXd3QaLpKbjfx4V38yHuzhkSJGB1w9CqZCu0M1ExIelaeD5Nrbq4FLgpveXbP0warTM
hH2i+7n3BQS60UbTy21PblGCs9RK6e9E49qBcTdKXkdRUu4vx8EE+ckSygvNI321bhvDQrN50lIe
7VJzW7ILhPmRwQxrrGU0YBAJsAixwyfEwugMQAlaQVyO89X5iP1nPHX2/W84aE0upxmjbnV1UEyS
QosIKkuhvTitHCD8YT1xB5NGyjYLOqdape99KmBxQJZ10le7dGHsIi8ZnkGWEqAiXpWcVCNRIMef
3ikK2U+kI74wJ3cms10uEd/ONaZUlfiypNOa8BnO6PQd1ZnitdUMqlNnrcCv8GwUBgDvt885mFp8
dpOW0mJV+eRNEDqo34UOMprwo0cHx91qj+c0Hc8B9+KGiWcH+YrLHIG/GXq7Do7dUKkXMG12l2bP
b6yEEr1MZggq3HyT8h57uUf4ATjjrnpeCoBXBw6gm0gmHlqCe6nfDRj/owlOwfa+IfcZue0jyE1x
qmB998OU9mserHoTqQLFXBUJjSA7d4y/4wHoC9GTOjSkBT6cqcUfmRCks4niRXdavAn4ptBdT3w/
rD2Qv1zmqHr2ox4GpeZ1ChchniFn24uhqekBp6jGqRIVajdRPM0XdtSTt2+q0b29oNB9PlSNri0m
ZBO7/g0z28In3YnL7tdT2Xus0iENBPSTKQpl/LNRSUeSYrCBWqLm/B3ccf95Su9f1I8+YJ6pGlVC
QnRGGZ8bEujQSquz8/eb3f8/IAVKkLDgGUMHkl7MEN+zozTaQBYZbVIQktyX6T0KplAkco0ZEqFX
4FpG0hUOdfVK9ulWMeGvso2EbHlDwtwmH/83xPIe48lc6zMUfJo/3Z2qTGyGaPflzyWbWyfuHKNQ
8RmCHbXPQ1S2iEcAnBzIchRjpzRqkrO8ram8aV+SiAbLkG/RwqR97LDftXcTnqoMH+wH/+ViYvYL
UXGcTQGM1DpwoVzTED1OdeB7OQMGUZ7Vu8X+rjVBupywxJEkBeQuWea+rG/Yx2lRtWF9Jp573aeA
ei08GecoPULiRKg3lHnF2xn3aEjpOr1VoyIhRMO+U6+DGVywYFzh8Akc4J7nzK+AfYUr4nHIfHq5
h4R/cjix3XPQFBK8XSzP2bjLSHAjto3xtOZYKPmXhpwaMQQ+9t/fxkj6E/18G3nxsK3xFJsKWLwv
PDRNZE3n7grGvW1GOeEPIbkg8bfKgjlEaVNvNwZE8kfMnJAPWxMoEQDA8PWl+yOTuHSDmQAHKmd/
mDeAHKu5Gs8YoClHRyev4FJm1wivSC90kfJU8hhbkVh145c23FhNFV3Kte8/d1n5e8L42Iu4NsvU
QNp0FXndZPxQ7lu7E2oLqwhtcmSyKleDE5AIs/9kT/YmK6lCMAs7pa6Mx8J/ycYw5RnHXMsHvnkk
GlgETjh3Q1pwx9HKtYWnmZ2GfK9u23Fdh9spnz4F71UoH44XLHJUz9qIGBVDABsuPjGbu/cXFcmN
iZpfVjZzbKI4qx4+v86ZFsNxutKl9JC3raWPuBY3dMTitiYT/UP6brPRP34KUgitQ8KUYL39BT7a
QAzFNGo967TLkzRKPzkXdk7tSDoFFY+egK36cd3tTGg8u0exfkAh9jmBpXfulLtgJdVBylJW/S9O
4Mec5yNOjyWnvFSGKovTiZQtr4syzMeqDZb73azE8mnnTuVoUG0Dsn0iqAJmuliYmE/aSyW0TeHM
b2vg3JzwoVSQptmucI6JY0YLcfR73/PbtJ0yuaGbjnfLAY5wt3T7Ol7lK0MLXp0H3e0a3dDa3Z6N
YNrB356CYtkoI/Pf+URDy6OkI45AudanI7WRv/74pjjicITQVLwfL/2vNiv+8Xkzo7rx+GPUeeOv
7F91ZHROp2Sm8g7FI/pnXx4J9F+EMrARNWOGpjFTvJYVzeTVvtJSzH5KIsVAZ0u3hPPkzMqqavfQ
pNlXKmnIPDiliq4z4q89uAv1xW+/Zew5KqwcitkDzIy8/o1qkHhNXTHVIJ503TMc4pHEOsJJoVxd
cd8ditPFPvpnAX4nrhrsZGl97T+KxBvlwrJ9pc3J8ZlIeBIVSx5MEiy3DAN6NujSbZ7j2uPJglfz
JvFfzCFB8tfe+66DMLY4D6/OvIqFaZ9N0YpW7Opy8knZuCx7lJ3yZb4CWHI8F8gScb0uBz1eGds5
PVdWhoPxNhaG6Yxbe/iLdoDs3p8BYb5zpJmBBOLFvLM+EMljuIzTOGJbkBgmMhgb3M+Igjajkav2
DNMiv1M1nmRJtjOWWX3uI/NqjYkGJqqdd3wRBGacElu9/aRsUYS862bIHO+lMnxPF9xvvy5oPOT6
QyPq5zuOwgio/wmzCq72gdXeV6P/d0Mwce1hF7ceWPwGVX1kNCQxtumIMqaSl92t9XwyYeKE2EbA
UXCE6pqa/YqIMfmrLx2s+ZMPjaPiRidwe06wRTO+ptF8xxVQx1eugbAtcwiNQ9RooBwVwWHbRRTg
kpnUFnMk/kR8kX4Jg5TyuuOelU03JLtn0ZLhQsBibN/cwhtXtbvoMKq5CsNDNMA7GJShrySNnc67
AVU3B72oo+LMGsKkc4uqLN6NaUyb0QZQAKrYArjDptIgb1Qbesm6AEq2Q0lPIMF3SOzoI9E+rCcU
jpy4uxsA0+FAp665luIsecvJK0CA8eUyX5HAwAtp6MtKQG/F4GyxZWfHWZdf+EkgZaVPRv4kaNaF
wUohpD9iSeYvPLq0Pu1hTTPd7MFeB8LRVD0DN9sOvy8bPLSwVDB/kpDPsOfxfApy3QE23590pbkl
jIkzTeSwW8nWrOKs5y6/HgCdVzLztqd1XEunYx1UmxAqhVFj1oallJ2awzL3j+RZgJncy2STSO0C
SjsHURN7KTulJOLTUaZo4YVCiu0gCrpqzWAR2CBZDo1of8Z0NOHCsbwcnLV739uZrSd4tlFqhx42
K89HoKLbG0a+A/L6jGjkCXmx2zrd8CcvDmraCJWN7DTLICwe7XzY69nc6AjHfjuPitepW700Pd/m
vLQJLe6qTtpr0N16+NRVDIZ+iRguzNVQqjRfLWRzPWP3mc1IHiZugBKXvLKl5XBWlCK2jDZRKFaa
hV0uCn7RyZVKUx7q/pXfRH4Ugoq6sFFi6dZbDXgItRI/A9qW8YX8UOITJZHpe5gOrJVXW0JN/OBS
xjqN2iGDrXs2zykLc+Ec67PGPv1CM6Bz7G5aWcjQ2XK3NXFNxZU0moHDNglmUUlnwqI3qnitbV6A
lvZZwY5cAEDaJVIn+1BwdNThvZJa2DlhkYGLpa8okKkEng8G60iL9iph6mhr9kUXPdiOZ20cVG56
/6bpcd7oxVlioF+U+aCTc2Of/+ETMdFsggKz1wVaA3fcTCJANZnDL+qJU79Y1PHJMp0updxL94g0
bopVEvfF2yy9e3T4pBJHPnWoMWpi+1KVFgBkFhPnpi3EYBQylFhMqXfzIQ/WpHWwiHFUJPRjH4tU
0EuaLz7YPRztquapo6i4WTYPsAv4gL2MJatMm1Do7MPVCHQ65BMgYK0QmOx+RsZzxJoSeE45mCIy
ezed/dYbmkwQAi0aDkdee4kVAriqefPLGNoJBvc6v3vtq/15i38RctZRbROYUY70xhYnGgrfJm61
4nJerEfaQUttDEOIgpx9GjM/beisyd/FV2Xt68T+6y8pDXPLQv3uZky/Mjf66FYKgxWNcCVdi8b0
Va2/mY8y204ysl8FN9qetmh+wTsGhOJ8b8A6tcnSA7JcajUcOLiTe4wjuh95qMOEJNoiiVG8rYwT
pdRRFhJ26RXr/jYsX8//aeRznMhZGXGWRkcROfizRAjuO0+hKkAhGrK5mIxlcxuNBrbo9+htfLrv
+dfx3AAsWEyliqzjGncAhhwzZdFYvsMcDYrDOqbpvrDJfh/hwhLRSwOmFGvqazuWVPRqvyh9Hgjg
iAQf3XkC1q4Vg8J5AJBVidxeN3NeCwsU8xHDM8bpSht0JuIwVl39fuW9n+1e+s0GHL69jz+LPaiq
GrL+sPexBP6ZVDGGMN4lHMe5HLCDuaALQDwj8mFvZokM2ldMgK/oR6cR+lAVLpT8Kszk2pkUKq3S
qCgdr+GGAF0HZO3BzUiQDw6BZd9n5v2cZMZ89pirP7/XTtkfWu8mH3KFiyrEt2Ty0lAIPfGzk7OS
F6HuoGlHvduhEA7DtHrgnke9GFMq7DH60mCPwr5iZRDYOMZClKPzZm6VNBr4VMtBbSoOuqOWBqej
YhIOYYODxrOF1NIgULU5gK6/0BN7ppsWnR1Y6Jrr84Yw6bvbQ4MOxTa7wvwyZJB503kFMOzeXLOS
wov0xuMlby5dXYz5uhkW03ycTuPFY0uElFxtaJcxHpYOxKv8M1ZTdBdeyggdAIPrwhiAneWAXuJM
HejsvyhlYtacxIMIL8kLHefHlBydCvDgyB7YXo6YYALJA0duIfS0phblY1r5n38hr25uAVycvMrB
AGWmeVTVOwj4jnLIigI6ZZHHckDfZLtYXcBOCgTwXwgrv1i2qpReoQ3NQOT8BVGDX35216Aq7eu6
81ssyQ/0AA68+XiA+xCXgC/B44BH+3Bk+LjAHDh6I5xLyOtsKSIx27sH0BovkjODjR67FZ3pC1LZ
fjLzun1YZISnfiYkSk2K+srVcjbF7cmDsDSDOtOrOr0sJiHhqDggLQZI1aLHDXiYrIXg4fipHDZN
3P10NDKwYL9AfY+3IfQ896slP05h8aU8aCDLldu5aOnYHVWugdWqZbIWk3FAaZ4IeVIdFNa8xhfD
AlfjgoOu36YWR7CVr+lF1VFw4HEb4GemBS2E8XztKRh1FSWWyLq3FsyqS3JXVpzCeSj5NIclAwI9
ZArr4ER5j1JfjkIYdyPvn5nSypHSlqANc0UItAX4vI4e10KrseBJ3KYgdSArzR79JEyZmFhHW7Ss
HvH+PigZCnQ5IBjF/bGisGvSG+AmHOalGI98AXLoqm9HiyX1IN15HlGkTaqqoYJeWgj/X7UprmBF
T+A/20QfDxEK4Patvp8YkBpPDpV0cAjzD3gSjH30vTiPw+a0urHcuDJt2KgBjUzXfXKpfNiyUfvy
CXjPtAwcSMrJWRcQuI6s/OZPQulFkb0vYkqPHMyOS+g8nBog0kDuN4Wi7FWaXm54FGoV7Q0M0Qiz
8q0Q13TJKBjU2t4J0AniQmQ2nSgSbdzOUZ6vKzXhoKtB/NjUTgEaXSuyK2rqOuP2+dVL/yCZk0z0
BKTu4kUovN34vWCMFaWlK2X7wS7+Ze4BhSgp39edVCfc7K4hqIdAr9nKdXmmJc3dobyDbGnVBj1M
FHvfzwZnJ40y0Du+pcxSZvrSpTUhYOqdAt5QtJE9h+WUWXJNBZg6F7NNGBFKSz3X9YxpO5L2aSEo
0Z7Xgtr2Yw7RyKIsHWMvp698VVrd07UO9Lb1ZmFYYz3LIaPqP6WDZZzjVPHLFLwkPw7qGxWNQKtL
Kkr7r+Qgj9jPIeyJy+C9+JuZUXOz+Jw+TgsRiWq8ZvlWK0u7vAshBCqZXTc0AJeGfu+bmMOejEVT
jMl5BcVD6Yvv9esLTOJpns0zF9wXtCtTKjiVtdoNIxOEnSm8QdWtAqzd1OVfj7m8W+/4/C4ZuKEy
t/gO56sDhbNQXbhdwt+y+HXgyBWjtYGAuVIoESnD37zy/wTPj09bJC8Z3nJY0KUmkf/N/yMVhEr4
IX/9JL9LNStRDOdCC0u5c1IHYvU9DwONNF9XY98NuGgUBKG9Vv51CiUOFI4HSSg/Mp+z03iq6gsd
CidqX9GhF1rtp4wGgBn8v8PlTCl/x2iCRHOBEBl3PPRO1nztVohrrFwBPQKWo3eNarF6HnBOq/mW
UhaTDv8vGUYeoQXiW+v4FQ8yEvxrP7Lsnr2VBrBMYdb67+AKzQSq2kOfD8G1amZuRptuFV0dO5dd
qKqm0GhAjZZO1Ks8efC2RioUVsNxpWxU4p52Q2k8yz0UZ0YPphandGhAwo5K6dzc9I3kPcoUHw9S
98hKFTkNrUYjh8SOj4Sq20tHRDRURrd6l9SROgrvEcGSWSSWC2zG7rxMU/P15leGnD9C9qADQqpg
K9VN6rRcODhPYgRKb7cO6rdu3n5K9/s6uPiUAb850HWtFp32rUWO0gQwk7qDaDy1mVI+RvpSgnWc
1XKxlmsrWHFQRFGvx0A6Ld9sS+79gG1fcy66kaooR3J7ooTkXwflzY/Rn+Bi1TyRwwbDTgOwnhJW
SqFQDM24ywwI9CMyZWCtT3lbYeTMjxP85fLQDQLY3KPZFNs7G/KdvMENlxoAs8My50o968oRHPg+
Hpil8f8MVpAOme1ShGp5IR02EBYfdNMk982FmN30ayaO0x/9DZDIN0nLdsBDzkbBEmDkcOVRd0VX
otTSZVkad7nuO96jy1GRzsqpCFaiIJbAVlYqW0HBUTx07fkm20l94vpaEhoTq02BzbLpI1yd0zYf
N8qAsgcXN3wexIok0Lnd4NQ6FD8EVVqIcEOHwJyMeKTXoWMC54KUyfrPktHBqLPMH6Tcz3qPLvb1
5VQDy4VoRYdhByqPBEAZPKnxBFCZgKlziav8b5XzhmfJz1i8tM9rTClBg2Xb5ycCXp+j4Fb9Q9MP
HpVt0wWlmHEAKIZbROMCWsDnpsgjBMwnK1BoNekG4fYBdJQZMS4576d+qP6WQ+GRdjCof0E3CSWI
yPnkW2rTE0ERo7NS0Toblpeo0Ho88z5JnJRslVtxn7lHhQ48P1MZfob1MrYIX237PGSOCSu30q72
lHoi+cYVZzmUibeaaUnNe/NAuJGXhPSpIvuIc4Yr4/J7gftQx09WrsLSdzm/Rc3TEuWlZGGVdnOG
j34l0O+v0ovHTEP+uzM12ysxEl7Q2LdehtFf0QwZVSi6mWVpt3JMYlywOLE1xoA/IVAqxstj3rtk
Mk4ijheDXVn2JGvpCrp2KQV7r0sOUwLCKshWEk011zA5ojQ2K1+WzcTkKaWOLzntCqHaCOhbKkrR
LgZ7UqoP3WOsMGRk/HLV/FaQlMkwtYjV/zPCnhhRzQr7tYfDBYZttXaEIJt1Dxfet3FEnIH+9fqL
6vyagnK91ypED5pnG/TlmIwFG0AFH5cRdvAgkWhH7uuUFzcpmMxJPK7PjdayebyhvVsQ5Doi4GdL
rbWdIgTDZZhjglopFpviEl0TsTbvE57mhsdoovbSqc3nQn1BD54bheZFYbAumqPwcALiD826moHd
wZhdK4tkbG5GsQKW/DRHaQav9hxPcjaspJSEjJp2lJuKZuxC8i8bo0foxJX9JoUNuN+eficuNmte
TYdy2w/oz43UD34ukIMq2J+xDCDXFA2Km4uB4NU2zW8MKnxYCr7497aOZYKH1eMG17yIdExP/fWy
TTrkNkMVGvi/sjkN7ky4xj+nIEoHGqbVFP00yOL7SIZGwYBFv76gNG1onSQUFQR4eoagwewbmPNg
bPGHAeOnrU4uyZYqVjoa1UIG6MdcATXRrvcgl7VDZyd7FQ3OKrhCsSM06JDd9CgfIo5jn4FaZCGY
wkmFFlBPYCiPJR4T/BhcpB/wZBqeah9I8CyTG+S1UiJnNQVC/XqN3QYltMnwo8I131j+ZTuDZMWg
+GK8yv+7XD5hz00m4v1tUhZ6dlzdAozBGa2TObz1xNLZuRlxHIQzJQsla/tvENEBlPwZCQDJ5pkI
9XN/127Ug7/D8FCO9vZMXk/wkyjt44gwfjTqN9t2t8YeWkd51I6n1/LhU2Rf8NQqYSt+5k4g9ka2
Y3mobt0/aeP5pB8Vm6U150gz90EAdxzCvH25E4wqEAMRGdKbhsjybPfBXVIVumxo6m+c7dM2rocM
SVXhr3aV0FJM6A81398bqMxVmfyMAnT3VqIjyorW8GGMkuA/H1mw2fWqoasG/eUZ3DGpot0nCCz+
C8hvV6ftgqo21FOXmjYbG1JXMj/uhPiUNFy8n9ILrx5Z3nHbmPaI2AXFZr92dQwm/bgS92J0IPT5
RQMm2/S3rvrY3xB/SIujoZ8JOPAM8k35ymTRHgt7zkkKaJ/gU401V8RclgyL9nltQ/ceoDGZS7Gb
VwLcnapNJ8oN33EDz1W4ZcQdRM8IY5E/Eda/i/ljPXGtii9C7SyYk7CS2bYQmnWHFFWOxfVdMhIM
c7a81b6xfrgCCNRHiNkWw6bMEGhJMjr6MP83c29Pcihbo5VBg2OFlC0gF2Csj5X8BQgXC622fVe0
Iu4SViU3NPgJDpgGbDDyxWKe+8BmdfauVnvULYjvmPf5aDx8nG1QqRftMqZvN9MWs1N3LzUGLCy0
HstNcwudGlqcyxVltue/EkARslLXbcjmRBwmTyoaLsaa+PXqSfTNEMChl3xZ/uvRbDSkw0u9Igjr
1TQEnjac7fR3hO8TTmXGktwWWnMUPQK23Drgv1GGIVpsjDTf9dc5WaVEl9bssSSsToBwC+vFaly/
q+ExguOELwv/IaJuRwdCPmiLrjtG+2McvNoPb+0BxglbtamM/qIrflRTeqGozJSPO7KD9NYFCIXy
RIYEOKa5pLDS3QhpWGM4L6V+FXo9ejGgI9UqYNX8lbHGbsQvOwr6XgTsQf53iIg+u7oTu66qjez/
Cy3j+gt96rykOPK6THLYi3ZIdxhtwhZgBB2NuuqAZwzwtmWRedAAr2IntCt4NncBxBLy1xXHmeZh
cUTPAMy8mNsAghiLiztP9rsZ28pzLWC+Q0xC3Zif79DHzzdlAJamaC3krU0ylTlQPKjJjwjtE+M6
8barYJOmV+NPnhCsc3Q+IjnXqTCj1DNXFCiC/quK7glSXyFCP6SyCTDVaTeI5oJh7pom9yg9p896
yjx7gDFaO/VakLesxD9Rw/iHbwAtFKiJNfx6afvswgPCOvzuFi0y5Wqjd7lgGmuyD8Wv1CV3/dr6
p1/Wdkxv78f9AYyMm/iC7Lgfp6sHvcn6THiq4uPVGqzr2bOWRjD7OTzQAF7AlVpdJqiU4QjlfOIS
kmhMbYwhrQNV4bVLUPOEycARU2GH+N9WCcejzaVJoXXTIEsJY+JkMfKPygjRD0HJPSiB+Ux4It+M
3upcUBFn6lL7RLeRRIOGwFPOE0NKNTVl8wrg1A6ilRD7dVVUT2uYIX1qF+U1z4QiLAmEDTHtfNSR
2YTdGY90ignEMYs/Pap1G/tA1DJP9yJhFmKRPm5v6SDSsC8dU/edU4+MEl6HlSatBxqbbCCGErmU
5OrwzSWAJh3yHBv46s5JdXAo0mIARK0SGQlqWMlOlVmoVTXXLVdU3QW5YDHlII54aH3DUy5j+c6V
5jxmpksSEb1ZVMT2QBCSlEXnVpWMLYTgqlr34EM9aPMC2gEj+ttGrf3s7frsx1CGJboXR0qED/Bd
KHNs7w2RmHhpy57CeMskwxV0fXXkmiuV1R3Lnpc68K0+zhQT3Js0qDhIezN7zL4uMbSBbVvWTe/T
0ItXV8xOGfQrHcXKrIzfMyWz2A7VgJ4bAWMDuRpmds1Z42ePh3epaWFtFF0aFqgpEc0zuhBVxlyl
mXBA+i9jB6kC4vGhMtlhGeFKpTx8gIk5NRSSn8/j6WDED8f1pD/Jj6MYcUf3AQ5akANwhgR73Ubj
iNxTkQ21tMIK1aciWo24OkRWBslkKqdbqMoKj7w0UIchkGzDuxURiuslXa505UJX+0ssQrmuxb7W
Ac2Lo1zbOvco2OV048hVLZKVZLUKSTtbGyYEJpasgrt9wbK70SkTyzdFOPMCKvgkUIL33K8ptAo6
I4ywEcTKBI1ysF1nILXTetp9eUEOe3YN+5HUVITQqmu9geWDPjMtCgTn2a0YpvOy7EC4Jol9SOQ6
TFN1fk+EJflRliUpMmF39j+OnubbpfJfb5rzfheHjUiMxkrf9WsXbArC/yiJCHT0otLyAygSHQY6
Wy8LZlWLhhlYCgKeLC9MOgitgw4XUWxX4l8oloXoq+xzE3vvSdrwYQSMTDfpXb5n/zRhIOB4HJYl
qno87T3SnliWA+WrW1TJrQVPBZzHhYnTkvb577eG0JC/Cxts7XlB6h5jP7HhKHKcyFUL+xz9iTm6
rFIB///EbQN0NkbJIqZZCG+wnxbaUy5Vh8ibsNiOmyfnjUyRUYfW6G1xR6ddElPyL6/+frwoV5lC
DOqTKPxtECPXeUJbuPYNGWNBaEOFOu2fpukmE4aLoYHts6YmKkNHMA7rMdzYwkjFGOYBiGx8KBkV
CvTDciMqVhmd244ifgqiJ/o+Qem1F6kScQJvpQzGbDKya6wq94QnYPh7Gf3KBfcseGKEmRQdcAdT
biGWPilqy7R0l6jWO7ESijmoopLJHNk0xYWDrOfdBZbW732WMuGtjA14W8gDB1MmX8th5Gt3NcZV
aIogO0TLaYIKLPRl3V1njX8izf1sv/MxxvahJT+MEYSTBTXlJ/jVwKx3zLmO3+4i1A52VOQy/URc
uaPp83tqZrEdluwXhCVjIDJgeMtTcOLn+BUYrY41fms5Y6eMJrMsvj8M9rihYwNInZctxNbfkAB2
12YEo/XwGWqa4oM54O5oG+4cAXDo8Fvjm/tz1tmN0hF7wnAAeYB1wIEuJ2tVz0doNu9bH80IXhOH
115L4fFW0PYZFjP/+z9XUY5J0bZcA89nDuNb663GvgDHyyGtiaK8B+p+jLP5RWBJ/kq9sRlpnENx
oa1i7YjdzMvrh4o694rHZlsp2HPWeEozMhVpSrFtTusZzw/lIC7aiVay0beqfWDEmwXjboAgM6WP
2dSIL/af0X6k5miX9dSg+Ep9HzU3HBmPmQ1Ox8xUyVnbDg1p68libCbFtPyflix5K3hsytsxV2Kj
8D7M8U6gIGaMoMFZzFQp6YUgHBP2OOcz91fKqGNWUZA10UY3z0/4B5+kb2WMhVJn0ueTazV8aqAD
3YYjPiRyO2kb51RMHiRXyP5PQYDZAH4x9ecfq8SJOfj0iL9BsMFw4qGdeMJ6Fdw55P9/qN+rbWTl
7akMnQjN2bF7iltrmIdtV5IIcQ0F67Kokn/aJlzTOrZmfm44lHcLarlJnN9GM+vYmrVQ8/QY9bVi
MPwyMq/5OFKlTtSyOqXKn7cpeQoRRmdGxjkIo37WTde6hD8z6k+P5DnRnjRwC4HDXEcdzWV6o4vF
OaJ3AuuueCOWeSRYfah/W/M16rWQCofUDXG/IOHSD/cyT23o6D549SrLxe6FAmGggqnJa8N8TaGB
GI+7R3IH0L4Q2zOUbXdTTX+D/nT57ENQ2Yc6A/IIQg9Ud872zKPgg5u0uopSGMdT7VRx8aoFpqYo
1x9mbhCN4jPjjJ6DEHU8dBxcP68PbhNMU2/+4ISnD81tb+8AEPa1os2iZNKCvzcKz2Zt9Ph4vPOu
Bz6c9bCy4H8E8boQR29u6D0oDfG8rLUFwthZV48Iw2KhcjSuZxDUVobimRctPERfZbnk3DX/0KtA
l7tPbMjylliwm+FCsY4fHN3Qy1EDCsC0fZIlYoLBQR04aPHi0/BYbEgeW0+i+rx+ArLvucuzyDrV
SZDNqt7Ri/70P0kKuBvOpE+OfRBE17+sSkivRlDVBAOgIENXCpfVRYn5dGidl3KZAR3gSQdqqT83
AuaFmOB0tOv5R5sF0mGNmyv2Gleic0iVaWZ8wXx5cvsBOaTLpUAbc5v/dx2HSlNZ9Hmgw/B502Vz
BYn9ze3EW1wFVMKr+Nz4YRKJH1dY6ARG1wSH6Xur8ID2MhpNvbet3vPIGK2rCvyEyibT6hO0yOLe
C3d3p5R5Gi0UwRpAwQgE8QifamA4cO9Tc6wAGn4P66Lx1UUIpj3dOKAiJzgAB/nLP0mwdK7F3RHb
B0XibxOG/0EOrQeY0lmluPOeEW6NcBynPRCl7ACRyfn28uNai0ZvjU8KVql6xYD+XfTrr4DN173S
3MwTpKg8/VP8/9IwVE2xfFThPlzX2cFgsAvZTwR2CeWA1UL5mkUMymmUtnA14tg3sFuKgOyPgQLF
9rrZlZuQJjREmHTb7O3iSQylpUegCbEHZStE+xm+Z7BH9uWpg3Oy2fL/m44RQjmfgIzJF1eJNe7s
bqqLWyjDPQg12Vyg1nNRpL4XIiB5+2TR6OPSmWAvXRIgNUXxJYPe8DlF07Dmse3wEpOLpKKnoTED
oO+EIJU0yXRxvtwUebDzZ6yw91oKosGAcSxkYJ7xR+OW5Uv151smr3mMKQio0M7WHksuIG+pjTMh
iNyVcFXjIjWQ1naUFS3cMMuPAHOG5oVOop2p6DnkR+EjEvvY3+z3ppZUJxmzJU1CrctQAAUFei79
wJMGYVB1E9vKWAJcpT+MzBqdrBpoks5/k6p9KMrhVwzeFMz0GLqzgWId6+W06YmQp7pPLSm+8woW
3bFfvO2JNWhh/g2CuQujw+31K7w7+rEN7SEcWC2ljO8DEw57c8qkd3Dfnh9cEavf40EfvJsBG3UX
CU0LTqZA1/OHWsNtt6yNtzECoun90e71lkxof2HINxNMELrw7w/F2DzFMisGs3igs/kQuzD+/ylA
tl9+1clJYnPc4LqbDkAJSaTA+sOnMpMYSXmAEjFlqOXnDWnn6VEk0fuNcADakUwjIRaIbzXQFWd/
MV14PyeyJu1n3XtdJeWsH0laEscyxpsUKvOFD/PGHjao/27azdhR0zIAzicLCn0FQN4wsSzgxPD+
CAJqrikdPlaxcQ1AFDmtf6kM6DKO0nYvz1XbAUfEoMMaE9CJJtcEf39ecVUWX03nsN7dnqwcAD5o
E+0uVOTafgGTZBTuEPYWtX6AwTKc8c6UP5dfWfU0M5In7HmemdOVCzMEiiMdfTL8KtND3B0cACGb
NhakSzPX4oXAdcrWVB6hlbmhax0pJ+nL5RggigwPwJmdSNIHDvMi0934EZ/+RFi2V2CRE3K0/25H
uGzhMUuNGnuUXbSz8RCM1EDN6bdANv9TWVzPwOnD37LNWXMjutVWe9Adzq/XrNJEDwZsnllnJUhZ
dZ01cS9daAp7/yc0tqC/htxnMeR1kevtHiv+68N1uakhpS9LeSYXz49Yo0rIaNLqUOJBgSmIMzC2
0kuvDyO/GhjIFbBDuuAMcw1C7Clpc0MIMtuXVdo6VfQC2l+kthWfrdw5PN37h8bYCUSygN50bLsn
y16XCiTaKC28tUN26Plimv0GrfwNCSDNifaAXBmInbxiJz6rXij4kdobO1BEw8V5aDUtaQx5F13e
Q7ZsO2HAW4OU9KK/heiuWvyhj5jEHbsYucyRVVf3V4k9fdmY9XpphnkubfCb6Crwhrvnmh1eIaDq
ua5hO3RNlqgbURk6p+GkMN4NthhqWAvmUy33gp+zDRWrI2mj2PI8AVeQRhN5knE+1CFLtaGNttgw
AjL1EDZs/FEmEwPZQD53xitB7kptHEjRyfLoC2YW2/mfsGVCRnTZ0h9Xc9h/5hwvXD7uk0tHSXMq
JQVyk3wK6gTZuaLxuzPg+t6xdsdKjufkh2amaRn318ruoZQhzUvkD7hbkmhXeRyIj7ziDL1PSeuS
eeWswn1Od2MMMkQpdkCqSDq7ROPBvbo+SmleMN/ksXX6TPypYyNC7x/pf9HBxsexnRU8SDS843xt
JUxqssL+/YHpUNkKU3lexZ91Uxh7egWJFi55BbrPVrVjvAAXJ03ekEHxqUQCpS8moh5ANvheayB3
Vny5X1oY1mdifOurO17UbwZW/ObHcbt+bQZSwPjWjVU4QnjxE61vZ+dFe8VBG5Q8Kx9x4UWzH/t6
ZOP/6la85KzF0gSq93IYZhxLirpVamT0eDX0Gz+IgcyWf/TCcZtzmzbSOpeX+wPquLEvyMbz3RkY
TUywyTWz2fLJh1sZy7iNGPIZTqI0ntf7ORhi1+r+dTD7EOPHnyqHt0V46qIYkpFRsPyMv9oMmPY2
Z/RmQatGA/AyREyg4iiPEN6g4lvS+To662SAVrEo2wK4VxJAIta7pDfgy1QPLxlRWKOBEaIjk68T
uq0SV6mfSwWEe/IO1+LZ5eKoJFal0lBMuuCKtIoGM+84/dPbjSCCO/4gWXifxbvhbfTxvu+/G0jz
OWV9+b3qJLrHjZf+s7iE1ux6GoueziFsGDNC2ibc1FJww8ywJq0Z4r2+OgHEdTtgFsdlU3MohZXj
PdMRN4FCw5soDHUTFKz8e3wi4OXHBJq84F3uv3NMKZdIjZOPYIlDju1Y1bjPog1oVfMGFP3fvKBz
CgF6Vtqe2YBVxgPT0ekAy6sqAXcP+QIwuh7iin21jvcp8Bq5k+6W4K6vkWDwtJYDfJ+9yL/JZcqY
hJepW/2IRmrqtVHN/UaNOW2bYFWVzjCsGWIJYlCCfdfCqCg62TJ0WC5FgdVxkqwiJlhMg2WGePJb
e0S2xkBoYXKc2KfKNsN0Bcra5UAKdtNUgUasulc1Y7gCp15Kh/IfcTin0CnV2pPxNj1210uqNv/h
0n9+cGrmU1S8p4Ee6+94SvSYEXki0OeA7Yx3zzyBLmIiSXRJem/2mPhq2JbKh6rR5MD3BQM48NkP
a+0+cy/0KVHFTJBtSPgRTV8AQ/LckmIMX8JLxzgpAOkhHCEZDvhI/8ME5FoqXKq4eu5ZlZnJ2PY9
Ak8XvfUOSYLPw7Qr1PnZvAYQtgR4fpZQMYPVWrpr7OY4B9A+ai2Z4bAt41DiOf8HbZ2pVYtFMO8T
iwJxcOZ8R5s3p+Qwfrp2KNvSfA/dst4NneKTK/AuBu2AV/NmyeYdCL48HFTRXBuVbIm0alWiCcQs
Yy4xESiA9xewit6ylKZTDnxq9MD45bWi3IXekNdYd1Ns9/V2EyWzRsAn/bQoPHaadg8ABjiR+yRY
lVsYcHmHNLfvggIjZ1Dssg161wllaa+2kYzKFNe6LCrP4m+psvXYLTOQ6DIZvChQ5uLNfms0fSx9
2myfd+ff7k5MhNHm4wvBrExzwWDQT1XV80lRGaTa7Ek10dP+jKsPEmz6pudr+De97D9ABO7tlDRC
6r5Uk+OV6Z2vas9d++N3gomh+tEwVyh8ty71ZgVSt/UK18H4jGpH5dmYBp5RXdsPgIkSYxdt8cLY
JZBouL8gmOFY5YLF65pjFvnGSk9alJ3g82pIIgiOfMSOhrTWYRrw6VPCjKwGw9D0fYpf1FC9t8MS
j3WOgjnhRTLbAzxqTcUacUuhU7dNkeh7j+aoE73WiiPJ5kzH9kFNaoCDLoPIVsHlKYTMgt6PTZYy
tOOjy44Sc8f2cESzsycsO1vpfnFUfFItRbdVCNfGssFHLeGx9ZZvjBb3bDdFHUeAxVChU0r5iJYF
LV6tk6XJY1fxmCB3qC6iB/7DNUl/B3kVVYeRd95P/MrsXpuwtD8NMXPAs43TnJxK4p9PwqC2cTcM
htSN6/B7J8cNrv/yTQZyS9MSMN+RIgyAppPPIONEl+1UQL3oAHjMWZQyjzxEv8GmvXCLVKpMVxtQ
tCULs/0mnjSLcgRKh+iLdmlMXwlXz3izaqmtorNMErJNALJKKXpuMAG9FSTn5M5xnJJdWM7ujMkw
ZpN+a2r6UYMaSuwSmfDD5bf9PndNcnA6n8Horte6p6zUBB+J1O4xi3Xn/JBDCHDjYb66BUsTK1wO
6cMWD6Qr/mRLr3DzCEb0uMHg4B29w3C5KxwoU+mMvBuPq5ZM8YnYbHCYKC7hFe/C4Mi0F2ZJfrrN
XnREoI5wVxgyKkeBaphl/hEkXUQKyBNbJ8FmGy5WmvP5+1TO7v+5yBy2ISEIas9Oeeo3v0LFp9vE
ztxW4FsEpo1pLicrhGqZu0+pOsB2vbqKw+5VV9w6w/ChbqjFdH82k9qNijQ2U/1+lxNm2/R0pClO
j+Ibtq1C6w/7EUt8grN/MvcjfZmHBe2y7gatpRe1J9b8rYtV3zWEh+kiPV7SPvehN+crf5cNvfiG
FN35p2Y4AUVahR7wv7CSzOCxBfo/WT9700tRG9qKOeCrB9Opw4Nlf0ZPo2qIqnGPSHYWri23JIG6
E7Y4LThs1+K+wGqBu3o3u8E6k5DlWHbyXAlfXQgFJpF7ygDt51q7zNhr+/5Jk5lr4iFZKTbQzaXJ
tamidaxry/KFbIUqgj+hnU+3PjZ7W9BoiFPp47DzBfNNTTEwiwmxFWwPHgPvR5B33phREK1SRIrU
VF+VKWUFKq3bkJyw3Pb7fqE0U+zLKBpI6nTm1PooHVLVNS1PjSOVwFiAfAqweU8WkYrIrdGroH2o
75RY3pIndp0Gk/MuM89laGBtJOZXWDXNUunefQdpUbYVMflSOrLf0auVSCbFq+VmRJbHEUGg/NRv
zXltObn1FABfQ4sKn+qFqqLuYqDkJ/nzZh+fYGdpXGUZ7lTAB4GnN6+sRLVuVHKey3L4aCHpmMws
vZpK8dCwss/PDVh2wvbGIMRPx8JMIb8thFtdNi1FOVuxEnU/4LbQhTGRCEGrKo6O2YdKtm6A6GNd
93TOsa2lu1qvogKJ8sU3kAWnZmBa+Vj90uw9cuH9BwD7AGaEC94Fhc4dqOhQTYl3r7/kZJ11nSuo
F5QnVDS2dEUoHor+HRvwmbhogfwN6h86QRfNV2s1urIpyFiesVdCkJEeUemnT/9yNAjfjGC/uoOU
osqgL3jvYmunANtFK06joRNMePypYfdVccONOcLcOxT21c7wyjV6iqd1D0CQt1YUuORtwGk9btvt
L5NgGAAUK1D5gDnx9aG2XJelpPj5nnvgL22GB3TLTWwxoGgpJJ/MMu9+0Xy1snDBctX487Yy76lQ
9xlyZoN5+ZZ2uZfE47AuqyyZI459g4MZkfLsRhI+vbVZgWAb4i4uFgHv6BS+RKHNNQAkkosOM45Y
Tp682HsglwGRiBDrf6GLcbxjVrOfdW8SxVh+bThVZAr+yW9jmf3S/TgdDhaOKGqaEDvTg9V2GjPF
ZxSkRqQ6doGIjbVrTyAXXxldOtvZFAeUArnzFFXn4qWd50y17hefVL+l/i0hTkKTfui2ZL407pDV
F39JSX6PuE+VKVW4CgbgPRnC/oRdXuprR1/g7YgYuaV0jO3vQliCe1ZKVWlHKW+Q2pxpv3TX2FII
1I7qMIiD4ZgJcD4TjaVAAZI9SuiR25ZvtV0JzRahtZMTq/p4jY4HVutzt2AW4a3gYZSdJaylyYEY
OMAKwFp2tjcJ9cL/omZ9+tVE2WCZpTbZqAMxCmg90mCbZS3fsmz7cs37LDPZpV7BqlAfloctxpyh
uehTvAIKsPc0Q3hA4mR5EFy2+b+0ZnpHOcnDJTTYUUzFjJ+4/JNuWanY03Ys/lHlPr3MML0P9GHE
az7DDLIR2a1ufar9KpjAMjqtT9TiNN4xddF1z7di7pCOP6dV18FTbbXFczdfxeXTRzs2nvVJKMfi
CT4HqB2zJop/RwlHYoXTxRos0tdxwrbxvDATle9ZLj7boNAbR38Q9ZUUeWkD6gC4i2310dU5E6p0
3kKNFL3KStLtRlXqBRQzYhurap63AP8svY+sAQ28sg8xtxmOuurPwpEX2HnudaNYmKdiQV+xuiJf
KYvmwYT+bdxLiOm9hmGrRJ+5VDuz/imatQviPhGAOcSW9p6DL1qBXknWZX5af8aOpkVdelrUi3xZ
yzqQu9xGKvFYXwXZNhkn0BEcON7vFyCW4AL+qVvtBzMiOJU73CAXun0hnNGgVmZChKbIa6jPEyyB
L9YInUvNUwtHm/KXLaD5ZVv0ux82j49p7njjZqM5/JuoruQDosCOJigsWUukrEx2CQ36IFeVoT9e
kf2aVx2uwGSwr/MBCbkB7vXte8x9aNfDbsLY1H3VExp9//AWvALbwgCpr7f4btg7TZsclVNn+yCv
LGWMu4LiaTFBjgvYwT1I/y5KaXxy6odKB08DmCL4AUQXv9Crtoc1xBXCNAeFWJ54QjkY8HAExYb3
NsTzVuT103fmOk6cYrC7CUZYUEhWiPYMBTS+6icW+LnX91HNfZH9F5yayMyNNLGu2jJw84CmBmbY
LKVaIMbSlMzN3Y9JWFygBYvxZVLS23K3pblls9beUZP9cZSZAkDPG5MwjpwkJRAv0aFwHsIAx+zi
BieCHuTCC49XGaRtUnWqqBv2gSmD6QoJLUGdF3dZLMCZ9nKjAiQCh8qp+ME4GcaOQecSD8xjGvGt
dP8K/RlTR4SPQTMeIKw9PB9JTDcNW7qRzP1dTOZozbcjpj2XXIvI89yFNaJIpk8Yj9yweI/yV0Nm
d0OoIPiZ4UHhoU8fe7pJLP9XZLIg0PjKfQ8z3smJVEYUe4zk1iZgyvgTUdYDCyBPd/Wur5Kx3Zc7
0y0cYHuxBM+E4VvRcn7aM9M+gqAePuJppHvczon6qkTt+YMA98KZvDtWutTcwGfOPkYWNEYEhHjT
uFTk6jIdcdv/OcsQ8Bd7kmRZ5ABg8TGLOfotwAZ7WWZFa1KtWOtPViJPp95A4/RPVG2fSBYn+QPa
PIvhsEp9hvgPHoTWI9LkAn+cfXY9neYxILCkyr+puUNHWN+BnQ/NW1Xg/vNlPVF6IBa53Kj84XYY
VF4g46QcweniKUo8gaStEBM9yeKFaiETcAS2T9Qe+ozJAhHIITufiIRVt1nF2ntCPr0x9KjO4vBC
4fO6YH74Cbf3pN6TtOr3Fec6r9qfs9mZVzyjd5pdNUa5H2CKPrQaTo0/bUPbJcRCFddg+5Hu6OlM
1JC7Fkiv8UVhvc4zQl/HkEMGNRsBiCzVnMb6THQCXfo4rX8vFjVraC2exY3EAj72XtVjhv62g51F
s5MqRyKC5O/JdxIsbAUr1bqD8GnX9rabTq6rb01tKp7jclFKP2700Tu0XQ2EKq12ARfIcJGN5jdI
K10cZe+on58J6D2ZjCEpdRRWsIOi0GTdNlQeP8ChUBuHmM6asEHG2Pnj3O5A1FEVpNmp3OSA9oLB
cSSuTWtfrR9RUICbfMHDdp3NvC1Q4O4xHY1wrYV9kXPjatdROiPF51HHV1KgeGNrZ8cRe8J/pN3Z
0w5H0FXVwGe4Wrr07zSzKka6albjLjaVrLJdWP7tqqU/WBAlAavyUzSnZS7ww6UgLlQYr6EMu1Ye
cNVounG0lBzUfHazFXxWkOinSmYRd6hgJ4YUjorVAvYX+SvinQfJPkcuGHIvir3TT3xM5B4SzfoS
17DGqvxg0y6pnbPCx9L/QqR03RNLVmGkyJ6TZ/ES6wgvrapvJ1dOV53m02dg5zQgaMxJaAqv0bgL
z9Z9aiDV4N+kCbGXs9N+kLG0OwsWKVG8ZWd63XlYA2PUB7oXkpSeiMNLv7RQafvjFftjqtlpY0wT
FaRvqFZQ80oe3pwpae5VcsU2xiEwMyNYxNrSyMhpHpgNi9pN57B/LAWfvcJm9CQ3FbQ3vazrDXVy
hYqcUmq8nbisMVhuT44sN4aYc4tRzYKfH/c3Tn5yno8F/JpCsdS1qma3c/yZ7TxLJj2gTEQySZQA
XBLbAO56oUx92XsCC/zpXx8wcj0kZMPN8+/Mcqr1WwtmJ1d4lE5xFLLsQVpzbySTbnDufKd/u4QA
ErjRlTNCwssCOncHJO8RjNKS3eg1tu/gmjKurgfg+mNhHJREgtfCI2h0Fw51gY9qPBXje6VVWmFN
+TCwcS1QgrSeIdQszI+k8fxbdMpINsD352+VSR6WxxsApocoi+5h/Eb7VFKeuvJn/JavH/NHFHnJ
GPE5pjx2tg/8h0Ty17FlO/dKikyVqnzO1PaHizpmYpXLebpBl+4JmKfydEWIM08tnjobaCM6buNx
StSomFVLRxumVtckSgw1pYi0+50G5QEGjDtqv2GlJbV/ofUq3GHc2T+D/yhsuao4upv69MgoTsR5
HWV6aYIZJ2v19k4qdVsmQepdHo3yrZO4BkTbmsxowzEKet4Z1WMBViu4x1k+gagHOKd/6RPE+ZM8
BbkdfAalTvX40xedRczChtrh43eiiqDxdBIzdj8s74aQ7T9aPJFV7gqwloJHCBfD9TFIDrI0Y4G5
76M6FwG+eoA5bC1lGYQpGgpFBnqN3MJO1HDI4zkEgwThQzJCOmbqM0IZxt2LNX0L2JfoCfB8OURS
gNLCJgf2HLnRYmzGb0o80JBEkf9Hc0tHufVhXB2TjY4FEKA90tb76JmBKazTdg+Fhu0DIl9KGYeQ
M7iMUaNaQRlzrFvWY8oPWgd39GenObi2j7vaRbNo88AQUqbWJl4hVjiqlsSf94Hq6E1TNMkZWY+i
8HW/clZXN6QLc1YTtOk8N+A/9gFqv5zqNl/q4d6Q7UNznkaduXS7t1fTmFJYOFzXxWG54h/5Yaa2
ZNNYgDg5Hjt9oxTxalQ6pAVDQzMKgJTQnd8BfwjDY3ByEkeX3cCjBVuMvTnF4mLIHujXyE1FWFxs
Gn1DkU28Q5gVLP+g4+zS5m9xvEKNtQqwkG63uj2f/wfOsFsF3mA9Jdnadja5j7KpQ5dhUufhHrkd
kc5cukEaOQckVdyFbIqShhTWcWatCGZ49G4VgHgk24sf+wEki+4WXh22gLP6stZO8rTO6U/q1V25
4KxgCR6x+ItlFXB38509XRgwCOsNvXj+/dzvfGHsQp/Br/wEUpDRmy6MEj/YaYzo2mfHD7/CdnpI
bguBsGbOcKqra4hw+TUSlBurIS7ehSzXRQ9ceZcOW7KE6EkHPBkANmkFUkKQ9dTLrumc7k9Y+ftT
lgfnwOFl5Y9qwHbSNVuYdqz7mhcZZUVq9KKPBKPh5yS6M0n+f0gA3ztVTI79E4ZmK7xn4NFfw2+w
XRjwqxXsxXMyGcgZTOcOqG+L/OQ8v3G11UmJwcFmDRo/eladDln7mlbf9bszPp0BXypRIIEkFg0t
odp2Yo+EufHX/BRrqFBs9BvLITaLt5AtmASHQGNIq7Rs7a/T/bbByGo+oyqHvgOn1gIZFRoBcNnL
+tW9QIX2sAiLl1UwGxOOnhHsCSCJE+XTwvUB+kRyn1sJlwTP0rcZ1wgtU4WdsI9IbyikGyg9TSV+
QYuC8YYRnMv3KG4qJ14Amnu9V1LU/vdv7usJ+01SKW/53K4QsgoG7Ci3sDDQPWnn10qtE7lFF/PG
yE0C82xiFdvtDbfVTb9vl3I2asd6mBVh7zAAGXWR4wNgINYkyBAnfAfbrEEHqcIeLaICiCmaAzta
gQ8N6QqvTe9VyC4r8hg9diPGScwdFcrl/S/P0sGBb/SG6S5heGweNWBePL3E25ruh+fJrcVroEx9
oeryiipBNvJ6y7qaW6MTtOnck8XlTZLg2QVz7/f9AKFQX12XlTZvBL5DVUZ8+KSHeZ2AZB4YHFfc
Cg9bJo3wXJe2PIdiGfJzi8yzUtDkneB3g/Y+/Vqr2hfjvV6SKxEYzDERZpfRYf+N8YHwx9O0fSH3
Caak34DF1M+BrUFWE05bNd7eK3Sg+pxYC+ACQSiMXkZHQg617HMZyk081GtZSB46VsTjNYCCy47g
a5Vjt1pGZHHyYKLnDQobPw2Z+5nbxWjambUl7AxHt+hEhhfeRA7FmluDz5f6Bmxt0Pev06w/9N5H
OtJmpGHnBVhlEUJczS7Qe2eVJuqJ7zPWyABII8g7MyZad3XWsUmLfAt4Rjep3HfWPipwIBERVLyC
2lWZgQu0XIIFmlB9p4RgSYbU4orhj+UEignR5tdi/q/9s6ck2g7hgUEykAUf7NcA+hiXy/dmiPvW
yBP6OpjYPz69Lx3LbChxErjRdYsCo8uzd+RwZplpBDCBtzcpF2xvY86S5yKN8CTenTG9xfpza9OF
4noKz0HUjRQCJNroWGFlsB4EOVld4Art29iVoshuMDgg4hnqD6DY+QphrIq98AFCL5pZBIG2X8ju
KREnvPxyOioj7bkA6S1Ru6YEaw6sFIFaOWT6aqZTIexUVZTHQshx0i4dzrpT4jMoE70vlIWMMUap
Ubsmu//K4ig0dxj9Has6grsZXLCdvsz04xHvu+3hnh65AEqglOMqBe1UE5un2Bb99MtuMxDWhjR7
6DsFE6/Tnrwx0xvyacPPMvMZo1C62Bfme/e3iQr+9pwPAPKhiQOCNxrSGO5G7L8fXd7DiG7y/SXe
j3fP7Y1giYxHpyi5KZwEsfQpD7sGq9W8uTgtdYXUYASrqunPinA8jJ9TgnOjxl0X/QSdK/zNYkNN
ZXpsMwVaixc2Zcay+rng2EDYMsVlx4rwcU76A/OGkVRiqqEIVbD9HuSU+kdKuo4kIX7njZHZnzi/
cKx/l6W7CuIdfN7Au+ES+872zN4kHSPwjOxUO8nQiYIa270oWxFl+Eze7iFXKqE0XKr3qhVYsqm+
F0XYh8RsCRVRK2JizGPreBlMycjbjslTEVLtRVguWMBCbwbyWQXcdcAsk01vbA1ilAwnh9tBpB5b
rHcai2vQ0oVKJ8qKFVXvdo9XCjq99eO7yw1PNXWbXggwbtVOuIvXZAl3AU41AemOoLxvosRzgvbY
/0vmb/CAd2vI4UEBPTEZJnYMqYphxReOg9Klfsg9CqaavAFlzldAgrXY6xZ8zixqXN5ApOsUoWfd
kvan0Z/oj+/ZDICNCH7YxddDa5hLAGpX23JRUQkZVARXb3lMakphBay8rXbfPQHOPA3Zs6icIzPt
aNjYhici0tA8O51kSf/vNw+cOnLC35Ua0azcIaCZrcA/0ok1l57EAgM5J0iduteuZJqwun7NCK2j
x5JjorIMaREafb2NBuxMqIoP1z/yb+gw9Ubo1hRvm6mtjhM/OGGMfNNALyNatRaJCOaF7k86FeqC
xeW7DVId1i+wlu66kP/D5fZaRH3pv6Z8SfVywt4ykBE9bPrOTISGVmeB9aUp/lrNyOSNpal3RBwF
OdH7nEsee0YSjkBKEToCbFAfp8lMcscvVl7ck0UVglUIAtxFO2gME73AvteO7QoySUvJFP/qjG3S
YNq0xlCgWMIfKp1GYzYMdTvV6LEveJva1L6f6ltCprgWzDKs7SOZh1j4zFwP650NJUxF4iEYxY6W
QcxatAZ1iPsj4bVS2Io3YhcdGuc1cEBBPs0Q/YrZqDNpYtAo2khv6L3CqK2ejwEJXSQtoCS+UYyE
0fLKYtB2W2UpVLVjkgnTZVSDEM/PxWOCe8oNscTRsEd08qTt1SyGc5M7oF6beFr5Da55QKi+LMdZ
/i1gMxTCwsrdBqBkd+ma4Zf9eOY8nkEhvtVJ1Ay5PXDwolQ3Jh2o/Xe7PPjHGwL8CKyiF/YgfQoE
zkj929A30x2rMW40JgVaRc2zRyp5DvVrsc7SgwU2LkzP97FIu6UwfGxnBkuEBkD1SkZnL3PX2MWT
ODscR2ticzWTQVRRRD/nckRPlkFfWWj6eWZ46nBk1WP+8vsMn+NyysFhIfGMHU0R8uUNia21LPh0
RMl6hGGsivtxP7el7VVVUgpLGM6F939h2TrNK7MjRsKcOZk9DbbYdMi210AkG3qNy7kmUdwLZk/E
ohiKO7jz/earfLp6MwKqygfI+2qA67vNqmjGLY2j2NU3cxVRgWJ+df2GOR2ZJ7g4QP1r8iB4mYjC
TcefxFrewLJ5AGyEzDvw21FYi9ANjNETr2B2Ius5W+EzBVevbhjfaZ1fNcRfqpebozKad50vGiR0
ZZ2p7n3VVOndcIxciiNJwKPavigECXFQB9hP/Q3xAGIcAj5Ajyajym+1Kc7HNTCLdZEpjiQf37pp
khkrNMLp+gpkt1s0f62btZCJYbY1fZZhrPl5zTx4VFm34q9t0KyXkyQwOMW2TmzoxkrbtgvQw0YY
+SflA7XuXquKUDLCqJVz75u/E6YbVbrTiomGnXoiZbqLZLQNHBEwJDEFvlZ6j/rXbjxaGCBBT+X2
LijybBGkBNRL+maUDi3UBz27s3/3ODTmQhN3kYjG2twHiE3E4s4xOX36Td0JiBEeRrOZqpHIwXtQ
Kt9oeSda2IyA/6C2vRA78cqnwthRGCs/JZ+mCxg9dVdJhnNM3zndxXRRkwLXYIG9NZdoJdPit+MT
OCaoLuJ/ch7x69PKPU2G6cf0kFAE9DDr+vXYRByPo+GlG7VOk/3gfy7clPod9uTlOtP7a+bH3jwM
HRBnfWuNlfgEfQhqaNp0pi1Isto87n4s91fjfC9ikNQ3o0ajDFOpZz6lPX1nhvJs+QNp3Qf5zFIA
6CaXH+Pb5lE7tgOYYobMLw8tvjN+L1TDl5HEXmIhr3NdN/XpNlq1BEEIzcyEMRHbxqXBJ6ajJYg/
zDXugd1xIObyfvwuiGJAfeAybpVIjxmpGgB/THbuGZjnsBX3KrlY+Gy/zNvzyeg9+nRKv4ZtGxLx
KnmMphGsTPsSjwWZkpX5QZZ2SUAKQuK9mqxsppDWkRF4fR3027AV9fm8kyM7YDap4+d7qCa6zikj
7RC7nCSTGSiPnALZy3KrOv+xQPwCtgu0frMi7GemLy6SCG6ASQdDMOSSgSazhgsPd0eoIJPDwvYH
uXS6MY8atfV72ozvSF1iGzfT4ijceWN2/jzeQFbBOYG5gqplC+NQwoCY5dYlnS2Z4SD0Ekanhvlm
oe+glzxr86BaBDxPq17KfJM4441fZzeLgrzCEUmjfCyALZdBYDYdcZuLvS4fYEjZU/s++pdfs2AL
eBOB875MyvmF2Xqcq3y2erOgxZQm5kAD6M8dcsa6gay0DDma+MUj4hWTnxfnhpXXxbluMFIBGo1v
kVdDJLP52GRd/eiBEBJkXlhqu+gsogcYmM2Zqf+Ojvcw3CBoT1xUntUosBNXGIJ/J1pnJP57ouLa
LJEPZdOH8bKntPUFu69RHS8iKLprfiLXp5WqnFOxtCMXi5LdqCHcM5bcqRGmoQxIeY2dDDGeRVsg
hIfSjzR/U/0f5zUxx5zREpptVXaNFmgYjkA6/ElhsOXA92S3bIUNO6W62WAiP030UA69J8KrJQC9
8z1EYMI9Sqt6WkDqecehlLiM2+W3sbOBLsSZTLNna/DHAxbR9zyuIneKY3FiZGHkRinYykFLW4gw
MnoUZcbE+OJgXajpgqJfY7bVQTg4/vvTe399yf6qsY9bXOBp8jwaR6pak0EJllilzrde00f13YWP
6i1G5HkeeNAEjSt94i1stiFeOBpVSdM6HL4p6neNWjEM4LvaKRI7nq7ITBvfrGSe4bIxOXhdFv6F
HRD9iDq7AQ7VpWIBoOe0SGIjrXbditvg7Q2SQDfWsvlCwjZPrkSaa6CAhXdtcobbGO2f86ti1PWZ
PM/D70rXpCzElStjA7fkNEBj1QqCBVCKojwVxZv2F9N5PVjHIQA7qj+JAdzxmfCLKQUcmzCR51SQ
fadgLKFVyoQnToGSS1c16bCDenX7TIQ8D9tWnhpkR50bXgOOtZcHcXFaRmyk2L7fo7wgoaWGbP7B
LVIivO8j93GkDdnyQhG38lkMBOJ1uJbPXevby2yymeq5kC54G19LoCUQ5GS7shmlnv2gJVajV3Jc
hF0KT2H8wMnEFZqx0FsB7HdLEVIabAhEU88zs1ZgzpF+7+zIohnTaI0FcT9PhdId/IJ40iHyG8W5
TONlBGtDEPkAaGaLL9wWHqgvGf3KZP5aSXLQY8PWjN3Xib7/KabFRE/zJSbNctyk1wmkf36sjHhB
xbiaF8rRR7yP6PHKq+8amWQypsS/0UM0fj23m7vQH2k10WQ+NbZC9P0pfPINW+ewyYQIM/1xx98g
qcOkbe0PmyKRHrxoU8R9Fai+etr9XVLwQUUQHBEXN0ChEKtEn4OamJko6zGv+uZQjoknpeD8PwfW
Ylygxyx2VKkMriOU22340r1kLYAE68zbj8cr4dg8MYVdSjSrnqf1L8jY9Mh74R0UlE7BgatVSB7+
W7ypwfDAxc/9Y6oL6/LpViNESPLgldkcvNLjDuwNUph/YpnmsU77fUpg3mWDaOV6yYqVgz9Sa7g1
mM9/jmmApcu2R9rhi6PvE+3ay9pK7VgoosS+5BdejVQ7zcPcS+UPhTRd3+Eu9pna/Fd3tchvxm7e
vIAasHRi5uhZEz4JVOi1Gwb+PStUivh7tT508WZic230/zHDBeSsFyeVaWQm2NtzFh5YzaKxVC73
xYISjNs9xuVS2JZcq96dybyKM0+NXGvgOpG5Go/VOm5GbRMPMJIfM5Zc0nm7JeoK8INVPxne8eeX
t0RgfUutd7rYGG8Fp6cHucoqeGHc1Ty3JXWQKZkcDWHclJOXQs6raDABRy6iSfpBd2eLX6ndA/Yn
jRlK5yArRsL/9ZCCBrgdFSgoxn6ZyYT8q+1Vz9LKdmWE+4DcGdXPbXocnc0aY3bcIKcqpBu4Pevt
CHayPqtPZ0AlsWdyQh7Y+XEH4XYoQvCpuzCDaHvGynmfCM7tXWZMuYvGmF4uj+zn7S7QK4ELaP/6
XKrlbCzbe1ZioSyAWzEQQ1Tmq/BVD6kU8EjzsNv0ESwS8Z7LookOK+Z69fDVgjmLTDV45veU81st
5HOYmRTJH+SMW5rSVw9nux5zlg1yEL3isLCuaI9WoLZUUSvpYieVOGum9creQVb5rW9KWfva6MTO
g+Hu96jRidk5Oj+xt70C6PNiZZ/733ewQnQn/JEu+CRj8EMkL+XRCme5i6XQFn6ADEJbFN6aEK7N
NM4x4PG8+3WCohLBV09epZ+shTDPbbooyf1MmqHDBKRi3DU9dNKrVfeMN5l09e6K9nPym0kk4DL5
ZGNjxALkik/6ZGPhnUiIffC6gdUxugaZhYnb0Usp220giuL4xd2w65kUub79jkVQtnEn6K2W7lsv
5VAHDTIdJ0a47dx5Dfdj2NYks2Tyf53rWNMoifSW4uaVKzWtgExLKbBv0j9Udn7A581x6m5hBgTW
184b9imv5Zn8KI4jZ2OfKe0npVxM9jQgoHPDGtGRy+7dWBCcsuvs5B7uJSsvqDESNays3oXPDST2
tovhfI+dQMfVO+4D8mVe3zE7Oymhj2AYEC6KuOPOac/5vx8xB99PH8TOkEaYX/1J+2d5911GZWbR
TkmyfSj6fxP6ZKShE24iG2aQLoytMyM51r0tZYqux52n8aDkuahux3b/mUYS6V/FsZ/abFAp8CQT
HzfCApjOB8/MPt8aOIJOweRaZ/YUQNkyhYtyqzVOMKIedJa0wes0mVU/KuNK4iibUwbuVAXDbRxb
RUXa0b3hcYwKXKa8Q2Ruc4CjuLh79/lXEWdSJqUinSMMMUbkLE4oxGL5p00RGfZxoWKtbr8zYmG5
mFGu8ykO1F/x2ndPsW3/PTo3U4O0ln+prElSwVnWZSi5UK/FJaQGRVIXHNy2Owaw17mC4TQbz/Fi
7ZLxtekiS4yIZAsvrbbMhtHgDMAyG3gNU736b8sUAn+z/CK5lTC7iz6PDrwiOUaIypdQPvn7UY2H
gCtyczi9cjAKjON2Xo2tY3duvv6lC7K2WD/h+lMaOkPJqo8/tLWKxzYajBdM6Cjs7cGf1q3dahUo
b8OCCSXAezcjFRb1K7KRvi4zhK7DCPNcZwGrv/YOR8dPH126BdEe5eYCueeugfIlH60n91s3VKIB
fclCYHNjcmG6BYsCaYAxBTiEOGkhVOX3Shqb09+PAcDfXftNjvB2K9RLmCYe43P5VOmvYaZhwkTB
GzWpG4msReBwmYVZ4sA63liwyuCSndaFbJ0HiRIxEBUnXBZUCRfIACe2jh6Y5amxM3H3ST8tnOwz
wa8JKeHReNs+NgA9LVWTW1nGYzMD8vdwaVGZBceTrOyel54AYv5JgYwkA0/231Uydw/JZyLKofKt
o9BFgM2AR9iyiyi2lxegmyUZUBUTVeuFF2pU0xOpbEsUpV8j7xOgwilUwW+sJDdfK/4zDFDiyqp/
S84X79pKhsd/gFtpT1wS9W/vdpFLvdNRTB16bgpLrIiN9Tjcszy9QV04kfknd9EeOUgtcBUQcCps
MVqY4yquRby+m8jaTVaalqUqVMjQIsE0WNu7RO44bAEGPLA+4Wh74zIsxMj48BsO9bNI4UIK76dv
reD+J3KGdHuh5rve/HK1G9zEhN+3wKp0q4qgL/PZ1feydzQKZ1HT+groPbmKFmiYl0iBJr/zysrM
YalcSpoVazfGtd1H4K4h0h7FLQa4mFr1mXrWzamup9Nk0JHVHbEXs400baNyzfaM1+mAnfJQVfbL
1R2utKI/bPiw/P/hzml1z+17YFqP9E7LAusWPlGPJF40rnOXLshPAiHSKo8WVqxnuW+eFJ38vacq
4oZXMx/f7uK18MHMHrPbyLyp/D8NNud4qFM6Wp5ZWTEyvf3p9zEn8uWR2jl8LhLk026RI502Y2jc
N2lH+Hzn5aT0744fSSUatsY7TdI2I5QAhI4fu0bPxyIDrYxL5o+tAiGXhRlCYJ73QMOw3JgcgHZO
3wmxUzlXnZMleLd4db2TZWRh/GTn3ccsO1rZa8Ob/bZMQxykr1fooVLCikmKVO6v9ddxlDEDOD4w
9oEO3TydRLjISatFq3pzk+TKJpuSHjRUjq+0ByZWmPjOKTC7NEEIXmmxh/ozxAUoKHQztVOlpAFZ
YLRUowKjUsrWXo0G2Le2B4FWO3vFIJe/3zC+zBWEnF+pDAg6hi+pfILrTJmYtBZkjBAEZLcao0S0
EprT+5AHGl/3ds7dCVO3aOJbiiV9pSTMjKlW8pwakeYYWQjgEBtFZUYuLCiQNQGLnLhqbtYvgyh+
NDCMPA5GG617HKFqhEfskvTZUcZf71kShbT4rlZFc1e/gGGrwLBNBNhht5fRhmf33RzH6ncvnGwc
xPvZjnelkK7GIQ3uz0gtdea3P02mImQ7iccULU67eAgoctd1AjjyV/3J11fZ6tlEEroHI2moR/Y7
VYXQgoOyF0HrBPvWRBmD4UUtpvHxyLOU+HVyyFNYWVQkDpzIvR2by9Jsy+Ss4Kcc0GP4HeTFfyMR
X8b2YLtr140wTTMV7d+XddPaEw0EDYhFFeqq52ZWmAh6VVoJm1lXknnXnRpqzpX380l4cJy7cWQf
ta5DrICWH9E2/eI19c447uwWJGW1Pux4oVontfAyyj6eSqxBQtVzeOd/ADKtW80C/H3rBnj/2Utw
WBJ++5wsoIkZGoZYJLJ7Ol4ib+rECwe5IE4M7mWa3XZNPkwvpB6cvMLyK5FURy4O1Rejhz+zLtaf
NcojuT9ZEjN/Bs/SLikhN1pt0vjcQe178sHWH765CddRkiJEma5999fnDyQ0iNHK2G/tvIezRe2+
iHtGa0fkryg7NP/z7W4t3GcUsjuch1/TZOOLTmD2eCZ7NQ5UjYI3V6D4XBuGXCoIh4nN94Dq6sst
XZqQWvgV0RZfcePtRaDRt4hkv7UApxjSGhoTOUeKWRG5lcMQhlZAvJQKTmsNjxMO81v10VCkgYXN
sqETO9seDVrA2FfVRCueDEvJgLU9Db8c962iDWgyPoPuVKJvyIDqOTAaGi3wSeGv3dHS69BJ/TQO
D7Qd+NQHlGnikMFKkaxAml8vQ+aBji0utGvY5QqAwQDmN9jPig2e2JqvdSzUhpXhAdVPin8aCpTc
s5xqz5GL43A5cwZIw2V3tQ0rWbeePV2P+5jQyYrP1LH3+v9kneKr5vqPk0W5Lv19vMKxQ9QJCNrJ
AbNY5Ux343Z6fyJ5NgRGEzNsBZwsW+aNAoS7OPikpuRsmn+CWM3nXp7CkeIIx1aRjyYRQnNjoUD1
dB0lN5jPH9PHTcju8EVYkYC04bC2qmeu1LJOVJAaaCRy/z2Y7WL0V5o4NB3CfnU8JgptUGOW4wU1
nEGMCs19HkTkIvo8kQf34i15viHjfv1hCH4J/he8CI7XoArJYTclTrGdVB1WRfmKtLlGhoPIPYOx
f6RP4O8A10nUIHxFkXn9ujhaRV+gZl08hEpjIDUAnJVClVaPlHOoJUc+Ehe5dwSfUgPE7hv4OJ7k
fLoUgEWM6OPLDUcBcVRZOXyfBVYt0VTyaVqUB8bx43gwGBAnNNaekduQ+EQBEQRmcIn90ppMdsJ2
dbvOBFQXPh4OPsFJW8AE5EVcerKM4bWn+ObuZ0ZO0D/bH+m2fFLIzGa4UMYUVeF6z0NYaC0IU9Ah
T2pEzPObfThRA5QacQECd/bFqeAmPQ8oHZqBB/NFsuV1wgg3K2bUUEVLL1huKTmMDqPYvO527DDY
9Sb9WA2nsrDqGZDr0rqmfv+3vBmwCHAHEGCe79uXGSGXogMAJx+6zbh+X47N79Vg6N70Qj4CCz7q
yqxjmQUHmKc/nHMoGkcaVdi6ZfNQTuDeYJKGApP4rdnBtQsQSANWtF1N0h1H8aLgcnFgyS5kLb3b
Xuany3VM6chh/J+zHnaI6XU1ACzaTvI2N5ZCNKCsT1DKoD/PxUNyKQqc+yXfqukq/zOCa03VcZj1
1VF8aox/Y10yi2w8ba+REASmTd8CwvUypHnmaQHYWSpbPXsH24Yy/fkZ90o88ckQOVSvbSs7NT3f
A2bZ0hDcKXOy2NqHAik9RmNrxGgE44ePphoDC5eiKBp3uAtUYHFg0DlJkHR7EwRE2QDgs8okCDCh
XA2eH3V5TPTQYtJ+qmG2W1oVPb3fqODPD/k1BPrGVyIjLE8057N8hSBljU1Edq0JFuUyf8ooEO/4
SADyszb6RZjpAuXnxkIgVuIAYoOEbze9GXfOfR4oeWRFZyYBHN5mlak+or/nCW9FRlJulGTb23Wy
/ZVtM4//M2SbNQ7OjpTC8fwW4tj52wVDuODZ5T+uLyDcvRqloqlRHr7nWj+iqT8AUdmJG6H72yYo
FLfkJQpNZ4AHqzmBSZJ/jWWgWF7fECvtJmSV4flZRbz9XJsA1nHcYZyaxhduojztolIkdGOUpDQu
C5XKVf5jLPRqWQ2xe+fCa8899pEbtM4mi3OuWCq/8GAKg0TISJhoGzrDtpVCnc9E720/QDh5o/UE
OW7ySej2jymtx7H257u0ULNc1HZY29owjLEF0KoDIHl999OryRtq/AQNrMC5QGeDNQtFeaY5oUdw
YBIcULgGIqohUuAOPYKOh1mEUc/rm3YaH/ZSnXyDmeb24fgAECnIbuEXqwLHwQYsfvG5VvYgsvba
vMAvytHecy5WOqJqCMWpzvhha+Ld4UVipwD1v8nZyzxJJYSeDGtG/57od/ZWWVLs6L5msEEIe1v/
BbDwUOko1b7VC5zFEbRyu+RcGouCjP8jKjgIOq7Cju8xaNB4Tts95+/OJhbUtml0MEXYyHvpOmzF
lGHMJR0x8Une80sn/UO4F9IfhwCnOwKBMsvvUNx9JAfAa187TMspG3KXLDS7kCHhp+gQOQvlbxf7
9R5AZuuq4sFe1VXWEe9nZOmLzJH4tstaKzLz4NstO5cgoIRXKxEFwHHc4h/glICT8ay8AAos/Qt5
UINYE3eU3rhfB7ZvVFM4/4mj8/wjrzf9IbEO2r498iClg8ievrXt4Pub9FAIBz0HQBpIhJ2VgUzU
5bNvhWluwxuV4nuCaGEZVAyfQqRvev35/6FeDaxfXMeJMqt79CkXMwrsDKWwqBlJvUgBgCASUwfI
BW+DnkA1WxSj1oKEtyQ4Tl+BRXRJrQ4XrUUBlZf9stSliFeAZRR7OjDynFW70IAlFf1J2DrNhKXP
uiLhnJve7h2dlAhlZhUr0iovo9nvjfOVGhqQxfxUUtgbL9APwjvUljXde/0DziJ2TfVwU6uCnV4S
soUfId7qRbSPLZOb+YPeu/ti3r2dWRO9kQJl52I1C14VXlazRwoqOnVanGnWsIV40VJRiRtcsR68
DucABBJCkhjFSXOqCYvMV0Nnr5TWjkGrT7jgsRFIecagJxtkAs1qkZsVzhe2LNQC/g1DsuyZhtkS
J02FSpJuXXJ11wximbT32ChMR/rKKR7yp3tqWtmwgXFbQdjUGIDmZuMylXq9jI+XvT3eFN8Ey8p5
Dk4U41VhbZrH+ibH6x2jhiUmhrd/Z7G/qIPgpoQS9kafQWyZ6pekmkQIPQjpct8ioBVgoh8S/Esk
5+4IzEVH3B21/XSRvMGXScxJqJoQl37hqoCa2Oj3aUTHx2ztHts6faIYnvcq07BJ10piHDtpZ3du
Oqk3FsVFuuD+K5PyKgHnpxqA6JAecqr7XKWKByNXssl8O1G5bT4JQlYNaAy9V2QhRro2Dra3g9DD
ulmVx0xvlzrrcPeDOOU15NQpXEuDwmCr75F2JpCjTekWHIXqfofjso7wpCbKrz9uW4YqYYfvrHWH
zEAsRq+puhtAeJRu78UyYv+02K4/HR3dUrjqWW5P5iU4RAH+PB+fZbNK3tPn5FEEgVPhRNvitDSh
zPEwWE+HGsOxqFcD3rqjhDPTxGswlyV1ObqHOVsfSfnMeAKepNFgpvMBDGGU9mfRdz6G7wbvt3fN
vWXd+zg7UblOppmUakSxY9k7TsUzeFGdc3lZFY/A+yUSyeKXAouhbeeMKjL8/0k1vkMbeOdlmRhs
XWUTkVTJkkIo/H2yi0U0jGDsVpUZI1Tv1ZeZ0LUnYA4GYrYX5TWrJFcciZ81pnCKyIrUUocF0RJ5
HqnNDZu/CVOonenWR7uAJvcFKj3o6G4KqOsJaGKidxlMr6NGT3iil4mUYQdUuR6N0gLIf934IRwC
966IsQOQKCagiPT/MdzPn19LXTiNXIjrCAgC6IDKfyLf/kAJaDNExdTnwUX/0u/sXqZUXNqxT4wP
IpwesyP+F4s8KAGAfDkeOIMTGkPVTLJh7jGm1xCMyAmTAkeyAr1QJtklp+Hr4Ta+EYZuF65eFijg
esoSl9qReANLIFYDAUhLXT1VGmaUnHaA0RP84Ut8Vsf5Rg2ZuTWlWL54e/2zoONmIhWFVo1EYFez
s0vsp4glPXMbraDG7eIder+6ew5HJN6jz/N+zdOdD5MqTTkTmX91Wp9il41DAqBNHanuBkC70MMe
2SLJ60DOnRIFazy1w1NKVDqODdRBYq5TfFP74ARmyMmlkmZu5jBqFwKQOw54e2+rrbg/ok1+si6t
HNZUJucqeIQ3IzctL8QZrWKe+Cz+1zHWxyFCz1KJuwG4UDPjVvY3cDmRnTM68eeWk+0VkZC/jeCf
l0CnIHjuL6zpq8OJOxsgiXWzEP3Txt5UgvhagUguJHVg8im9M0/qIJd6aKVTGuJ2YyhT7UYPyMfj
spt11EpS09/cn5Ij/WbG8u3J513hm7Nvjo9DVU7mTANQbyZo19Ve7titpL8Nwd35DOWtIjYvKAcz
BzDlSD7mjRsfF9z3cmOn78Wb/Y/pfwkynI9rqdMUgkVyuoRd8NqYTIkjyrcu/4LYes6HQyo0AEl9
R1+5FpirT6lQHZKpZx7Gj8uS0w6nFroWzdTDzVUdvACdrbxz/qJiWfrxeijCagdrkdBZiFsQpREY
Zucp+AIcXmAu5j6T8eh9fOsuzQfvG++2dSiCWvJxxJZAygE9ROmfK+ms8TH6dj/EFJ1KSSNXX+up
GN7TifZkbq9p3XUTAZgxQzWMhX+DQfVRlwHNxydXDeNpeLS9OL1h9AOlvbVloT419hd1IMabqJ5B
MkI18927VvyfOtlUZjHYfy69VCvrEZOskjtZb5IAFKI2gnDhoepr3SGFQPeqI5v3zmpnRZieOMh0
oXBYfpdEiEofOgwiNAhotx6prK6Q7e9W6eQFdgMZZxA9LxxxuZ9W1afKclTS6+o+809FmSWtB5mz
QItM1iIFVZ6bo1CpT43MGQUMAwvBhjW8CRpKpaqrcPNc+Bx2ht1vNHQMhmXbH/7GaXI7TXEvBnB4
rBpTRVQ7tsrVf3RU8y1n2UpEUUGUkJf/lDM8liTMnbUGX08UdY4KgJNuDvBNaK56aziuxtHUb+c2
QvFUIhr7ICY6lwjXlIEv6QtFn6CaEDOu3GklYaziJ10TNa1fZxrhRMiOreZLOH/scKtYkqNTzaWc
ZAO8jVhN+K/YMNppJNRKqUaATtRGIWtp96OPZYPQvMaYX9n9Z2Gl5u6Naf415VVhG2uxDoMMKlQ/
WTc4RY/W/QzH5CjRDN2I9fslUfYhFu81BKal8+snc9EioVEbQNX/Yg1QllrC52Riez4rqrqn0c9a
1fxwo9bVhu3nl1toFzCpCroVp0YYBa0ijXQRtgrGAfPpm+VEh/SJMOH98JMQ5pwWQ4C+K2yHZeos
K3HfAK1vUJBw6xV4DJfW/ETntmetoA6VTHYb7YC/vui++JONCK98APo5bA7+5GRjGwtx1Bxl6A9/
PAmWHYWRT20qoC/M3QyzlfmyG+Q7PxRO2dVDurl6T+InsiEp/cr2frH45E/GGI01U0uWdERrD+HO
Pzuon956kgzHtrS9g4JOO5po6VXA3J1U5ePgvO6fpYrpM8WtQM/LYg0IYo0nj8Q9O5i0Us4xxVri
mrB9z5IRpIGYgKJtvZbWcWqb68vY+ey7I0hoec4gJNVvK2Eb9t6MPJEUj2zvjlM6ZEp1QekQX0hM
C+tYSWxhT8eYN8VWDpvU9hZD5FLC5RNnwwypUt/yd5juhy476DXa+5uNETADAmkQiFsSmn0M6WHF
eq5/esBXJjwVUqE3DIkI42CTH3EGNa+Uj4XoDS+RcEag+dV/DUie/ANhM9k22wWY5q4cN4v9dvFI
qR+gChN8rELiFiE/g+IXAIKVqXVjUmBUus/MjauE0ccQ27Q6P3RGpH8uGxYvAEOzyzX3llSlSe9C
Wv0QfvYBLKwy/LeCChG/Dn795s8lblzrAJKkE8FSVxKZD/x6gePbKQJf2BIigPt4ZnoDhjB0x9nB
zQJGOdn3OnIfzHrP6ip7xDFmTQ3GiF2JjR7oEZOkTrGYDiWavTGL+LXWtv7Gl3hCfAixebpLzC/c
tuzE/qUs0+WFuGUldT/3eDEBDtHQKAK3IvdlkFUosbbdijLQf5uz+IvdwpYNKAmRySxC6ES5HUMp
YHdGbKtWb6T4MU2rpGlfXOHecRdNzTV5LQvJs5PWlGXtnT1M/nOyxeRS9fuGuIZjAjCH6I2SXyfU
BxeaK9zCDHeZF/j3k1PIQwyKdWN8jZ9swO4reBkqBVyuN2/Sh47Y3+mdY0W/RjEmUSBKVOsveRhe
Y3BhnhrDar42Z0HmSTz9jsbi97RqJ77vdLEo5bbILTPlUVHDIa79FBjhGmfg3LMakDNh9YGbKPC/
MSMGxlIiGBXOgF1tQ+6SgO4JLc9rLddPkiS91Rny/hNr/Ozj1c1Q5VX1Athi8NA3s6kyjTlIVVtr
b3Ax8Oq3GWfLPU5fWU7kwYnyn64v8niFq5d7GKp5iPCM5jmt26N0xTMBA/aVtbMGoamW8TAniwDE
YLpE8vnxaQh3IxBkDVdUEc4itlbTCjFxQPlzUSEEcjZB23Edx2VdUHVcHTMMLVacO+Bv8EYgCX0S
8sXYQWxqaQzdA7os43u/MhfIH80DLSKgkLNKaAKS5uwqK3T6FfA2sgb+8H45N+4QPgoeUhwezgh2
XyxxmBswgT3ZrivHIE4pbY3mwFZWIjp/20T/Z2FTlb84qUm8CLmUzcHJrKieWr52p/vLqUJPOhMh
vCooAUIwJ6aGPsQ1aqoyKw9k6EpSAkEKqlXQlO26RzXDYjOABLO0IEo+z6vepo1JGLWImy0KtgC8
9MERo0f0iDtVfmt7NpGZp/hm9UKIDyvdLLBdsn5rLh3KuqQzvcxDDEbB5WnWg/0zub2L6OpRbzaH
uDr1wkLSnUFzTlhTCEQoUaFYEOLM+PxU/8F9XCdbIosG0TgsTd7mchqZUIs1/9/emwSG7ThFnfF3
jk266kYQ4Zd5tlbMcCA2VczkFHy5anZd5MCxSh+RG9qpUCX7qZ6GLTRGFnKdJo5az10lLDhJhXU9
VFEARhK3d3pZC3O/XmXumiEHDQjKB1OVK6XIsJ2ZQVfKumvYQq4R1rxGXI28sH5+ZLvnAdcroxya
Q4HeK5ePTphT0OZrQLBAA18q7O+2/6PbnZHZ83EXkQarRfREwCoQ4q3MPlV6fY5vOfmEdGUJgVA/
j3cxm5J20+LuGJZTlYk8XcORC94/CksbsGI4FZOkZC19BW+MwQD4gyWqUt7siWhdx8l6/Sjxd6xm
3XJatfMQw4Dy7GTB6F1dFUdzm3c5ARueomPn2Cr30HSkdGRgXejAjOkichRBpPdfLbPzppyOMaLR
MFQnvqDqPGs41o2B8V5eEcTy7t4v4/uJfbjl8f7eSNlAhQhIJRBdQgRCHjYIGMmBja7zDvxNtPHQ
zwBeyoSneBifJdCqpddvi7vCNu9RyDS3ljtSQX5aujldDyYut3U3iv08ezHfy+hRLLT2BR9wFEaC
IGqri2pG1nVnQFnp7kGQXUPdi3HZ7uUswbGPWijtcp2zx8eMx4a1aiRQ1RwUj/+B+ook0CKE5RoQ
NN3SCMSgtvKnBs8iFW6hJj+GC6YCStotNnVAwwx3888q1Foq2dkhqPePzatgfy2t89kBSFKAhSvg
d+7M7zeVPYrHZagbQ1AdM9EexArGRUUwwf9LBVE1/hnjMRWAk26+76MgLujQhPGnbYLvQhVWXAjY
UD90Ebywhnf6NpDkcR1XzKgES2Uwc1j5/B4QYLhwLpllVzV1Bsmc4LYV2LROa0aBU/OEneCsCYcm
X1tvinbOwjS7Ba9KlH3amOdntLa9ImnFbUt5gDz9uhp47ZPC+z7Ht36Rh6+1P14ugmuSHYXHTCwv
zhHdIVLlyMvUtSDhjqGy2nGyhiR/63U0CJDyx5wTKM1gr2OgCEvXWNk35q9bwrETamZTwQdlSEPo
3mLhm32GuVbVLy43cr//PJwvSNuVZStgYtYIKEjwTrlBePKh45+l8AMc7jt4/exxZ01poimqpeK0
FlAQUI2T4TBuIKG1XimOxzihIOdC8CN2c3LySTuWIWnXnJAd6Bu4Qoa/sclLWVNHsjr4MtOESLE1
mBXg8AhYiqPUxfmG1guY9ffznepm9MKGigDO68RaJt8F64fNW5mvU4HmRsSE6QUuzSGhn/W+h03k
JrBx31SOil8YxFyF+CMHaCcK0f1iWl/lFYOigoIMxuz1D012w/710iK/6+izuGzjeeZFWNd16pBy
KlHRj8pZwbLHcOetLUVEqgjWzXIJCUrWnyCk089Uus9lb6R4ChMJBiTSnJHI/EuWiNkjyrT6EVO5
NcQhwECU9csnBepsKppPQCZfcJ+a5SLTg5vNp4s2h6SNxbhvuRSWtmC3gyWD/G/ujaYzZG5kh50Q
IVTOQtK030+D7zS/5c2XxIPoYMvgLBb8TDHJDWo/4zeUyQhBGwh8ZNu4/zbOJB/26jVV1JpaNj2u
gvfUJsZGpfOzrYU0Oe/qbgUb/XaxPAYP08eKhSEM06mQJR0waGO0OzOssdDzd6ROaZP2syzaZaV5
RVScfFLUz214o9+VEuPQHXcbkIp7KP0Wm8aPJBHPYiT2M0pW3QtbQaHr6uaOTifbnodKFJJUtdKQ
4PGbsgNno8cph36pyXxezRlrULvljerFxsT9LBNQj7hsauIIHpuYPNXEKQ3Jky6gSdri+aeqqK3b
Oicm07+Y+sa2gM9SY4sdoqgQdJSuY2us3AdGz5bbLjzbLJMG995bSIkoIBgGa5uAKFRi8m7JnrzS
20I6+K9AlplO491Ji0N8l9QkS6TfQfg7q/ZqlpIVQLKwzQ/EE5zQMt5uFEYcwyqaDuWqt+lSmKVz
8r7Wn9rE/d88HrqD+dseu2/GYDYA2vOu5KoVHpj5upED5KLbiBK5ibaSGAVw1YA8Xr8slzC1gfyg
ga81ANRFCPXyj/q2n8suLLcIop3uPh5makXSoU2X9KjLGfd3WGQ0Lna6BiXkLgtwpKOdVRyFMSuU
TE9hCoARyrCp5x6ah2f1h6ycyKHDD+u6r0BtblyfwTWRc4CnwjgEqVNxXzg7CPueLIEZnFr1J2/P
vekg85qAEY7sNkwWQ3bMk+rfrYVlZUAX9wdNVUzly4+dE+3Fko12+SAw8mgriGKrvmz1A/S/k80q
8BCkHLPQdOBUd8VfvjAfxYFwgMYFaiEKAOe8zhQ010yEdsSw74tnEj2TV3YPL2RQFfgj6rijyCvP
/ZeXe9+KUF2LtjzLGSbRtyCqN6Xw5d8M3M6JbE9axPT5EQEt2iNMW9zsunPp+EN8ubjqe9qFMyop
dy/sbyu2ekDaNkftIZR/1K6zp1V2yhgj9JBd6QuhK3pG6bE5iFBuxJVSiUehrUHr6Kk/wmZ9Li4M
TIzv5qaG5oWZra60b9y4I6QHDVOArOoXPGzay7wtbLU6eUUMKPina8V1bBcDmVtjZI0DkV8//WhU
KfoDclMDCHgOHctgsifrSLAfNnACDFaXLozpKcZv14M9QvA8QBOCpmUEK4mhTULkydRwst3lu3Ah
+/6mPy5Mvr0U0ShVYmdonAaoVtsNst4TN9IXa3FQb5oFlGjD0fPnWFPUAe0zDMBngcJxSrg77ATL
GDHfBPYucrGnP5btlT5vfdrVe+F8Hyry4/v1sJEXuRISOl0U9jt0be/SA1EMpokLl+2TW7P7ec3x
pzNwaSKge88I6hZdEBEgCYsOHR58XOkg9Q1tmRu0ICxMD1dWg2EYZRwM+L3JyrUE8YCGy6+anw2f
MR30v5CnSxmJA+9YOeTp3G6niXaoNDfRi3VT5rPeLmX/4KwFluD0+69n2Oj9wP4RWyG7TovQp/FT
pR9YLSDXibYOvAPRHpqjiwJ1rpHMkA9wT8vXe/GEOEMzGi/N4dFCtMMLtUPyNnOPL41idSz4ng+9
KZt3GRmunVlKw6orJs6ne+HBgD1XxEcsk9W+GT8tewHquMO1/WtZXNaxlbF9MmRTHOdEO3wlVbLO
7GskFcWrts+JW7+rEGr6acqm33Vx4b72yx50nMswYrWSzgK45BJfHhvyRKBV43P72OTQoQCCsch3
vEorqrLMc+0i1foDlKmbjHB+NacCiKkYAiM0XXpoGGcWF2tIHNCb+1I2kh6nnzULn5jU2Yhe8/qT
Ts0o1u26j4QR5FiFBO+6qKQhSjyRA89Exr+31LBGaEdq1neDaXNqPkz19qzOmobWVfg59sgHxMpB
0xQBEO26gIYKeKHYUUmM0w9XgZXJYUfKRGoVzmq99+NKBWG3spG3yY9QDs1BacRnJdKgpmDK/9aG
KEwSaGNmnRsRvj90HajaL/Ae/PlJ8ez5I07fnlKZtAcddpa7sCiSxEHBSa8lMbKlWr6tz8k0JevI
8sfQr0RiliWPVNKi6mZIuLzkcPmiaYIZNyl27aQSSW3BGxkHVgFkwvsGzL33FKP0cRRG1zb70fve
c+xhmIQ949WsceXQ0WB8vtcJ6kJute5jnz9qTXeF08G52gjd44yLrX2BNnZrgk+7SFFCM629Le2S
TkTKPpA4PCYNDuyVK0TguofddNyDdJGdnBVTra1n0VnFdYRSAyUXVe5gEgPHwV9qrJbEWz8L/dTD
0cybd4hZv2roUacxD/4hc0x6LA2wjBB2SxVENpy9xS53j5Lwxp+D7H82JPH9QwsoY9uBQ81zEiex
ACAKouPA160gBJbBCaWcXpXYdadY+tSe/kGFbfwl2z5MqRuGJSetQRmgQa4riGEx71y+kuIasqDf
b9fZDtCTNrCaMhSpe0G9LOSmQZjY+5weWBQZG1hYtSGxcHzUUaQ0MrAIjK6qK/2u0vHVD/alvE1v
s6y3c3GO5N7hQ0Gg5V7/YkLZq/epHpV8BeLcs8IuL6b97aQfwzwfJss2qkhm9j40c/FWM3WRXGOQ
X/hZzmIiVlN9vJwo50sL8CG1i76xi+iV6AFTrLe0We50eNDyNu9D61IETwuEYxllpj7s24ikxdtg
6w3Fv90VuvqWfcS/Do46Zp36BPLsnByz4FVIE5TUjbac7Hti3nDFjmOGqJyNIrpGy0AuAXH1OQ++
8W23tjEzuDBJohsZ26ZGvfNA6dyBb0fBO0JnGTnd8xNGdC7EY1EUu76kA28ZE/PRRKT9kUPaFhhi
BhLZrbKteTFJAv1SD0XnuEyox/fb8CnOsjoct2E5MqTpwvHdI/7ga9xVgRHJTJADRMS+U4K8bG1f
G00Le5UzSatWEhAOs3OK+a0amtQ0xDLkyAhI38RLDdU4HKvqUWwfRNlkzU0cU/GeGTYzG3Xnohgr
EssCi+4gCd7Ys5Xkeh6BOMrzbfyoFXWsDJrs0af3HiG0p3bTJZbpGL0jgswqYIO4Ah7D2Tg968yo
TYTzCX8u6+H0KImQVZ1FlRJ9+zXZqfcR4hudk6b6i20KNjJEyPcJtS/5a6eRN9oLNJimsd9UF0oY
xnxqjHWnfjJdIDHTj4MOVvhe7oP91Tf1Nn/NFyrrGkMEpjIE1fwo0ttDKtLkttdSrwbYE3eDx6eX
YiYx4Hoxp9dw+pg8SFkKG8y90XO+0qvNgODOZtOArmjEEdN8lQe0Pfk4hthwfm7moV91iDBFJU+q
6oRU+F6YjRtbTjZ4RFwi+nokveaduH+IRJlQdtNGZUIfPMta6c/QkCDruUODrWT9H29QFnraLWDD
fdO4Cd0uoNzVki60yhV2JsA9Ktb48UZNRZ0MCVkTqhZd6yidrf24WDE9qAGHSNeS51pfxCCzt6Pt
bI00w4kNNap+5aR8+plkBSeWsza3S/Q9jUc337hlUy8YOVw0Ex3zBy7zLh1v4YFuXnOVq8x9JjfK
ko6vwIjHYFqN+wb6CnrWACReWTjEQHeAP/dpsQhUfpRqp34w7SqeZxSPHSrBpEDMpLqPmTXHfHQ/
q9QQsDYpuKb3/yO22FzjdMZO7pIwIrgDbboWm3a4hF7YyxCrgss/1uHlgcVgN4CqRK9JLIFOBN43
/znEvbAqWVCosKNUHG2c+oYpCiw3Pc1WFqXR/AEz/SdKL6BWCJeqzxho5cb/bdlIvAbgfnKv6eIm
i+OFgVPTiqNnlvrebgcHNjTnIsffFgMExNFhYLsOS6irznV2AS5e+wtvPoDcYn17ShJ4EC+WaIjh
FMnDYDmZS0kdTMWbJuBA7AoGx49+2QNh2fmZhDsAbLKnw09lNLNsdr0IJoWiwFBdm5Na/FDYqE/Q
I2epUF1p0tZFZ6GKZdi4Pt5Il3jtOwEvISCicgNBjcZEZ1HiAtZ4TUxXifj2OY63XILpkoHF45b0
Dy9FOzbK/e4bsqDGxGqjSSBz60o5FZpf4r6Gdz7CnPcixAH1qpKdh8cKoy1XAGnvXN4o2CXUOBuK
SeYxpx1NSrkJ96pmM1T2bz4i3fErzRHTT1Ghl9Ye42vuD1e9i97IJmWI9Ybkv3h0A7pMUUZVqUv2
Gf/rufHRtD8nFordYc8R1vBBW7k3x7mPnIHlLHEf2pcBx2YpSQb6ATPNl1WE5hShuUKl4pL0zObj
PGi45CstVLeHBX+7hSJMQn1ylKUifTT8kIncHuPPmzIbICkUX/D3SPpXzlpb/15sGra6dJAWiUO7
wMN+87UqBIGpMOywZzeSFU3pefNJJxLxnTl+Ga11sIiEi4Qc26r/BNODyxqGkmpfio+kdhv0Czv+
T6mzljDJHv/X7nEiEQ3qxD3FX496q13EQoeEUEzbTkX3aJ7+iXysoUsNxWHLSHRTp+D9yKYD+Afp
lYiDz8YqY+vyNSHYEhzdl6Ag9Un3FTquWB8dDm8Ua4WkJoQa/BY1iM8ohoGGx3FfpPAJjB4Ddzrk
ionKQUXteW0KEP8vUqM0CXm31lFeidpFNgNVUkuoqm4DT63eC+6WzSDfJqQ4BATlNAy7V/XNS2G5
Uk0xYcHREK+kNrWEuK5AXwm0F/7vguGh0/R2cBHXlXSPtuhX+svJy7lD1IZybmlUTFWHFb3Dk7R6
MfmuOoWuNdXmzoejf2VQv7mQQFFVjzS83/7xiSOVIE0L0UA90x+PxDA686ENehxuO9hsXBEPIr2w
53zdHhTlpQ8F/CmdwQX+Ern5Z/TnHSJ5Rlp9gPQ4viSy8uvsdmvWkGJFpyzWdmogAMkwSdJdlsqx
DOnHZ7RSEVnCIgddpF3XgBOHu0pHvBEGu+k0lAkkKe0+YOT2ChippetB6HVmGTopy5+4BCpAbQlj
nShBmAiZD81gA+VKRKXMTS1o6KLA5Nca7KLku0d7yKX+PQSrt+3ZRW/lv+7yL1bNPMEqBLBhEwnp
RjH3aG3rn6zn5Aq7PvKicapPWQBU/fbz2JiTp1YS1kGIRkuIxcBK7RIhNqu3ANDHbvoKCv6/Aqo2
/WcOwLk3ikSkUc4LOCz6a5DOx0Nvj9seHPqLYjTbxDY9HsM+YPNGTWFB7VYhBsa7NEZobvurkxXh
fwl+W/ShfrpWgbuLT7d7yQCgb5HqmQY7YTrp6hADPP1OXP196IcpbJKvxmMyOrQBbK2/sS7di1V1
ArhVGErBgh8xm6THJwUpYOht+uMh/MRzSQub344hAAdXNkU/ShhqsUc2UPmQdwmRHB9zWtTBbTC2
Ze1addJdk6NspkxTnwwEmP3/v1mIRqT6o5qbsGSHChhiaXYVOdSXLoaStH9lFaHYFtjlAyjGqe1R
9Fl8Uvf99DOyEmSYpx1HqK/l5WCIPQvFozjN6hjtidIYz4q0xO9twscbz5nw5bo4roPEcyrhzeGK
lZVYcVpn2/q0+vvRMELyJkwNhVmezrmFFThyKfQl4vN0O0k0lbiXVJ3qbLFI6PY0r8GHeSN0futP
MdwLgwnBrSq2xT2sdfsE8KZXx2CrdS0T4wewoAvMiekzJLXFOKsiXR7OzkcFPk6SASn+xGK25thU
JmIg6pH9e2peeUcX0lJQ+kHhQhtyQjLnu0+DwkHyolihccREYk8dKbKBTCk9EvL+S9V/A6lGD5oe
0wrnhbdjU7FmQw72BdYK1XlLc7/KigUdfAOE7wRoUWf//1z8zVASnWKgSKAUmpZP2DR0Qcc4Jj+F
x5jNmns3bGAPr/sSiWpAVW2ughPusGHmU/nx/0bXwpMPICxOrQV1yg8Ss2TggOC/B1p4wuZmDoDh
wgD2TTE9bswnvAfrLby1pBk+sfLYejnL5b56QjLYFkKF8FqJa+WVRbjuoZemIbra5tfXuU7fDPc/
wv4P4StKMTXjG/nb28WvKQ9wd+AATwQK+m49z04sDP8ld3pDBiQQiLkszwJ86mho888iBfTTHK9w
dAafI21/ea3KK6DDLEwxptEofiC44BSFgBylzN7s8wfPNKuIEcoq4FnVWjS0e3gilhgG3uSfofdO
byeK7GvjYXT811dyL0H87A2K7lkilGTpqoF2+RKOAFelHZAlqM3d1eGctMeRUqJGL2Wv76lIoVnL
BKqryhBQZXb3ZZSTRIgVT9+FHsX9EqVSbsOfgkeJ4WonQaZ3/+CQPzUj2BIkYUxaM6BN2HSZKNKQ
r5AOCFN5yaIj1/qB95CU0GQ/OcH7wK8p98hHUycuvH02aXC3tK2UyMyrbO5b4b02otVbOlwJ+vKK
qFaYUlOlSduM8ddLqUgvHPFruW/4WpRjrZmIe/7IoKsnhS97/u++vjqU/zwJ3XfebgJTSm65LU9l
6pYrV+x4VLbkzGkHadSz1wpCugLPG0i8L/DkzX35JrM6miOJ7oDXW+Bv0lo37CwMbfaX+CWRMO7O
2bTyL7tjuCuZiSDgd/JJKlYIjcBRqIFdoJo2NcAmPxQ8Itloq5D5NuicqmGLnve6mb2ZA3pdvLML
4amx04fYhB8sfVAfBU8Q4aKAk+7eQc2E9vQuFs5EA+7dVyw1z6ETgkars8KHrz7QeJvFpA5OKmdX
Le530i1JnzBRj/DWEvfYaWrDdj7YP5sIvVMmPKksKtISAbNzk2i9i1oDt1G5zc03oO7CWsqOccGT
h++6FCzq2nafqbbfPa+DlmVA+8us2hM2L+pBnitf4yUUgIsiek9tmL3lR5XeaTiWSpt52wAuJtZo
qf1rInRLxa0zI1bcA4cvVAwbHcg6XGuCueY/cFX4lEFIJmLrBbHGbqm7THv6VzwTfPuMZ8z6w8+I
gaw04TOTx5hmUdpfEPUKkS4maB5vz8tsTePYXROSbVN5BinNNKp6y5Ntlcmcqqg6mpPGEgYSimEQ
esEIloampnsCexQAxrALqI7oFX7Qty72r+1umM6BDkUltSp6KuTlu6fGDrhUp9zvgxfET1qqfVQI
csz14TFwsKsS565odpMnz0+eU0X8sfXHbOOBwhcZGEyuETOosAWpKRNAzuYQqV6wKEXhVHM+77k9
JgF2TmTbd6IrQ1L10WCQL3UG7bbnTIZIDXD5B92MXbYz4GINtdGozkcANAQVBM5pPpkZC/TEpdoz
Gx/aVR5jgG1ki7vbeJst+Lcsf8JyvzE9r+RNFdQ1YO2Qe1pnbBuvNqmhNeo0KpTwWxWapxuB047Q
Q9ok/yrkeUAz8sDEzQ5aqh+UqiWsyuczZwnKXllyKnJqAcH6n7jXQYmaSbjvqfZP33Tvji3EPQ9p
irMRwjK+zdp3NP2+4dwZCXYnOMAuDx+GpnsanMkcJ7TyCFzk8M/s4QEYUWl/rOj0qg9Itzm/nw26
8sQzaleXinkErro7YAj+FOCvo38/n/kuAFqgQSDn8c2D7dB3FqVDvCbH/rUQ8sF+ly335fFNxlfq
lZzBma0cfWqNNlaRZQI+tlGfQr5abYPjco7FhYRp6O93Yk7XK8roUGm11jPi3pnQOK1quBcTBa+u
7iTRj1VjivyMtTJ4wBO8PVwWZY8N6+Vs+90f5P8IQMHDZcrC34uMPHpnRhJakFydiq0YFqt2pLGz
TzBpRDAfYrU8I9GYflto8mjI2e7FZ8yp3+WnqM8fzLATyJrJ3XzCLZgSOiWSicD6otBsdVkwD5Ka
l/MLKctyvVJuGMCUeqyuisewn+kAfjqgZAzsEgFyz0xvyaQO6dJo1VVYyc6g4ahnG10I7o+m5giy
hOzrGdMXZxD0JsBJ2Bwpp5wJaP9YoeMW4TLtyaHprIxSeajk+L0uu/lJWED4ZhOQATRZwMQij4UF
Tc6Ujge4gEI3+K/8KEIU0YBf/eSaFeEvQ3TRhBVor0sQqJYnA1ItmGd9VkxCO7FPBxE7maEzRNEt
7fWeAzxN75TbIgYJAIDhVOhrKIZZgdHAOY4P60h5lxBPQT17/4i5eEqjDEvPU0yCrJ7ABPDpl+LJ
WHeD1RrDMRfqXsX4E82q4k3PCIe+zHnTshJSg53kZlh5bD/qPyaLVV/gMMXYtcVGgh+wryRK9alL
iyNv9/gz3NtS/HPXQ44OiGaI+xblePjxkxJU2hfYZ24qLdl/oIU+Re0BLZgErLwkmEh67bsEVBhs
TytA+WPOXYKj7T7KMhD1U4M7Snjz5cQw+0yLIeCi5rVPkSfMXgdGY1QthRTpo6CtV1AHEY+cJWZx
JkTQGu8leL+pSnShmocCki8VAVZbKtNPRZCF/IlVfkUdp/6gRJkeLEQxKvW9StUDYvIl60QCKkXH
gZNmQgTdL2HciY3bjchMebhd6TNLjjKQHER7VJnG5/bLR9KcJyjufPQ1QFmRTOgxbzpOPUaxlT/M
OiIU6TYFD+8GY3pxJ/xutdxpBT/WWdGdReYWvzr+QCsdzoUs/Ck8dUij+WSDZ+ZE8QnMlhu463wZ
TIZgkZHdWLIeeRA4IiAbdg50TjAgUt+I+Sz7tvKhENJ1pA0N7jkQ1qN40iAvV/YpxSuUQw0S0NTW
Lmpl92HsBIGA/KtNZlcabna/iu4quSuyhMvyAKulZZGplQAXXGKSK20M2dVHwiFq27NMwdM7ZOJ5
5LaizcFgljXW0d6217hUc1KrWt4c48q92K0FYkLXBxbK4OstfBSjiWCeC0HsyIqmv2cRPKH1cg3c
zc3n6nFAIWFlkE4qQyTN9IzVosbAaErIwiU8ceRleTOxEYqS/nMEN4AQv24pT2MUAg+LP2Zbniyb
5L3wt1jHFJ9cptoID5Dnn1KOMBONmEzcGCKzy2OP7G0Y3cdsu0rkcJtTRwwJnkbDeHUS1zuHEWxd
6qnndlCXmR5zChPi4DB6KuSTG2mmouSnniG7lr3RO4nXsS7HhUycNgzf6dCfd+dOs3qSJzVLhUNk
AXput6O6fkMpUQUn8YCiEEhm+m6wkipoBSkOvTbEiFblov5BjttpKyzfuNl3C6PvSXWY/Cbt1fBw
t2O27sKsQiCWMTmoHRvEKsI8LSmYsk1O9ykuzCRhyjj4XT2DxthzVB18Qd8LkEHqmEPG5ydY374t
NvjFLUQTNCn8F14DLLVR+ZosQpAh+65jTPf83/KZ0TtdRpiBmlkv4Yq4x8PAHiEPlr3l9yxU8A3w
gERg18q8KB5EUexuHyY3BLRBCNN8bK3Tbi9uUnuR3c/TE5wzB0U9lVoGqx+rX1/8kAD432G1rAap
IKrImGfQptSnH0f0CybxPyYFpw8THXSotYc0iyEEVzo50bWqsCcu31jiCJYol1YhGLKtOaQQDcYZ
6trY9AL8ZA3Q99oIA9xQz/ShbHc/J3NgLvBMo1mkUiSqmdQ+OosDVnIK56hfOL0WlzkkWrs86JkT
DAE2vSPCLbnyTT0WyLY4rxhwmxRLXn0k0gJWz+3lB/j/9B5MHpBFa1Cy4ApNufoCg5ywAwf6wl2/
kwhYkNHFtvlBfCSzInn4O5Gi7F9Uyj6+l/j0xy17zse4M1woFwnmnzaWPIgctTzH3MV3k50whzzt
WyiINLVQPCLWfeoFCsJlDM/zBas0oqkUHoHM+MyQ68JWzwUFCTZdfJfLQR1kS0045bzXt0tx7bo7
C779YqbpoYgIzs7Amn8h6a2HEhB8i+m2GYPlksVo79AKc7rjDbq0gzHoU2fe6d1OpHjjEMzVO6/j
OMtlOU4fuDyKuOGyNGoXwJckIoFmQkJrmrURyABGwakY+YS+okKEZ2PU5hMzYwLj0OqG0mQr+4Yl
mYSJqI2omLZqJn+s9CAIdjmDV/nD2Lp3xsQeWkyiSpVWKcJU98+nt8vppoJHCBep3+KF2rdN4HgZ
9NO1BJazipNH+CmiRHsngLHFyHYU6ER+JIDJ59XqSu+mrInS1u9jB5d0L0phkkRERFHpMtRcQHPV
Ju0BKy7E7fgIgcNL5j13GogaqqF8i83tOGur/hFCU/sz5X2IP7yclt3TwaaGvnWUM4J5Fqhvqpan
RCJ6l+/AIsGlojIAVGWM3ct3W0ZOgqT49JA4IZ8r6ODL7szxeuTJDVeUe0fNysXfp8hmeCD8sW5Y
KdlIXzrwz88s1VZFm19BRjNHo3xaOAVPoqxZJAi+kkp7PmBSjZsqb/fR+lPCUxplnBHAVm6ly3KQ
4ji4MfMqa6pRT/sxFp2+2OYbrDoTDa1zw9aiiEcuzWPeIt1yUZhVxrKav2K+RZzRMARt46lGWnnx
9c+I9cGwXfzJKt8hZF+hKwnshM0/AGmfH/gP3/erMOjCvNcBEqxNY6SBsmKpKZj1b4RmvDQ6Ki6d
vpo6hmQivWe6qAEoLcGjICmVdndp0xE/4Q6hd+4JodrgtJ7r3z8+0bdTrfyu9YIGksDI9khqWQhQ
Mk+PPudJHR1p+u3LG4RIzm8iVg1zKpyKYt7Fln7vsNpycuIt91mNA8hZDMgn9wE9baY6r+Q2geMt
ltiT4Zcy3ksP+BSe9NVX3oL/uMfCIaBAYajlxi5tpPG8zB6pOeu3YCaAz5dTQmm0nmt2FtvzEHxa
4wjEgtYm0tIJbu5FArF5BW5V6z3hIJsqeDi9v2CxYPeZpgoeOqG1YNU9avJtGyOV6T98tVpqUPti
l87A53iWuQ/nC4tT7UnH1vpTigpCuC/QlPxPIF36o2FTHcw8/5PM++RNeGwOq5VItf/euQs6Ku4T
SOy4h6GBTt/DjEU/Ld80RNyQ8n/gRBrWWhvHoG2VIKq4cP8BbyWaGzEaWckwZWd20d6D6O8OX1lF
GLdC3SBcAG7j8gFM+BB2Y14CqQYKVpAob9+0MlNFFpOEZY+GHPd08IrIRKxpGFnPN9UfMepsza+c
YKNDL5/j6VaxX8Brr+xbuSC/UMrOut48t1/5Je4gVE9Lc4r02YnbJnuPLYDviGhO6Pg5YzMt8n5t
hmKW3co09ZhvrD6h4W+okqqJT+4RS82mzL5eInUsJTuQCaK7aRrDrfw3yTOuLJ5R2oIL3O1sM1HS
JqFxOFfiMBdm7JSUWiRdDk11rH11GJ/Ap+yEb7J8mnFbpmLBRZ+TzhYEr2g6EBvG+ZgUAYQ2kjhw
wgOCa6cB22gjX550p8P67aqkRi96n3dRi+MpQg0CP26GTKtPnD+B9yfMmos29bAKDRR87FwRUn/v
OCaf3eQ6/okk7jJrxsKVOORlPCMFFON68P5bfgJGOvlz1YBG7f/GRckb7pCneX27fK3Y5wB6VV0M
Jk2uf3bljCe5pRcjjPd376CVQFU8ue1RLMeYA216ii7QCRp34ST9kF4U8bX5jOOqvV5GhufHegnb
2Zjhkvew+FfAy6XF2HgGNBuzF3pgvfAXcSexA+9TKKxWoOAk3FVgCMMHDlulf6qgY3YJcnFwzDlA
UBJ5UVisXeaWyW9nKkNSN5Zuxn3JQ5oQTWXDsQ0/m+IFIx6n6xGvl8zPEuPBlCcJxQUuWrOhz1XL
AZEfK2sfi9mQSTJ+EFgxyRBfrenuRxj92U5dKzZ0S9MDaG3HQI+HTg61pdHwS9ziPtJ8Jtwk7g8y
HfQVlHhh0xmdQINSXqBZNXn1Le1TRi27A1ig347o/J58hpknTUDTh9DAyZjk8VQziCHuswpNnDhL
l1zbCXzECsWPZXWVgDeNXA3KXRq7k7hruHEwka/gXaX14bsJe8VZ9aaIGFHfyGXPuKYbZ7ivnTVO
xDc2/MWwKHxBzo2NO495u3iI06rchdBJ2uenv9fSBTj9it0BQiwZ46wVnj87vv0AsbkNs6HswZ1e
NpRfitZcHdGTzj+W4hxj7Yw3OPRj8RcrSDAI4jQzdomxc3/QeFIGwf9FEDCA5KL4Ow/ImMObhMPi
uEW2YQhM8VpvcJAi4FkF77RIXnAl5cfvNL2jVNIU0cH2xtBO9peQkBx8mgpKpk0HqOm3o2DtutF4
p7ueBMNajpYUcRDigP5JikJx6RWRISoiPW5gmsDu5OquqkK6SpJu2wYB5aCdA5BvnQIkDdlrE9Fe
DvSnR1LYB/dIYsIyF2alSfDyUEbJGYs2k1dVZ3uLtFqWoP+FR7fWMeezmLIsfdn5sKGLFLLUwMFq
f422L8cZYY1wXsplhYd9+KhgSYp2vNZ56hYJYwwyo0fGUCcX3+Ygu3pt7XLTxqGS+d2Wc24N+3XX
dWiUGO8215Nnfnm330khLqSIXlVgDwGF5M4cQB39UwJg8ysZIExIqW5xwL1gbZQQf1W0MEqpux5X
SUJ8ZoBJaEAhDFXz8PTA9O2YLqgZpSgk09HHakxYu9V/diyWe0SNTXfhSy9+HrD7pEEAfpI3L5+W
jNZBVe/lqBhqVo6ijtB9nWTwZEXoEy3AStTe2NqhpIQUsa+dypbl5Sv9gljDyniTi9rURpgZN7lH
ThuZnpW+X1zSZgtNCzBxQJYaAtszfnGDfXQuQ99kA5E4ClLJP8IIRWetlOxbDHlwzkrfbwjPHcd+
th4w+FTKMLWTEbdz3zLiivrGHCEpiaIF7Tv2yZlQzZiwwT5BXslJ6w1PaP5fbkDk/5qtkM9CK3Ed
kK0WcaMq9k4uh93ckpvtc6av7A6SaXQLNG03bxGs/ohtqghf2nuFcdCovP/yFtaSWBMz/r2wr1AV
Eh+T4DOI4Tg9EkrK7EQhF67eOYEo1g6Sgz6Gaekixx74uSBJJd9SkDk4QXdkyHKCLEjE+KR/rMYZ
In3ZRuGsX9x3i61GrQCa7PesiAUkOvWMXzRE8zAy7hV1682TLnoS6WXPFBd37mKj78p4z3LxxgRk
7SQ6BeHtJQqm3lUgFgXLR0d/s3xfe0CTVaHCKRd1GuM934DAgwpM8uuKe1YYSmQmzLDQqkWrmlWy
KvWGQrKZPYFlswSBmHCnAuJWDs42S2uRT8fAAjGDHru7WmQNaoVR9usVihb6aqOExZUCVFcS0uRj
y7GaONX+8lt5PJ+EKOD7rBNWH0Seov6BfqiJ94xqbWa2nZXLCIb0gXi74DFhQFDsZGHaGHeBOX9Q
sLvP5/hhScJtCwgJIWQ39WkEq+qD7sdWGdDQuruOXYxGdWFYV1b8wlx6JYUhHKr+qg7lgVRzLYfX
v6wnXQMRKGFQnXr6+BdCIgGMQbeUv/twrI6CmLO8QfrnXqYjZhbrKou4cky6T/DZR1Lh4JAgTVZC
+1mXOyiE1cUPFlw4P6EEjkPGdSw//4ToBqKEeXZTRhDF15KNbl2XvIS9VWOnHr++qfHnUIebMV30
ya2NCGrIVl/mmC9gGGFZFqj39JO19AqrTerhHxB8unIe1n4XsTcWAvZQ3jNoi9oOgABo9W9s3KLi
YYRN5wa2oWmm6oe2Athyo5bhESCINmSNg4rjNkXfH6h9H8pXtjOuuSLWlnMa97cCIxfBygVaJzux
g9gwRFyXZmwVx7KyUC84SHp1VuIM8qSQU3mFWZu5Qgtd+0SpgPx8cGLnD6ZDbAAmUL65se6WN1vF
OPqkTilrdMg66cgaqQpFYlJDSuydhvdOYTp8p0PIW4YwAsjhA8LKHI2/wKPHhiVsOxPfcS5fmun4
IS4QOjqRXQlFc/zJPwzvaP0MQ6nXUJbPieqROucMV9wFRfrcVzc6Mw1YUi3drygsvaJnJjqoh0Wg
48bzF+jjazY2nwWDJIJdOyeXLWSFQfkFh2ADmbGEZH2aoSgFo/orxaqg8Qln73OeqlTBUnv66vYo
VCAa1p2CNSEDXmT0yqhJp0EKNhsV75k8TDed+oiJdi7m7KRp+MrLBQYGbRa3bKg9jYFOs395K/Pz
3k9xIWx9EXPp8CD61kOunDoArI2/8wPpfBTeOJfGaM6jZe5Tgi5LJkf1MoldFnFHqELVjSlH1+4b
7FAth8JAwm3O+wdvhxXw5CPKpnccmilxNRefLczQ+/PUFygv0MKqnJFxyed1JFT3ha1f8vuMCSsS
EDjVfrTH2n1RAS81pS7CSWDrjkzT+ayDS/44X1JgSeu+Bh4MkUflR4vpLwCjAhuE96PWWvsHytgo
1UaJ/LA9GQR1Gzsx4oRQ+84QOBUjrMDSx8zwSw2wlwEjUW0LmIfLLGqvnvefsIYfzQCbpxxl39VO
Hm5MxKSqFLYNOBpy0hyP2L351t2Dp8Rc1UB/IEn6DWXHFn3kxCNmpxAJXD1h38bsvitKmhsVLegQ
Ur+2LdYhPBbanezeNieKMDoIAqRDDTrnLXne84ZC1pvRH7h/OHKqAZYQ23XKEC1DIf3lG/6Zhueg
n/1qJmNIqaAsaLP/hwt8qWRxbQuPvh6qtwTPtOHl5BbwNnCZyouF3W77CuIfeCpZWZVq1reJGBA3
gqroaTana2dlsH6arYxwRb+Lhi8qrNV9Ggatdcnne6WugadYDxXJQzfmasFNBIz1ZRK5eO8oiPRK
XeRIri0OOwec2K9i6hgJr4GQsmpqIvZR7KCbO6Ee1i5ZYCULS2pvowWzvz7ijhFIGA1MLepFPONy
2T8XZ0hfSGgqjMVwsECFQ2LFO+NdtceAYOfJo8s6mJSXLI84Zdk1ou8tCCoU0yaY7dkOTUh1j4lT
eVZ3QAY3w+uGQhTzCuGAFI0t4lgQ40gdGaZ6VBYpa5l6x/IXl2yRkNYkjurXPePT1mSpIArOQdVn
s0HDWno0NhIQmK+lz1rfhZIW7OHd84U+MSBDPQQal1BvbTyDajkABnXFfYaypdDMzK1JzMc26JME
ioq3UOkwxKZ2Si9IFgVG5+2U3JDM3Y0wK4wZl4b0WIpZckcJNNoijxdy8/1h/rrZp+qTAvXcGXOH
RzRm9S/pTB5AE0nHq5oCdp+oYs7Sqo0Ef2iQHt0v+9Vi9r0KvFORBzEnr3lcAJUyxb6NKjcBpKGU
4QyypC3KVJhxQ/aQyg4D08imy2qDwDV+uKvkpU/BzfCVQ3N9Gf5qpoVQRA+wwZ4pxSwQGMzB/mkr
PsW8l2PsCIsbZ12pv8C5A7x9a/vlffV0Jp1n31JsNdcnONGQ/8MjD9FqNNJjex4PyD0RZUi7jFh9
sjBbXWVHF1RZWKbbZpl3NLMQFbSJTH/5y/OF943jSuQWr2NZvPeClFbj0bGdie3XN7O1NacdbJEG
YcqgsvPHElPfhME3lt4ENtuWC1JLoRhT17eWmpG7ndgqY9zowrkozDVblRAHmOP66FfH5zQJNA8y
cbzU8pPP9ee8u+pbMKXv/MBzL+vvMpb0GtGemmVl6ur8ocQxwIq7u+Sgv5u344jdl8eABnPdSCXP
LJst08nbU6Cprjqi0iQw368BUs04/Z+uv3tqf2XdVw4IJ6KSbjKip+5Nl2v4J7pzllZr+AEqP4lu
VLG+M9YbVyde2b+9TZbebO3/s7rxpB55xRqsgrts0y1k5u3cUmtJtX+B7pqrgAlD3b4IAeEWacr3
Mj7kQu7zZa4fKaYeKOdEJNJm1r0v7duN1lsNrTK4G/+O6+cyLYxRKJMenmrY5GzZN1LnSE97+0ka
kPZTl6M38nYjdJ7SN4PSUAnNNS0TiCAgI15x+NfA1nBJpd1AgGdt8VCfseYEh3vsN+OFP2nA0vOl
40ifoyi1Qc00Lef0MIF0200fv6T/jldpyn91J5GJ25uFBdi2WY36ZOXJwp5K7FrM6PXpW9yzy+X3
GMi1b/1+FwlaTKoBoI41NKl8yOdH0rH7mz6PUwFAWN82bo2fzeBpxbWv+OHkjtxwcZKalF1K4SP3
GdZppXkOpdkJYkHGWqo7uig52ApHlyHyhIuQCNrzYJETqU+UKuQRGHTcS+C4IyxVbiDdv5EZbPXX
lJ0zj5ROIIJxnBIyyZhcGoH/QfALlK/OOt65RI2G9xRN8XjHdy7Pi/9kd5mACzcGPFcK6WyVDR4L
mVosG8CpjtI3E2b1owvO5KQqcvj6xw4OAM8T9vNMKQCmkg43/nzg0WQdhxuLhJXT2/HGVZVpR/gt
QtSrliKPHz9WmeLFd2J2HNrRHbburNmiWPt3pAZ9IIoY/sEE0AS0IdAb1vFsbJE7+8L/u4OWPdC3
MIUv4kGoFaK4TOop1bo/QnFbYL0edpV/lVAd5jAMFYJ8E8Ng5tz6kHRn9aFKG0L85WIDTMR/B404
ajMeZHZ2FMFtkpOOiPLbS6PHyAFWHxqaVpiCupceBBdUji15DxTqp62hjoLTzG1AH5tiEQ367a76
Xj0176d+VM8LezbtuQic4Fmd94ztDqDNqYG2y//7r6TH8g2rLK/yrNGWONxCTaHenUzi3eV/MutJ
EG3vy4nVmggTiqP0y8T9bF5o668ohGJbLxhanwNVMGFiXvTHcYa2nB7M3QeSsZ2b1TO/RNOrShc/
OWhZXcNdOKYAhHQjLeI5wgKqk6rNk20Ovndu0QnpdQZ+IYff7CsvjAi2Q/S0pf/eUZaB/nfBDB12
y3YzADKrUbl1EFSszfbNQtUxGQ1VCdbfBCEg1ahFRB1YBvdQGhZ+YgXsChKM6VLZ+g3PXe6uZZoZ
/dl5mYrZQJoZBlyEHc0EgaVNfNaJJ+Ov+hQGsV1Y1poTRXMSYjLVQmCvDq4BHQQT1rtps0MLn4FR
VIbs65DnqE5B8RAcxDK5aWIHMO+EmCIKWVMl3x5dugvG4emXshbu8Nh18REbGFcKR0D40vwZszoc
G7CTvHLXoYLibN1xWBz2OATJV25+yVUQdfhYnPbTtbsHwesnn5wyXDwFzDGzrQj8WDkK9PM4h4Ca
+V+KyI4TZfmqXSc0grbcy7MEQtWl9R7D3U+JH5DXt5Vd7R0z9JxMBQ0TB818JpnN1Vw5WRUIPenX
AMhN9WSKPjP45Y15p+Q5OALEIWrRQ7cV5Cyr2Yac/6m/uGVdCxdsjtZhJYU7xvyxK8rTj7+Icisy
6/mFHtrq+FUGXhhIlkoklaGsVTxiwZ4Gd5vEiipRb3CIzASloRYMBLk1AqWuOCjzBYbyysArsTHk
eWrx/FX5xEq0b+aBFwPtHCaxOegJuFcp6GJu/FFVTWdbbR8j5MY0EVbwipa9O8J0Ew0NRqk1+mcG
sMRSyGIyhj3umpGLJ6ioQWrCdw6zJ8SS8dKMonS74KjeP/RS0qUt2U+vMl+YU4A32SAn6+bIdNDk
kUEANTxmzXezfQ0+3XGzPi3gXhcKVGXPsNKILBUp9+NiBCaY0kcmsNsj2ly6REqwKCu4vPXWHgGQ
kcs2cH1ozkcQkY6DL8A83woka2hxEnAgcsvboLsoRnMzaHNAn7RW9qqlAbzkT1w48tk2zKVmVD3P
m4jwEyIYnLCCQ3BJLgN4+QfRcVtHmwJnCy/PI47E1fRuqZtOX4khY+/tTmK+wMe5K2VEEilZPw4d
+r2Hk7sxA4JIw0aVIxOLsSC0WpqzhmNzx79THixXnakif1CIej2Bbt4ydSatLgg8gjEwsALCcV18
WmxLHMzcX8WNQeNicXtMxPHoNfHfKWqioHNY/enW+KkKFjX0KzN86ttCPm0xZR3wlHrblI+T3y2z
yB8QMS4LGo/1zQXlcoEtNJ+Zj/rEuV77VVthHuNcpszCRD3EAQ/VGYQa92BUqb3LCtZp0uE1lLwI
3D/q2PxM8rZ4/wVJrUQxHDlGfQSf4nnOlkbiG5UAH9OJBvOqEhsLPYcsClfsvl/9xRalk7dNe0vv
RT1MKIPqdcc0jnRd76yr27vfCMRjMUwnC5rZALTaU8GpRANmreWN+dIwRNW3N9liMQWnweX78fI/
gOF0zfuicN4Uo4P4w3ppmtdrRfg3k6zoqTOosi3RBWcgR3ghKNaHlAz/qXzlEOV4+fxkdBexTxtV
bOLBC0k6Q+69LZKlGxaHjYdqTEyoVJIrREL5Cbn0ebNGS6vTw7XL11CcyGJEhFK3AxB/pyu05o1F
8HEG8OCbumb/A9AT7FLSb+XbNu+BOcQHiKDzTCy2Sur2LyQbtn+AIsrEKxjAStHk6Zfi1hq2Ny/w
4AH/STdYMLSvlAW85gNlQBaTj23PY56jTQvufKDxt12yoK3xYVHCpyqvxusYwqPDuyqhrP30UhCo
rrb6RgZEpRZmPpvilsABzmfu/Z2J+mbRM0Vk9AnSUIPrlNXcYYUILzQpxUdGoziCigpCBCv0QHpl
MLjjhbYQFID7gIIsGi7GHxes+Jo3ayOjkAkWLS5hrBZeImxFVxkguoBY+0LKP4YW94upH9EkaniX
vTImPs8h/pJNCAVaX6aQFMb+2K0K0LkZxdGDfPA3Haz1t2oyQ1tj5SAZOXEkA7jMxvaPNvs2RfLs
gtX5c5hI3Slgkr1aDZXnZ5ZBZEkK7vNM2/MaoK0t3G1kaGhHL463Td2p4mi53359f6XrQy9Iy3V3
As3/tbJw1XkejWc2fNQNTuyjN/2MMJS6kmQxV6DBXi/DWfnUvuVYTH0Ke9/AZt5KxjxunFQtsaMi
AQzOWrvUNARNLgAEtZsWHqem4CdLZ6324MpE8LgBiupGQhI3OlkF78UaTUkyPrObfYlxh87QkmHQ
nqo8nNxfNEaHMl23wtXkkJXsFaSV5EGGF9lJP5kO/e0YcqxgpWydSiiCzdceEamajZCTjp0FiJ7R
wPctqYqg0pxVgD0CG66Gud5fZezBqCAYc6VQzZ21wEfcBkdPSSmqD5xCSmYEdU5GwuY5jKZp3o2P
CKge9Du6rdG1meyAqQ27W4qxMufb+osF9xpM8w/4KWxzArJXYoDpiG7C80fQKLiOJhC9R/Sv36Ba
0p4izHDmZJ46vGNbu3omF9TuDVdGE2IfK1g6Nt2f6fGwSb37wf+iH73MY9MS5PQssTvjj7cfSXUt
8jf9ozD/D9u93jHlpLZA16OOA2XA3kQwo2mUsljcTqWWC+Jc0Dos5qSRzvNgfpd2gf450S3IWKwo
Ms32h0JaROdTNGCWJ8gA1lsXgEccxrOpF5xsZYpIkCPKQbLDAdor3aQ+axRNgZywRZxjAetbMQ0q
eweT0Wvn7RnWtLJLYN6Ww8A8FMf+Lkz4BZIC+7RoFyWZWf2kaRGFPwtSek4vfeeDrQTxtN/wk/uT
d/3OagTSRUwfRWwHfrZaWLaukoFL2Cjm+KlS/4eMcOQ/4IEvCfbH4HOrIKysTdFSvbVnc9oa6CUr
HrBxumyoWXu+PWPuEvnqrcm1C2QLJV/BvKR3W93grH7f2xELcwzLLvrGypA62l4pTbw9AufWsqi2
IcDvdLlT9WrSzuYgayFgT1PrBPfY1xonTKvRcNd80ILcx9nBdjrMynBTQjnofGVOm03hOKbdlTu/
TA6z7BimTMz1XBmTPzIf0AKKsurgvXMVXDFWdySP5AJvknaDwJ74tPZpAtmlb2Vej6w2z8iMD2bN
NesygHHMytgzhaFlpvsyyhnMWhXTjMyV1KIRJttrqZoxM3NTDvsu0EIs+2RBex+CYMSmOa2PRopb
qTI85jliuQmb5mB7I/WLUWzpNmzHLkxEUZgAhGcl4k0a4g4R3vlbfn6fKBRJgdUEC2laC4v+ITIN
xQkE3I4XNcuJ/we+SmtDPQ7gEAAiKCyOVOFHvYDbgi7vncX4k6suS3SvzgaT+iwv3/0487Fa52ys
Y5tp1qrBx4t6A3I0K7uyfwW/PPjc+L598y8b66QCuEsWplK6KRcUMorhbOFKSE+ylFZmb4lJ2PBC
W85yrWjLu+ZhURPyCbpAUsN6ntDDCS1XtUsfuCkXOs7SxzSBJd0NFVQve5zWAVAhtmaV2jSrCtdM
EfK9DBvLwVkBx+rgXD3zhvqvmedYdRxJfyqlrOkxeZ1O55JShytsJZPAGrcGiiee+5XyHVxtYKkL
NWNIfsGmh+z1vnVSCg94TmApkbdwhCgnWxcFpJIdH348y5Qm7ZpUet/hRab87b9hOfhqfGO7W4Ez
+kedZeb4MiaE7fQ8S6eMtzYOxY4B74wibHjMBl9vkIfH9KBzDZXXQDh9dYX8WLkD0cBYNoux+oWm
h57DLRYZVmJ12OKAqOCzhvofr8+oGQOrehp6Ws6vsr7YMSL3WzHb9+ECrM0ZYBGtaPKe9t+cHeE3
uetqGtP2YkyopVgQgCUcFOzB5vElWjUA8lI30sWIIno+ZmnFLDL5tJ/RANXcYOXB0lp/8SbRxxyL
uSDkIHA4ukgEwo/d8n0wwa31T+MfWXitv3ULwqbtnHOj3/S1cdbk/ZCbQce5d9B2dzvhhdPObyKK
qVXIZNgX6oHqVMD/i1G4ADU/nIFdgP/F92QhrIF1wFhoRLHvWTvuIzumn2OdI5/DjYBiI6tuHCCP
pYDaj9NSangk9JQZrcLAnw0emWzDlCBo0hRPvgIgjqS8txF9uAsEOPgtbzlWhEOG4FLeATBkSMyd
VYPA3z4rTMl6RmOWxbr5nCDVyx9BuVPbUijTavw4IIgI6EsF3PsibArq2xr6gvd8SQBwooeR0TS8
4DVRn2KZb6iiWKZanaKo3qxTzJBDAqbNu0jqU/oq5eblrNhLhcl6ihPWGLqq8Y6oE8VSDdV51qVK
lqpE7iRVNCe4iUtEuleAFicwFqzC9LECmF/F1lek7vCQNneJYi+HN2n1pYtwOMJrW1Slu/g6ggXM
cykGCg0d1tc8VCxi3wk9tDbQv4bjVX68zo6YUTw2fQxOmUQTmZxcpt7nnF2eQo7NHdqfwDHD5WPs
zCpl9DQIrF0JMWy3QGbiursTf+VLzm1Ytvyx0qzFBat/MHETwAZpApKek0IKRpdwN0j7mwCXpSsU
maqiUstfZihqLboW9VJhCQsuF3G7iBPJkZWvAPCduTtMCWGO+iTNJesWuTzF3QopbbddXPpXu+nF
58djJ0UzN9CU2LEpMfUih5VuTIDm6sLE5HDc5l8+bhMX/mGsX7vDXj6cObPyc5jn1LVltCJbPQvM
/TeMxHi/3PvrCEOFdZLnhV3z2NzvnvM4zoHLyYr/9MxKtCc4Yl5NcxCiXmendJU4QpcUJpPDgUMo
+bhvv+RYHwnrScN2Pl8wkUXdnQkySuMKEFTYuVkeRajfvDIekMwyb1nExJfNU/iyUU/K0S6OMisN
kwR6ZLXeCAOpPxq0Vv2hzSfD9e5FQYe9yX35i23bhiH3T9DN4n3pZ5k26G16TRTUHMLWO8X1ZKNM
FVuilABXpYkFhxdJu4JuLZaoYJgyMWlDojvTC4A3pS9RWfQkDQ+ty8nNW2ZRfv5IV3eC5kMrqTkB
m7o/0L0MPGhw50yzSgfkXcxgXhuCUI94PHuIuFvjbkdIaqqTyEOq5pED8VkmzNW54g9XAZgImbe1
vKhnci/WAYVC60Usob5w3iZnrTCTiJZPFbwYzmX2gCRCr2lmkKZNUuc8z4DOZ/MfyPKNvSqGOaD+
iwOqw+H6N4DfN04r3BjHu3JvZei/mCMynXlJLyelygFzTPTEngja+Rf2mlwwM3CEh503oMqEjU/u
8QvXTt+UfjNFCLFW32pJKEWKQkquAprgVYfwd1F7iExKXbKoCWkjj7KVRHIzKwgl0tBCDbUO53aJ
wURnUkJsBYPVaayBOxrgneX+OWBcKdZmM1OMjtWWSlmK8k5n1JcahbU9JqmWq6gSDmvdJy7ujMRO
aoy2lwQsCE0S9/YoX0BHXsOe/A2cSmf02jjIZVXKoLFF4xVoePnqd0utfp5k0kJ4epkeJ25HMeQ+
7RmN3MSxHC9SwRzaPGrDnAzbHojZBpJ4KQXselldXIWGgGzAR5jkotdOhjXVTitKK9x/6YoY1fdx
4V7EhCat6Jou5Bdo46wJxp6b8ptO4+hkLMr6vgRjaVDfPVK9ub78tesuPQVSdp7gKt1cU3pqbu0Y
paR6kJicdFwxf+CFH8718llyGGgZWmFpuOq1eQhqofI8/t5t4n3paJ9WWjwR2hU0RThoMf6BGszt
iwOZuiSgWBaVEWAAdoCUnQKGhSkB6xdMvi7QPkMtFlGqQXzz7RK/TOCBOn63zytC/b5Ok0WTAsec
gRL0/omjVYXdPRB5TboAwbEw2mvqIdzdDA0l+SmKOwsTAWoTJL+E26vHZhPmXjWKiWVsLHQPSoSx
YHR33PRz6g4Ue5Pej2rIQESNgbrQnl+l+R3SFreceOKGa1IMmYbY543jb9S24KVorLSzl/4t5Mbu
QDLaX7N+1zfkQCZ0gmG0GJaWjaHViWeJHUaUOK8D5LXaiXh4z5/58GjgxKkIRHxKmR/zZ79oTjC4
y9QdB/fQERSFjx8xxPNzK7VJdibi7eCuryYZu2/jnh/sBjSg4i3wiAjJ4eyPfVUqQJJ9Ltqfcu8E
3eep8K/RjJe1KHqSgCkCFlVjmPi6fUWsM/EYhgFt04eXYuR9VYe3q7rX3WkBsf7uHHbGm/fASsFO
rplK8NvpjTEoj1pttwSTYao5bMecmenV5LjsE67O7lh0ooDkkZTq50zhaiDK2uHdjoqKKgETIap2
kwbiBWEzB/CopXy0YgvC7RuxwfX46lQLRXAE5ThzNFC9yWU5VAxequ2/JlS+UyfSVSyX9C1wtXv/
aFyijViIyHUQJHmAVLrCnp8Z9luaDzJwhxoJaLVgsrJXs2gl8gVaGGMSZVkAuCGIOO3GvlVkdGmm
nxdZzUvtSya0oE/WoKFw9AHwz2JEuydEc01rg5JA3NvgZQlKrdPcEkQEdcUFn8LAemWO7zGSVolY
WvxOhs7GZMeragzAgnp+KOyTzcSNI+zTaA35AWzlX+c4swxXogMXEZAV9z+osossds/W4cMu1YVK
1s0mPhalQMq7yH/useU/sST1loDlbTmYbrI5B9VNtLlBRLiCXpGf9SFmqT+XCw6ucCJrZ3F3nY9r
/rFGPtojDgwz1quZ5VHtWNzDNUh4EdBr50I0bN8GWMEAe4aao1WOpmeAuzaPL4e+PVcFPmIbchbu
D7x3lAO/4741kX42KSvkHR84ZL2ZCSWKnWupySfcVZ9GPyh9XiYve9COgvWCLSFntLDDLJm529re
IBvbezYeF8Y2W+ZLaEiYTzjepMCNP9MiQaTGmdpuxS7PVvjmjVAbW6LzsGRutW0ZO2QopuvZ0nWi
YcR2zdqonZ0lheTPHgC4r0nwZO9BRdU3gWbQ5MrmBkRGjlK9+h7HKXopZkwdGT+88MFNm6BGZ8Ms
5c1DycVG1PxWcLnkIRllqee19+qlkV9AqqcCxLxDooFe4PQUshYMc1nvvTqzONcvg1nzPxSYl6Jd
61fcJ9i2Zy90fTqMUhLDFHSjZpjcezUsAqUxbKKzUT5mYMBeFhfHgVamn88Upu9fRLm4Kk2UkfaI
IIWbkgHl4fAmmIJ1BibF9N73D1zNgp+9Xcj+x0OytIlZyXdr6qikPL2UNYQAbyn+U/MyDrCK35yc
PvsuHxjp2QVbjHyNjUIK6nHZNuWd2F9omuXT/tlfo/mZ4t/TvqbBd+uN9+DY4FmPEPuS75sKi0WM
QzIRz/LyrcGfL1uQgilYkN9rzypVzcP1bRusurtUMex5vApGhE/9HRPM4/3ODJCG7sJmPVQLX45q
O6nkZY86Gj1hfCosBN+WTcNKprM7aXLKuboRmnS8IjYy5OkG8DXNg9KC5uoZ8J10JId7N7MZnXZg
FTXNuzYKyfrm11wcApG2Gldkd8hJM5YmzQNho5NoPDgBeRGB/hGMnQ0iEmVxj3Dglnxvqg6z5PZw
Mv+ejdszq1L9JxRTHluhzd533Vvvg4jLZydYH0ZgV8YTZbgNHcDG2pF9jqxk2P0pczLHbp0xar/e
yDX7Uzj8hjNJD9rT2sjEwVFcQ/F3GrnjGRl4ueiykupRFj18qWHT42Wxqh0D7hPxhfxoxa44/2aJ
VjxKqIvYMdYuPajzvhta4hxDzKSIrxuTcTRuzC4wsM1LFO+d6htCJmTWrEUdMgu8NEgPLGUEqIoM
1JvCcdMRhieOe8ziaKGEkIGojFogQLnYnIS9AQvl6tKc72qrpci77Hsv1C5qE4ubZ/gSWOiNYkbq
uen1cCZYyPhF+uK0xYtFBC12qBiPCnxtBL084t5O4g5bz4EaNu4rCSmaMq6/BXMIyD9ivC3z+9aH
hpj/FLGQBHGPJ1H/gVR0DKxzW5/+9xMVFCrKvm2xK5tHX5CfGHac1NCAXR3eQTt2PZ+aQKzTSHH1
aQz0vaDk/+2+aJh6XgMRuPi0WQgez9IsvJg10A/X2eUBEKre+n9TuJ9so9lIYB8Yd9ojrJUdiLf4
m+I8D4U6XnrQanqbKSTWURjrwzieJOrP0hN/fEccdRNMYiphbiQVqZ6Uo+rYMx5BqcExQN1bADkk
ofF3kvIUhivTEYQ2FLkMVG+wRQ/ab5mbKdGcbncAgWqBpezag9e/LylfR7CejicoYf+T8nOTyuJo
kBYFUKc4ppRlpTIgLkwJ8l0AR8z3PIKTaVPKFMs5rN0YaCFgMn4RxMNe7uweuZBGE3FlNOE3W0rA
BnFj0mBYuRomc/BDJ6JpSEWPWqYU1m2B+8hm3XZi58C0ad6P7nAzUtHdJVv+gk9NsDa79bs+cZSg
5SDQy4/j3Pstpm359TpZOJtIukcq0U+Dk3ZvtF3f3Duvx0FOQn8SwEJdNWWlAQA2O4J7wUCErwiQ
yvCtkNEhayU01MZpsqMC1DgklzEXXsUWMUlOqnMR8M5k6MP24tuRzL5zM7/I5vFHsT+l5PwvZKD7
UZIp8IH/mVkbwIcDhbkTl3SY5zAeAhI8pcOESEJm+AyZ+IbqDFkzCyLnwKT44pfxD96D7IFHQ7gS
tyD0V49JWNJIFbcTgZaRNAfNY62LDpkuUR0QI9+YsUCQphzhIpdpBo52l09AsID8tX4wvIbxRY1b
AtTxvIhirzkKJV1WKT+evnIYSR246q3wFMQ5yiBettnNDg3w94Sg8wKauQfQx4Z7/c1ixhNE6iA4
REwHZKi97R2lNx3IiDl7RyiBcJz0nhi1a3S6JRi4Z2kysfjEm3EdIdwVjsMoyZd18LjxvESWRpY/
7pjm16Ckmot1HmVoAuroDGrtSKJXud/N1pwbiQhCtnM3OuFdhi/1TxvzOgruSgR4T1hr/iD/yedX
J+TEy5se7c62s3MJdp0becmg6dBU5+6mVh6NKahrmuhdteaHxVqubGbRBese3QcgXZf9jBu+Myps
Eha765wEApwKjd4nUKnLUUKPWxU3rord45iaQ7hYVWqRiDAI56OY/LLmbBXvynoh0pIEM8SN75tb
Todd99dF4JCoc7BCv5WJp4BsPfmczqh6H8ZgDvVieQTEul+qBc4McdXwi+sCMGTp4zfG22gaAkc7
VeH7v/nwBkUFaT1jLKpu44FofqYG1q1/budXs2xI1l3cO/VIFgomaMQuZQOCUlIeCzF5IiFRArwp
+CCCFowJC7z58OIk7fdMEpm5K+M6jF/QgzTQPfET6DgAnX/aBQLpN9iLPHwf7hPlsL7BCFdv1hXi
4GsF1s1Rbzg/omgd41Tx4tEW4AbjcaM2hEdeK0O9DeP4nf2p2lEYBOIVcVWN2tsqZPsNCQrIwBQw
9kFvKNTLEaiJQ/JqJHST5mWOW3Js38/n2tTrPqErccaz4JWbdoY3qLI4NH79sOBQy6bOhXGyl9qS
7p0zdtNbxmdxm8+PlNXW9jtyvG1/wr9cS5m20qNsqZnEdaw91BnltA2oKJq56JcxrQoHJgUIYSi0
cIP5uqHomdlP7WazZRsNnqoQYUzYtCyIOsaaEd4Vu77ZywP0ssYma56C4+T+DL64E2kb60JbKx83
COPd2Ez7zOf03K6ICZIUaogLl72U+FlSsIFzZxikZ3QnnpyakzQ0UZF4yangTJkzHzMTkVGi1D8r
hxuXDFhvv1p3zTtODt76+3PF2VFVtVrClRQhXfJmQj5LvzwmcItq9mYG+zVsLjHyy9RCMB8D2G5D
R8vQtg0bA+Zg/nLmvi1c7T/gOPc98sjgi0jt5q4hnm3oiO3hL+o+FMf8KkmreOGgkEMZ6k92pg9f
JMIE4/K8Ny1gIAlFmn6hkj+Ukgsfkk9WWXYpJKf41cLCKBG1ekYsSjZ0ytDedfwkTM+7q818cXUm
V1KjUcxrk5u8dd3F//pPpbhW6gw5jfux8hTFfQiDV0HgOU/qsVLhynRxTwUmppYP4OdnX9QqtgZ8
l0IYVv27ikU5NHGYxxGokLRvnUkNiDjnwAZjMDErjdZ8CgBUEm8KInuaPi/dixr9294JIgdRlU2N
tJ6pnQNkL2b748cvaaICCqeI1tpKnVxmPNacImAERYythjRsjuB3L1r+MBLXH9UsVIZWHPXsxq39
4hzP8bAyWFF0DG8umKPS5OWPi7lDvjYpR+bkUhIiNU/Z9pmgmAsKqF7mcOuVIhwda/9LhsbXCQ3x
6ZT25het+2db1lVCSSHQxh8ZPVLXeJRuD8aQdk0KpJfOJ8tvRw7gy7DvmbXlICZCN0yZNFMuA6GD
1SrzhbnG469rr9sGSuXKb6MVB3C04bM6EaeVq3bCdyF3N5a0XMyqajjOA8jL/jaHHHzhHHvcLdJy
E1v8PyWFjyCl91mMxYJS6TqiPkdr89goSY0xPpetNCPIZ3AkAZeyry11lchIGA8KSmKmfskiknV2
D0QBiXrN1U9RBuhu9/fXURFSgJJfKiuwSQHfuKCQ1KUnCPIYdyuiuoLUEapF0eDLRiP/p5Zt6nsG
llXhM+6SClPGY6BzDUJMopvCxtQtzXksLldDswRgAQ79gWTTEpPX38xQOUMtX0TXdRt3z5zJ2bP/
cyOYMikWaZoCtT4F+rKnrJiGGIeMbw+ydnD33dnbknfdOqRc+9YU620r2HYPRPeN95l1jOP70sa3
YRf8YKBVX81590J/PJsKrqi0ulK+XrDAzmJgkZWkFtnPp+S+irX2Zrp/YSHFxn0EG+2o3hO8CHJ2
FZSBLzitP0HJM9jUbe5rEjW0KctO71nRgolIxLDuKNnP912hdHe6dvXqUCqvSdQCz7FmZNt7f0q6
+n7kEWCWRkkm326rJATNbrxR1jS1+huGltyhbzyaRnIOlsSed9L+7egx+5GrBiZzDAlfOG6ul8pT
fW6+uB3xn3ORyYlZvES+2s6GTLQmRU+GdilCDZ8rt2DwNvOUrbneBtdZfMq+g1/oj00CPOtt638f
1plNMgFIk3OR6Bgz+NRqVM1LtVjNF4sDi+Z6BjSCjY9OJ/870Bn5JfIOBAJyGEvga0guPJ6Dh2/q
o/pWT96VNcki+EcG+dRUC/mxNeu8K6xJVHlvJ/ctas+qyr9yFwhr4BzvI5rmPCpiUyMADp7fmIGl
E4mIGyunvb1crIwEvlEhNALzvzKjxckyZoBbptjh1AaIZkg3mqtsABt1gGz4QnCYZtHsuYsmz9bD
V9q6a1rI6lR3XNtpGfcX022Ftdm5HDXWDOfc6yQDU73lAGXmfjrEamggMzAxTnfWLGbDMmBdWbJg
bFCdhRszA7LGrvewPiuACYQvhONpJXTfXyYO5MQFTNO/7Hpj/xm+hnnYs5uBWtuXQx5NDRNx81Qv
6AXYEPiGmpx+x+12QDmjDz42hCHSsBnMJr3BwnaTbO60iq9Jcb3dByLsIXLi9aXs96kmKeHz5C4x
ZcYZuvuPK3KUQxj9GSfazWSiQ2RuTQW/EaLLZ6Z50oPo2inMev10maDCkXZsFXl7q35uniNVY/pM
FS4FtHq8Mss1OCQpdqK1VCaXIDn986aDwIlw0kM0c6VGG8sHsGS3NI7QC4gejLjARGxX0L6Njnfo
tGcYwOn/Ao41l1/lgJAS1fFwvjCIMEQubIu43/8eqabYA/TpI/1ozkW+3/ANDD5mpAgB0U0jkT1M
6tKps+mx3DWRhbVWoNNfwHbrXKrg0gCWp0VQe3UzRmXsDj+3DmCQxY2Xe6OdED6GZy3aru/1cRRv
u0499E+TonFq1bmZ1ecZ7b3pwGvIiL17kxlSU1eC4T7f6rqNlp6pvuO6d74lqIgT3xVFE5QqBvzO
eX1nLzgBbdpUk5T6+gFns5i1Ux4l7KJrud2pKiR69jbdL1SPmSBkBNnAY620vu/IhP0ZZrx7wP/x
HEKq2L4lvo0m0jcmhLpgnKXi/QFTf1pEqRcYTfbaGtrEQvo4pJp/f8o7E3nQg/bL2Wg8TpUvgl3r
2nUfbt52RqO6v53DFL0Y1gTmSycyJL06JahbntR4/2cqDhWtVgtejqd6hLI4A2lXlPoicredSxoc
OhfeYT7VMU6lm94EJ9RAlOizXTdNxvpqZJYiuWf5ZSdb3TqoXziNUvNh8EMQCjO5pO9TuLNndAwZ
eecot7JT1O3vy6jieq5DhT8HgPPTYcoX5yTtMSjPz7pE5mvH9/IFcODy/9usLSdwmxeTZcG4q+xT
9CF7cPmAkc9ZMmC9FyElSfDUjhjDi54gRxTC/ltowdiN+FY/aDwFv2aelp5WibnLFUgV8yxMBsos
fCZZiWa8jZ1mPQYb3CG55UBoK7O9kRo3x6rOpNreouwxhAo9z+SWVQSqoAJ5TE5bK/sxBAYTbzlG
t2Ya61Wb/7MglsJi8OomcmjZKWr0KA2bS80kRaNz1aDnbgu4oVdkHhDCmK3lvj7cUdciY9GNjp+C
5xPNr70mbMqh6Uvd8MFc1Uql0TvPPwLkC/xjHwSdPfroCjesa+2jPEKmfzd6kwUzCIak6cZV3aB3
b7G0NYW6SgFLnAaIUmKLrSDGnf97hX6raiqRErxRsr7wePE/tQnpNcW3aqIqqAC5zIBFHFPsDem0
iUEJpkilMu1jcB7kYp/DLpRiY6HEZJq2Y5t+soF4eUGX19EKejg8j37rzZlDkvrYNKd9l8Z0icB9
BmxnAbJJvjVdxcDV3VswKuzHY4iLxPNrkIHm1i3Ql/6q/J6t0z+TbpUQ+/vuotKn/j9KE9e5UVEJ
xOvmIg6zTLdh07Ec01s+33FaDVJCLfbni4KQBQA8YEBEWgjls4qn+xSXt2N0DK2554g9kfLA2Y/y
d4sCqFdy+Q8QIrlJ2T5xJk77JIOxZV9G5afrc/47Gdoisf07lfk5t+/6OAyJ0qsztUmmdHoE046c
IHXidqR0Ex3ij5hdwe0YpaH/QDBPnUXK066ZH0MCchS6gG+3lHlnK/gPeUN93EBdTiU1+cM5IwnF
F8cCEgeyThEZ6dWqxiWGvQ5pcJkQ5b4zv/QMCyzeayMdeK/0Ex3vaKq+sPMsd+GBrsnATZySAs5z
Ik+t5fL63rQcrswyPg92CRWXso/tCvxvt8jM77VCloSpjCdoJz0phIn6jqGqtaedZZeVKH7xe/Je
xSOUn2Wr8hB4LaZwfRMphrC2Lf4ItFPA7dXoArinHXn26GvAPqt3mEnU4owVln0XOHtskM0I7YjA
9BmVJgXsMPR2HR6o3w7427mr6MF0q65vMYzzI1NZYx1w5HQq+XsP1CpYVevq9PEiNv4Qd5TCpCwG
BeimctQPvQQ3HaGHilQN/9hwHlBB6IIgpABHqHTYrsvGTbLOEWqEtiR73F8MxXg7MbRfKGFL/W+b
XTWSNRLGmlVot7kVQaT7RJiShvOm15S5pFqfQN0/g6Na3v0LSn1c15ggWPatjHkfQwozaS3kNEiM
vBN7VQG2mC459eqbLuSWxSnClVrsM/IyD9fPOfbVU9ZXMD7ZEQux0lQA+uWEyGWwAxCpk5aL32FP
+U5mx1g21k96Dy37ylEqi4/XQrydhiIrKWbU6GVStEb7T7qj0MYqX55VAtEd1tucIAViNmOTx4vr
yFgvdvMVpNsJ/rZRs9KPeK+n2XBMsL9qkJDAJanuWl2gKuykRy/762d9+ySknvdJFjvu6SDV4mHx
Gprd71SCpRCvb72X2odb+PC4tyiF/rcGr3kaQb0Cs9vafuH+zIjrXVYxZsexPLFHAegUPjm0/HHp
qmtFv7cu3wsgY2UckfvMT7/krzRMaUCeMQlA9by8eBRwV3DSubKcrnixBRMfva+7jjgFO+tjGP3Z
hZU3kf/apFoHGw59CeVrS+ebYU6eiHnrZj7VARvcS847p3ow6zX1wQOgbNDeGO7BHkZpSyQjHr0p
0woBCsjUMYSE1UajBQbfb2I7Ozuqhnqh4N7HeEVNrT3+XUJP+mxeIMPHb7Fg+DB52lA27etfXSVI
YXRgklXeEUV8z+82iVjevrpNlK1YotnDbJo6nJtc96iu6BOZQWP2D8Fr3HCpgYTlTOsfYXx+yPh2
Yc0wAOh2xRvffoAECjPpWQPfHKjl3i+va6XXAK6chAT85s5kY+4vV42y75+tHHuqi0KR/IrDwBj6
j2a+m1MrYSsNJgucylj17YYbw7NqDjsmD3q/bRrMC+W/F8N6Mxar62L4HWlAy+hK45FZ+UM9rCfj
Pfhm4kQfpBVu5eMXiesPSwUavMW10B3KPO4U33TCaQNlI0wyAo72D8mbA5soZ1m9gdvm1uT2EvoD
l7wU4M3rcoL/oUMYZDv1l0KgB4xXmLakABu+mSkPnLEasilE6igcOenkFq/K+x9t2f9bAc3Lv6pD
XRefbVOFZjm8Os15OzBZTde9Sl0XHM16W/kcUG7RvdqO8yhoJgmTW+LZNCDWGWM4oHSRLwA5CtJu
F+wh0IGNB4EZlEPMQ7Zh8kaQnyVacp+4HWpcLZaNpxtrzT+lyRqBrw+u+86Vp3dbkzGgzilwdKbn
BvNkFJPkvuEHugpQfdMxCGaUjxxogvGlJMmLdSBpJiH3mXEtHfEDovF4QA5sYUhC5d6t3sgglwxf
uIfxmTILMW6RtM2Ec0XyNGEPdg7+arikdOkML4+4LL2sL19FFrgSkulzzlxVHn0GF6nmILrrUrmL
hofJloVRe6qXCJ5jU7wGVk+hrH7KmnssBAVRtpz5pr1QzzoHtA7r5j/Mo474673Jpup86GYFlTkY
A6kFLA06JLn/PRBC3mYI8vSRKT7qZedoI04BpE5uv+XRKoVzf5XCmbWION7tb1tdamWOaRQOE5iO
EY5gqisa/wdmueZccKBfEOcfqI6XsDJTSpZ3mb49C9pEPyZo78aa6v97ZiTYvNeCF4zfHr5J43fW
TPQE1lu9zzthKMdrUUwDgt0Zz9ex5IQJ897XRNlKhFZBnb3FFpmBRTyQkBBAHlE3CQAknPeMZsHL
rBHhmgVd6+adx5Z1Ptpy4gQbduf3lef0bIGKQShf3TQR579dXAsXXltV/OZErxIaHpPbzBiPjHmX
SQzqkBvom++eYJtTKuaMyyz79KUgavPCWDTXD39rBhx6H9JIrhjpgcER9FNW/dHJjt1rNXLs5vxM
CFaOZpobIWa4THiHd5qC3hI1ZIp0Zr5s9J+sLJlSt+hHsR4jd6ZPiKuIaJZWwM48Gp9onAmHFPpt
zXRo397mKpRjq2LYq6M+G7ZjcsPaHXhz2rt0W/0AcRWkTwjquUlg/YiG5QzYeQcm52JYAfqSprMN
yDxYfx7NZHmWqCTGRShkCPUjcS1hx8QGEEFJXVWo0TGgTgTTYIi53Icl/6zVAyiua3/uO2WkRaGg
HIUI/FtiAkdCHv0iKJ87BM2E4OurtMrUdgwad+pzqRwXdh1q0dU+1cOddU0jZE8hPIc5Hr4lC3I7
/aXmTqOUJV8HgrcZ0jnNPQBd3pnAcA58EawsQVf9EMlTue1AjCa13Z/faiqGu7iOzGVTSQaOFBWD
Pxu2yEOtE5JeBLQR+xHhIqxEp3StkD5o5+aWPY+Pn4BtaygMwTf3+9BvKz0IftdDEiGAJfTmDGpF
uADzF1yMmonbevlSsAMqHlfSJ0kWREdRGSZd7WQGhu2oExydimeMiH7Evls2T/cR26v+FO9194Yh
VaGnvW7PyF5zHmqdHuH33LS2JfyWzLM4Zvyx/OfxIJayxwmG2Qy7YkQUaG0+oMFclqrEv/7hldbD
+4kodwbryt+TghR34HbLGs0VT0MefRMLRagyftL1OqPMK8QLrOSvUDL4FHC341PDMXjwmHNPMYQX
EzElgNBzYCkoSaW6v+yUj39NT/a0swPpDYiVfxQjr+xKw7hLLwNNI6sq1lfJ1ZJGayQeOHwYR/GV
c1/h6zBFgYkqF/Ek8OnG6SNflt7/ihU9Hg7lYxnKUg46/CyJ1kzPtz/urBtStHyFulecnlMW64OX
gNTxf6DxxmE57KXIJParDI/E0fOFfcZlz7ZDNKcDq4vIWeN7wQ+j7cMaKQ7gnay2P28dUXy3K+NM
gJUrLai58xJ5t7oqEoc/Bxtc/OKKf2WKBrj3I4nkBd07S/Pi50QiSlb4s8Jn6UumTD/xmw6dJzvh
lSjCqKB5BAyDUPLt8fGjg/dHAjoR9T3/xJcIGjdiJyk5bV8GN2ZzTnEAPQbfIsDFF0T/UXJhD2ki
nV75SWh8mvolB7oM1FpPOziA3Bq29HwMWAWQzxnLI7FKjlvtMVolslK+MwtAOwQs8mlkqCiPKhr7
IflLtcR1bchZ6QZXTiEBkoObueSVqM61Yzz4Km94RHnorklIoP+bwhMEh4KD5/qhGw97Z+S+6z5g
EYQmQ5oKjxQ7hr+GOHyfIPskBwotEExMXz76zz2ekzfnf7E98KJbWCzzyRETtkhzB4jdq+MRsyze
8806+HPp1ic1CDi356mLfIcqzljLeDqyUYPSH4lq/90UV2bVDSAtXA9oQ6BpVqYuF4I4Uu2IYpED
47JUGh3Wg/IQmhneGDEdoGyegwKiqYc4GUkEZzrK5Z1qWcQ+iIFQiTwZKwuBdhribWE0Ux36o89u
89+uVFi1Q4JaGAfnrrgblYGrEdWtExh38qLhIPTW9JX/ECo3hlzJLNub25KfLopB5xASxvjUJSzC
orDSzn3pdOcQ8ekz1f7LG4h3hL+zFuNAH3xSlnXdvR74r3+n98Pd/ibmsz7vVwyV28eyX7gR6YYG
U0lwpkE2P0Q9dd0QiojC/mNyKjTWwUpXnyUR+U6aJeafXgvi2O0BSHksH4ftgktmE/kwZwNvwwQ+
24HqfYHV6qNIQ56Un+lplz6EB8XClakaJK/+q2Nng7WiYKnu0RGY1XNuzSgojeeqCX2eHmHEYqVT
x0p0MZ2cdK2TZ4S399R3Nql8kGChG05g8gYv1FJdctXV7C+Tofe/Q9kQmYJZHSsHoJEEV3Cu1mFs
4FXGVGC0SKDfhHyuR25JdiXNtAe8Vp92mcx2Iid6rg//DG3NBskODXuvXesx3a5zQLUl+re2kZUB
Nozhg6Np3HJowYYEiXQo43765EBpQzWgaZTPEO7DQNUArBWErHowGCu28aUlgxZT8ERTCvX5U6/0
yPSn3+I55UXuwnbDs5FbWtMWrHn1jdFcZ1/QAB/fXkIBPTeuk3PHZ3PbE63FDDqShVo4cUjo+DUa
V2kYgaM/Erx9qGEYDS8qOnTXuUniKnOT/+vutcZ3d3EbiFt9i28OFOpICgk17n6Wd/kpBOhzJ4+F
QakX5+JazwqHnqBioi+5YpzfDHqDSyQg4Sd3HDCcLDYISxNuU+TXdFRyLz6wJpLgnS00UhgaKpma
G1PBw/tbOxu2wPxt7NaJq4MmPqjuKOfyAF6jG05A0GJcg92Q8oRAkoZ7RE5Du4PgOazWCoERHEp9
kDC5zY+yE+6f5DnsculA5aDqvDbqIiWWAQPf4n1gcEXoUQ4clL1LX1eXIm/DzOGwOVe5bXV4XL+B
dloUdCjpR2YQ585bo00NkmhcP8CEcgvYf0ODmct9FMx0k4SWqOp6JVOTj/hOmS1qkogkxoLyssBH
SVz4vejJP5k3NTyM5Eo7u7/BQj2jGspr27gBchl8xDy79/VObEy0cu5SCKFS/bQKfCttg/utJjvo
orwN+x/4nRUMyEohifEtkckV6naK0cWMBGekRs6O6XjNS2xNzJteuEpstClPc7r8xw29iKe+1cMG
l+MHy4W8wH8sLmYIih4RlHQXOaIr669EmqToWk5MULQyxUn/Vy2lltJQD1DoLU+iLZQ/2DewiCKK
Ci9z6KpM0DTDz+SBVtDREa+SYm7QqV9xKJQbsXpRFfh43Ipbqmia1JE7ob+Xl+ksdE4Y8fmTn8SJ
kYKfPageOwFdSBRbNAgessf8xb6rRaob8yseJWA6A+hjuM2Nn1cU3b88ud2Wal6aQwkz5nMYnt4X
krHm6XAAzcg586SAdjGDRJZc722MlBpov/gVa6v/G7b9V8r8sdP7FCq5robwomPTlHMq+YEesbgC
/rqJf3aMONnZOrvh/PoqMtDw2D7DCx8Rd3R2Yth6y3s2BISDMOp0CC8PLY9RdkIrtmUUyuslxXK1
b63EpWZTFX9jWwkqKEh5x9eGGu0UzT52zylHVkQvLeHMaAPmBFEnPNzyrDMyKXjcQ0u5hsHN5m48
Vo90yOu20VjbuG80BxVnS8sMVSthBlQuDIHCxtEy4ZpE3gm4WitY0kvIuRqAktp0fPBIMHBGppV0
CxNg9CHyntvWfvkRsEP+SrOQ11sBBMXZwJEruUX/l4KuKHhq2WkCzGe+cadVZ+I1y8d7IA+GPj1z
AAmMK6eV/c7uQVWyHbokYxrXESa9s45kiizJQx97p+zfqAxLHFBFwr2l37/0DAYXIZIxN5PJtvFj
xNVCcTKhZLFUe1w9c+rsGN1nmBi6RLOf6EkweX8uvhk7RsQrwTU9VeL6PSLDYqIzMnER6k2T9QOS
knNvQnNYOygyLnIuj4mYVshxQtGTgMvr2y4UQAnTWLNU7l7ScJO/uDS6T/J/lSl81j4fL+xI09RM
F092OgN4FFtal50jEvVLZhLbieKm5BiiWYHwfH1bS0WPhJQWTHYPgFJXdnTrylxMgxnRy/K+uNoL
pe3Vw1f4u1zxnz2dr3pVPPFeLWzU94fU6gUpArrD87PKRGr+NtGMMuy2jD9DK2hOrcU1sWyJFMTe
36wNqgUyhdoQtRpHudq9IUbxoMHsBMfB6V7e/DuVfGs+AAOPOwiAuurAc7r/D30t2Ldx9IvyL/YF
Wgk1/45cP0/WWP792fks3x56OyhJK5r7ydk/AklKIoLkLmAGAJ77OVDGqVJ+Kd0pHGJCQV5VYOz4
kg8p5Eq7TlJVspBC8iQMwrPSa5Hy5W27kQZxYMKfV6hd+EylWARzEwVWr1ydvu2Ol6ntVBbV+K22
oz9F1lrmGtg42xOiVKhKfjwQJ0l/3Zm2g2clwtNaFFLEtB53GDsCJ/7qUh3wnvdz/zZDJWKdGYqR
IJwH58kqPo7hssEn3e04GRZ7VgvJLUgp69tiYYdnjuL4VHiFUkyZpwvNVrnH6EAPnT7fPQpSj2Uy
cIhD0M3oXHhyhH80ijv15Phj+6jusowEY3FTlkS6WQcUK6YrsRiGdCoFPKVPxLqdnYRckQc0MeIg
ganpdZMGJaG+MV7vJGyNpgFRPGgzUXr/+7k1m3z4IjXKfH7IhpgtqSbJQYH7Y/oWZ+UTa83J5alQ
KHTVyYHQ7g5haVBMbks1YvrH3t8uDkUXQJ9m64G3DgGSfo6SQC5neFIgsuAFsaUSs2yNtul0ZhPS
UNXoZa2HksKQqGbSdTm7zdkfvhNvl6+KdsSA5SftKsb8uB/yO9KXd/7P0ax+ZWKoZjYFJH31SCZP
08sHKWQCHfr6cCnJdbHHEm34mwKSEwELPKsa8Q2llNmRcW1pamOSDHtWfktM4CBlS5wosfXbHdAm
1+KdGgOTb8nqey6sm3oAOQOZj2FfpdmklsoDmZCkB0bbaulW1cfJzvYR7ffL+pb65F0MDGwIOOK4
fJBvebrSKvkEqasOyi0bG20GU6nf+zwVfglj7nOEn9OZJykUAOFhiTsZNGnMhNu3xeNR/GpSHH8d
6rimXUQ7X3gqWctt4T7VRuMOXAIWjfa9MtaAAUdd+6nuijLTB4JyFRSg1tWNWuXTMHL3QPew3eh4
4Qr9zgh5/UJUNbTWTZhhtvwrG1L2WIc3c2M7aQ/x6m/GZYLgvnYfeirUKhkqsGAmH/xgoBhpsBTl
pgwEx5AeaTa8ZASvPwe5+FhhZBHYvF188H91gq34aEhokvJ8c0cv8K28fJRkoAWydPq1Rhfb8NdT
iYGs5N927DuLh5dCTZofEDT1VOSltWSF49BxLubSMEycTXySoxcSbo774dbEgUe9uRy5kHczU68K
XAJOPPA5/cnf7q6+bGdCdt0SFuiv+1IwieWU2juuh5QD3jBKzM9hvqQ2HiIHAS5v0utbBGYgQHmm
yM5YAJH60vzMUK0izKvhrGIE4b/XYi1ky2ki7Zmjci0IvNyi2AnuMJZPn8nHknN/uR5TuwTvjyb7
gLVb/1qlylnyx5aQF18ihlNYUZEPZOdFH3k9SKWjgCJCIHnehx2Jd/HPmfKadhTdX9VIDz4a547H
DiGmQ2R8UZMpC2PYeInT0y340VN8VTeBEqQpojfGKs40DhXAjT+3wqzDz3b53Zo8FRR5B2AVmmZP
qihr36/ryJiZxj5tUW+MGDZpzu70OohAN97sxs+YtRwmOTQdmxoix0P/DJ4pQBdwuTwdTXfLA8eI
v/VhTe0wCFVYNvPmqui4TNKTtjZHKJMGHayLo70/zt6blDRrszIMJD8evru6eqdqWjHUItwIIXok
pP4QsO4lPkXpEsoz3yd91Zm+miBPdgP/MDB9uq3nKV5MQJd/nCowMALLJs0SlVa3p9VeU3ADKmZe
UMAWX5u4BsDD4sq4UjmULkfPgSzh7m2SpKQAUrE8Tk73zWjbXrA3jOye2GWieCoOiBMDYEtYnMhN
hiRnQJQdrdLdyGUfHSF8kbCK9x1fimLXtvpCXjz2t0kmR//O2303Roa0vUSrAZilv/USQVdCuqfT
0J7R5WkxKZosUZGskeLrUpBqiTds4/ziNnB48GVpQ9bUKehl99RJUoEL0waCovKlSZo8PNULbwtP
y6cpXmZ9SjUQviWERBydHwKCnIci/I3rUZJJGQQEy9wePwKRvqIERm+2ASIlHiU+i/p6q53KVL2w
YRvvZN7BTEWlXaBx7/wrz/35HPhQ/zAWVLwfLbV/lMdKc8NjFTfm/dmt9z4R0Bln9QIvYLjqSIkL
06u5SnzAmQvBLFalVAhhN0xInOTH2HPDjDteDYINYxpWo190Hr8hMnRVrYB0DuU6Ap7ig5TcdxJ8
U7jXnmizLnACYp+nY4Uu+iWV/9ky6Z7x6vRG3SvyfhqsbnBZU+t0cvvD85inWl8eKvsrNVEgnBPy
CxJ+UNOS8IHPV6nu7qV/06PRDhM9F8KL9jGQg86mXET3dmu9H/4PZmpm12iSqMEBXTm2vgU9a1zo
n57IVzgQyOx3CCHYI4JzSLIYzwkY4VMpZAURm5NJIaQTIQpLqKWcJTZiCJjy7gtA0eilMZ4NERxT
OQR4dUIzWOGIGzooTO698mVfL+PMjxoyJt1DoYpLe8RPAMQ6+SXLcX8YEKa4H0f+ZCPDB5AMVu8N
uQr20vCkhaVEykSbSr+6vALezr0HAjxg3apBT2YkIJsSA+S7kyMBaxGJnQ3ZDs33YJH0wnY7PWB5
EYWdcJvnBR8QIVAJek3fLKXoYd7Ve7hjjt9v7EjhUgurWASsTETy5L3Y0zonjcol2t0YlO8UZrHi
ANduFOVCSsZPQEVNS80mEV36JNCFp0AmyiXVyUuheRnhCqaK1am91/3n1wbiXB26vucqJrtWkKCv
7ZFyEmIeAOhqojPKpp/XiCUsWva4AIwgG3NLCiKzf7QZ0BmGOUlQXv+E+sOmjgzs5xuzl0uBAH7I
/QcjotI3MgEcV4OLm80ihwO7UgoqSKGG29RQQc8pQu4ZYPmodRBOZXQURYoMInt7bTiAVIRypm9L
s2xdNSi6s4Lwxz08zDhQvynVjp9MZ2OYK5nUcWkzUE4Lz6N8Dne4cYF6SUtlY/YLCbwqaqLxmuZb
ogNzQ5TUI5Kp7dUdOdxz7ZWje05O1J034OoJYeIEsOkHKBjPKLewF2AdgjlMQeizVS4WX+tcqZ/E
0Y8Frn4+7mgbnJOaNVTB+VF2LnqFKdkMBh8mHv+91eli047AFpZ654KdmQ0h+TlPuHbm750QlhGg
7O0us6OloV5HWX1Nw67g85pdOzqBcf+RPyVgUrFi3cW08rcSuJbJdws/bYqrApsJPN55aKqIYx3u
J1pLIXXyAUv0EBEYhPoRxP6JpjhvyVfBu/V0SUVHujB+DTVfmwnbRN5IsMZo0N4T/LuSY0xUAlZ8
UQ0jhMyoJSWMcNZfmSMaYFXdcJjS6jsb7LzqH9D6h8GFUPvg6O7OaFmzVRN/9RsAFFZDqndnttSH
1CewANvCOhGqshKvGKPcZWGmTb2qwA3SNCs6tDFkctp3EQ1OWyytovBOMitw9ySWOItWJPKzSVFt
MiYoBqeVTxKx+Cyt+3hFFB7vG6K5HiUJsqWZ03zISIQbLB7kSQEoozP41s/iNiOMMxLU4RmWkfUK
KN/C4EqxqO5vqSghHQJzS700BzMkcyMsIhKOc+Zq5hfbEGcONsE1xUtn0c0JzXpTF//iQUTFdy1l
P/xQB8AUU32nHlXWpa2BZAxGoDzkNFvtCHvQo5tNbt/2obV0oTMnMBAHQKY/eBugVx2yBs9M2Vkg
MbHLDiXttrsUyN1AbRCTnbQvwCqFslYskjiaUqgoWY7teVKnnZ0b3tn02BpxVLX8jtZ8dHiEnUOI
TU6iVopULU2jr8vFcOYUaApHtqKcMGsvX3Azhv/qDg1dL6KO0galU9YC7waCQpJ/N37Z0NlJ8/ju
NV7TBpiCUhrbsjpPFlzoJQc9+DbYdCHvgXkZLCfkbxJTWn8+/Bn25cmBJClT0KBzhxq+rL+xdYBj
IdVbYabNInLCJCfG8KUqfpw5onSgTKnkUKbIkD9gzwdHmKcB8iKe6bKaVzXJ/6p+zwetgzHpeTIR
Q2bFBepz+ym7oOYz1nXVsPTpzsXT8tBxOfUYzEier8HupXNsW2thKQBDpIUtLMApwGuPx3DTdyj5
lznnkojfUXTp90tBDDSp9V9hxIt6BEM7KkRRiwtPn/FNKa2GecGt7AgUowCSj04LQk2xz80o9cbh
YvVtgVe/atRG2Y5H/MHZ1iXEi2fSwna/D9PSf4a68S2CUucNsPCPWsuptw7+jmhjaFYAevP2XtNk
SbMAjMcU8J8c01JKtjz10huSiXqu71eBtx7jMlH6z3uRdBBOG+vr4TJj/huHApzV7iKwMZjfLEDi
WXAEbZDgS1dOY36LlLnl7vt1sU6r0iGmcMO6HNV6EL5I931DQwLj7PnfTkjeupE/7wPXzvi6TG4x
C+qiZ1hYtVGo5HOU2sjEB6jZZhfDCssZBNkHHAyTnlHXRLU3AMffJOOJ6CYbr/BvxR1Pu296lEK0
pX5ysv/ZlQL/cX7Lvefw3TUrKY4fuYOTnrKdvdVz6QMbw5fOZJdXPWSPqLgO92WTg+MF9QWR15yr
AyHOcpwU0wwBqAwJ8NR5zQpOTfhHNQ1EcfrR0OkwXmL/Dq2/zUUvPAFebT6WPHiHy1zrOwZUjjct
yrz/N0B9Rzn8mgCIPBMbhSqCSqc2HABNQD/b7RHRJQRvOEENMNlIwvAytN+DGAJKrGYRrjgLJnat
bUl5/UWiYC/eMtF+VsaN4nbtOXYbfj2dZ5bsa/la7NxfjYeRV0gdPmXABpLpGV74lfqNe9Oh0dCw
qRNnMJ0CybkLruA8mdshuGKog+kZtgDnE2JLB0hZlrrev1Jh86o390B0kaUn/Zm3rVTgKvheT08L
v3OViP9rkiT6Akmix2lv6oJMD5QfmVvQijFIbUNxlEmwZITlE2lVFc07Jj+dtgT7iSLX5FLmlgA4
OulO8RSdslp5hSkWPB0zSlgLyFNYZcs5axYMIKazTCtG6d7tzaYJOK6oDkVhzlBj4l2OLdNQo5z4
9tI2IWO6jQQqRNQUoV3jgC5GACvjlNPjQnpRhI1jEPREud03j+/kYdPsg1c/KBjiwLFlrIJKcA7D
+JAEcB93h4eJ0AwPHmFQbc11y8lBfdu0ixwgokyrzHzj0UFxM0W/7Cs/WIqize/d1SJwcfsWeiFT
DmJPfpsdpkae93Ww+Gtzjq066FYRWLq9swpdPLOjfCqF0fQwQRAk0r4Gt8AZITJmq0wKA96c6qDy
H0GJu1chYcCHzYKepDlQ2ZR0rzJAXJzX/piSRZj+Mxwev18InZ6Ed3iXHLXV0fCEE+YA/NWcBIC6
RzZOnH9wtUI4KMeJpQ6F8bTcl+tku/KXrkSNlolk1SbPnQ7uAozm+RLjJheOawWWxapa8UYEgcLa
PugL/rsqFSRnnqBFuOHYH4ZeKNPPL40pmWVgaTJ6x8xm6pTdbjWLQq6HVx88UOYNN8Rz3z6ltGW0
hGcesGsNVF7HxkElQs/tfpVFycqBklLZR0IVbAPrPHeAh/0PXpRhVdBXQQOzu9BY0LNvtePYypMW
PT4HYBOfOxEIfWCfLRAqxYewRNYS17NDrYugIozUroiRDbSUfJXB4qNkLivo2gXnS3sq5gxOQEhX
oO2H3Xxjdhy+wsM/a/WB07jHKvxttzDtjhd9OaJB9XCaT3oUx9Is5mBWkqTcpuvnj8A6jSvIjnvt
lhWdUed/irUZTNav3BZokoVxDMzYmsHJgwgY5n898HJLM7Ddj762/aa6LKZL3ZUwJ3mySVjK4i6f
jJ2B9b5JqbIsB9qt9XbleHOXZ7Chh143pibpHnqVShUIb1vEfitHJvwg/LtE3UZRSPPtD+tDPg1X
KGlgq9ZySalGfXiKFEAQDOUfarLa5Zaf3YGUYueUQ9p/G9sXTehtzZ2ywOWhKfzoW0UlcnEHgsHQ
Q2JOIC7AgIywwiZ+PexuN+Memju+bqxCPbOkoWssiJ33MZNGArqYTuiz4SZj/A0XY20lnDP/5RgZ
zddOckmwONc/zRk71t66v2mN1DnqXsP3espzNU7mYXE58CIwdTDTNV8FbNpldCz1aihY5xiJ9+Ho
b+KjWTcYUTlmvg+9BhDEvh4U5kdeCV7VAttfCuwXC4jDtM4OP7xpmoS2+9lMr/DIN+AvVUll2xig
qPVvw25nK/1ha0yiPbcdiKoiiteUQdB3ug89Jx86VZXV27tvmMC3INrdeynQz88/yz2yWsVusmMj
AR0c/0bQ2Lm9maWus19xU6fcD8CJHyMhRF+qzFxLGDBt9xINcVLR8R24amNi9Uw4n83hmrpQgaCp
GK27hASHYdA+Kuk3yU6CruQaaq223L84mr3Yn+kIThsTKqPNfW7a0zxoLAzVAtFHhyGDzbchN627
GmZq+oppY9pMszKomvAcGgjw0xndD6Eaw2vh2XGVRupGUqXIuaFyoJHP66G1la+eRVreoyqcEhIB
28kb7IbegCkkY1Hwt/1qXix0pavX3ti7Kc9VkQXXFxuqIF205LiXHrXouXS2tAMPkPoTqMMIGHnN
sLsvhc1Xs19eL3TmKfk5E8p5oqVkGQwxAqbvhB4mJWlO2NuGmbx12EnILnCVVmdorHCXocIKiCbh
W81+NTxOrJs3vvQ2TeAoIvFey3J/xJwwp6F8hJo15YLq33KxGcriupSOPuvYfgYUWOnqjSNTc3zU
/yfl+znmtX0LX4KqxZ+EAAJomXLw6u2JxM8TwxxVYtxqKptERrclgHh+ruPr1a9hFACufBwlsNyL
9El2evV0AyJj0MtXCDIpCCAK4t/XFMDkUtI9FRIlocayTd0iTQXv39otPX2HKwkz3PcSCSSK6GSd
yoKwwn7YLZwAJw86Q/v53HrTK9YWm/yNaio6bWzAm+yNPFvR5ljnNnlvbFMS4844l39DTL3QPZwH
otZIcvD8ikfGqX8EJB7D3B0uJe2ZWBh7vQtXYXsHm2THaiT8E/eC1RCMOC4gYFDbRbughDjSJldD
JYchU2LhJqgipYdiYMzH1c+V7eZfGVTjauUiJj15H2smSZJZj1r4to5s/dFm9o1ISqiV0Ybh0E+n
TXvHUWtCCBXZc6apnYL6rnObDvUuCbv50MXWI5F5wiIBzX4+grnTKFB0KY9gR2JR2yRWntKARi6k
oj/qRTBAvNrkojLKyGYEOCPFWN1ttnbr5750bES7+bTTMf6MRChL6VkSPziVfWESAVNnLGY4nZNU
jbEzpYEs6J8snzRk2x/hH2MIQgU9IaibKWYN6o3AinrgcgB94ghZwk+mAhz5ysIouSq5+WDR1Op4
tiftlRaT6qlQRNLkuIpFaRO1doeJNEjP4o5K4yvLciu/dkH7qVMDQ65Siknw6Ushrp2fdyjNqb2r
5qAjxj4QxNTen+clhZOV7CMm+b7gpbT+1drzv6hMtsj/9BQg/ARH3GpkU6HImfmIy2cLMsTDHtq1
xMs+8nAH29TmqYFWCWG6Fq6Pf8s0OGFA5h2NpfF4+QZ8XIm0lScNbIQJdOiqr3g4L+gmQ70Hrm//
3piR71fzplSSsBmXnLUsRE8IRIgd1M4j1rRxzNf8g2TqKeYLHpe94PsqT3qUV5xaZ2ij2Q0Pc9aR
bxxwZByY16VCg/47zYPVH3+fndSvAFkROmMkabVDq31bfdCQ4Qb6RRSzJUX2xlVmW7eVh/+4cxdS
CPPaWJ9yRHgjBi9VAD46tngJunUxVIWesR/H/c4Q2BOkE0nNfNxzhVjI0VEU9LnyVLeqoJOTUkNR
UmbI2s+2W3pMVM6RmsGWL4LFDFCbmKTojDSVRZnnZVyjsuO17z79+fcyfFxb990vDOM9OEsebdXg
31dmZ0nEs4j5CY/zDrFwQ4AsZ/HIBINcF34IgglqARf4PHSV5ft0K5ysWpi9sgclSeVEQwIYBjPd
7veeDmUACJwPExbKaqzp+hX0gYbl5QZ0lua63+kYpUZSm+qtmglJASbLVPV/otdBa7B9lAmB/NSj
Qk9v85D0y1xCeRWQB/kOEkstQtWcAWrMTh7MaKB8G/GyOX2JraJQfVkR/SZb1jx1eL/cRQ743XRZ
paN+pX2voS6lAcCjq3QK8aM60zeQnblDw5pjOyt9X6zWskVQ/0cfUD1D8ylQv0iBlI7enjbmbajy
SwWTvu7uNJ5f9ndlixJWf96U8SH6ovMi/SLYviOxNXaLyfbOSuZeKhTG+pUL3PDSh1eSLL2LbHL8
uVxOrl22GpmPARcDB647s7qUiA6v2YrUBJ6Rs+JP5P106HwSS1SK5h2biGv1JbRMN6L27O95ZD5n
qeKYuvJkIiox3GS2xy41ylNYL9sO10Wy7AsGTLS4b/IwaNc+QuEYLcpWI0xAf4+ePX5JSDTaU3LR
MGVuxesexvJTwlT1oAb4Z41I8MgQ3PjJAk8v+VzZ6kTeaLUkVb8f2S1QDu8tC5ZWDe3MhXiCWHtr
R52UtB3UOz/4Gyd4uM9vXbzfbI5Ic3n27uCEWuzz3vbMeBbI4LTf/uFHVqbPZnsFDHXuFnXCqakb
DaPq3EzE+diGUWuryWN32BvYW6aCKckj8Y1xG2OYV6yyFXZUbvatvv1Dlq2YzRVqXIIXSLfv4CB9
K+tL//C1qD7kVQVVvQc2rKwoBcYdLkgfoEIp2kezEFTGu03c+SSD2VveHRBwJHB3tfM6uBS7Qsxk
A2nBSP9oePIX+aqPJklI/2Gh3KX6WDP2n+imil9bIvGAv45nWOFzql7APR/vfVa0h2vpLG+d3uch
AByod1aIdVmaf/9aNkcmS+Zvqgf5/U63tPIqZO69TVuo7wYYx9izAeW0eSUzyBJHSFgcYhcewKcY
ASYyngj5qneJXpNOUh31VjoUdNj23NnMkdbqwrOJ/X/AyfHRNZeYNKYaM7v0fsA9/sgjq5CQVvlx
Rxn8WuRr5ovyJWEe8z6F8JQz4IXHB663rMSl9FiRt+CwFCFl9RQPcnuEvQR6yvmwJdZYuovJklE+
Pp7pKdSgnt/Lg1eih7VCp56S1qaY1LuSCHrZJ+n7m2bwaRdWcXg0keCKJMx12p9+eLCRjTTjba5w
7k2AlPrMmxoqdFh0J9i776lef3ULP6XETFhlc8Tlz0whIBF618eszZ31MtQicVXwmXxGsfn8gmzn
QtfdLdk3eXCToKHVUHP4Kad3ANGspL6RJvSxgz74L6lyJSDqVIR7CRJR2Jh6K86hR+gTliCTF3vr
C10w4XzkhAlw5zc4a5J4KqGxRS4/SuRe0R8dSSemCIW09xHeewqOpFUJeW3vNIpuOYdVU5jtuhHw
77biCwEs6Dx7HA9/uV+gTgJezsb1AFdUWOEG70nUo01N4APRviK2gv3Fat7pd+W77P3jl62/fOwz
SVCXqX+8TOrJW6NELAhp3jV/hLC1wggsDq0jYMLJrEu1MXXeXuSEIMRQUjly7m1ggFQsEYU5TVbH
w9qAFZaDQHy8ESf4/7rbB/nQkydqtaeo1tyKXVLKqNG7CeJJ39CJbwuCLm+lQHRlnxK/KiOeVJPY
zj0GTBboTnHd1ABJNoR3kdQBZr8r++tgUD5MpajqyNCLPoVtlIf0cK5CEBqKjcUoC/ZZbEgX+K/m
MqVfqIIlEXW17jrpQhQNibP30HaZm23B2V+rZq15AEn3aTLnilhnTrlcKLwxv4Net7I9O6EhQ9Ve
VWyOvexEAyD/ZsULhFa6lnuZ1XJIrHefigMVpjKjRul9uurnMfsdEMT4k0hBV6yRym2FGVUQMJi/
PMwN6RovSxb0lF+AgB74lTbV88EHvUW3c5EEB7PUEunr0nEVBjwvhG8k/ilm4QPXJ7DsmLfdb+N0
lq/DLJHmbrjUdQhrRrbHhtdl2hk80bz9ORyTsqNae+eBtrOjrZDHzKkBMCJO47Dh3bSjaq9ccJ2O
n+uJLI4Ri7CT57SBRnX2HECU0okKtYMsHOPes/TZMS6U3uLWYynTveAbKcrs8jcdu9LM/UQXu9fD
U6vqYnR8gwBk1P2iPKcgJezWnNfj2pyYnf68q+H5yOKXAcA86zIoRjnVZxMJW+u2xYw+3FEKzV9Y
v6tsV48CJydI2t/DJQ3h1gLwG0JfI6ZNHYCsQLXExE7ip0LkUwPZJlEGbqE+Pjrc4pVcdmxZ0ymD
qIcVuy7blOYLRexGSZwbPKrKMOEv98IJR/0NiAxllRHqZSNJWcRyGJsGo+f0JYQNdTsITSEZ4bRo
1864nPXHONt81Smyb94QReq+P1QeI1HA5ubhP5o4yn15RbS5nZ8q8YUk0UnhUbjMGBqWZA3XS+WY
Az6/GiQN2ohwZAOBd+AXeUePsWcVnTaP4KHqZjA0YnZ+KERtKZXXoXVlPjsoqnOne/k5XkWRPrN/
Jq1ysOvJS8GOWfeZjYpOdGWMAQRtQjvFCULYcWlLGyx+tTzzaw+iebRaRRJ8g8n/Uuet6XVZkFyE
IyyYUkmKcMLDdzleZKzViKKpx4b2PBaGkV0YoBSxS3r4zQuDnpCqKk+1hn6Zr2Hk/CPotoNN/5Va
HFs+zK9p5duxhIlfr24TdBJJJQuptUibC1FoF6UkoMu3pTvmOF3DqIo8REPh4NEIMAr3A+/5uHT/
hdYPaENBi9S6m9ioNA0zWkTW1qzGADQHSyjxPsAVVsYLpYnKm8LRNkzRrMv7fnRfJf3k+KJc3UMj
MFoJZ6RRK/yBM5WPPqiuT6gsWxYnF2eNaF/anXeKSasRXbhr6eGWqm/8o8QTnmyhaFU7AiaP4dCi
BxgidUz1yEgEvqivl1FVUTEigA9mnF/aISUFp2UzdcqBGCYCfDnLZbOtfwNOAy3+i4M+0KpoMXbw
z44+zL7n8PbzxR+HY4coq7A6qO8lcBcrCUIfyh6gFBiXI/SHG4tPMNxYC+nWun5UC8KUP6p4+TmT
wFdMGkBaV/3tbm+IrG+eMxm6wvFpWqcJgY3H0p+rTOKMRTL8X2YzxSdyQ0u9TgAlBGG3pXaW8a0B
Q3R/kKV6Uf4HM2u+l//cPVLonTGj6uDSPrJFiAGgS4N696sq3ZrxWTC1zLtLkQ4ggCetFikcxy7a
wa+lt7HXPHpMQOlJ9qTtxQcRHM3ldmffyFeZNaGWQKxjfkohD+xYLAiU5DjIzyy1q41OwU3eIyDd
xNOajd3JUEKif5uG4hxMeHZRjAapAIIDJ44RozxppBw5gZgImHKbyC23Y4sp/zC49gi4VBLzsghf
wFoahjFaedJGNYor1UkRRcIfde47+91AS36/tRFa7ODfItrotfUcoCZabYGM/5yXymMjk0U0S9Yc
Y7V1MpKGNR1lUCZbh0piRbDtelIOjgvxVEMLEgzQeyolf6w5PdgdLyxY+nJQpxCOsDgEvdQ0rNL0
F2EjGLsR11pvIDE0iCnOtWERVAmukftMZTeqyj/8UNae4bCPEnoSPxFNbMlRyXAIEGmarx1/bG0l
zdI/xbCLd4Wq4yW+WPGAVTS9S+tJd8Gc3p6Tf6GM/qDzQMFYwc+lQ6Cq6G1aSUWRoqeHHhihIM6F
KqEGrdTdWV9TmLZsMVJNxBurGIBCC3xBL/Fi+0zpGkr5pkwisGfgWKc9rIyymjDAdbOUSt/wAaYL
4ddxyrkzw0O2F/4V5opQEUX9Gkbn3VRw4HGpton2ZiGkCRMumEBW4n5E60h6xbpCQcPjWfGMWhvO
N9F7d7hGcDdaJ6oef291lk1E5vKXUeXfF1P9qYD5+gvtiTsoWIg9yEyhgP1hDOm1uCcm/IRuYbF8
R9oiaw8SkBlkaFfn4y5etEwDXQTVs3qhFdkVxfls6SOFZGtBu9j0PzcrZyfZLSx8wvuyb5GsAR1L
9ovkXhhJKgVST/uWjaczFUoOngyr7IhJqZfJYQJOa+wXtee3brveEU7lbZlinhhw7WDNlYpKZj/N
YyZeb6JwtYSm2L/+KRvcZIxaF7TkOXeCvHW/Wmn1SpSATgqYshBeDBoipoLan9Cir98rfaF0HLql
lMGZ4r59O4MfWdqfD/jRcfGsU6bsMD7aTDSQfm0rxYcZFnj4x/08aySgzuEcYQJDMD0W9C7hxLXk
atY37NtHPtI4QlFjXKo+Uav+e5ZuJKsIrK/RttgHLjbfntnRLlPREoAika3BeFrXGJ3+DEoX6lA2
hzsPPppAmfQ/dskHBuoiX+SmAZ0gyyL8LlvmaIbpA5NMpYEGsyWQLGvRIVTF9r37vCV2Px0aGZh8
FqkJB8gd7zNS1dgKVQeZXbz6OBY0uhP8XItj0WoXpkhE053XX+uBFwlfhrKKkEkcnWoLip9tkXWK
YAfzHfcm1RIueLtPRT+25u3UDu1iYGmsv4WNY7wyZ0mbUGpapLN3gdTlxwfggFnr5dFPkPor981p
vjerWLbtLESYlZM5sQWthFckAbJlwsmcBHGzPX8qQRmWCptrNWrqWAN2xNGs6/HHeh0x0mID2EYh
GUFgGnQ2J00jXRoAqXQzC0rIVJk05vu/2cVPwLie3Ulhzqsf7GgplO+bSBO9m236nyHyZOneRT4Q
GICbPeQRYfRT8GjwSWiEkJ6UHI2pFW2OOyy/8jfcJkaQxooMv3bSw3bc3pydk0mfaF1Ol4hEmnKv
TykcxOiJ5+/4sdtWHQn7X0Dkf8G81BNiT7BoKwbAdtPPIFlKTVOXeXlhIADRQ7piq2FVwtLTe5s8
T7QdEIVDSX2N1loa6WkY1HLu1akM/9GKmK0AfA8hmKXeb8RG4SJGkAwja7xLh1UzA2yTgQigNHEi
HYyc5Ai9H0hsz9+tDvX6bEsywTraadH/6QGLH9rLhqM31UQCd6t1m8iNuYSvhzSnHZQ2KiBYN6Ru
nxllkk2GD+6a9k2rO9ACfjFXJ+nVuTAL/Io916Ak/N5o/xd6p8pWljgPZWU4y/38tAiCvlp9TGn8
Aal+eLVNBPlObkeUrGsXPxkVQ4hbIEDvUJCwGqZoJfrrlwuNIixP/u2TfmTQzyDj49WWBOih++Kz
U+cKHpy5w7V2Sye7lMNDZXP/cuzGcfOL57fZTXo5tZKb5eOuVZJI/3fEyrHCRkx2sjzKimAgc95R
N/DLXGfSl56daGCCHeKjPpXp2YH5UcTNB4henXxNVmdLf0sx9usUR6LJa4zfb9oyE+iUs6dUTBqj
VLhCEHYfnGaAGx17TIy41mPtwerYe1WSiC/EA5XCkxWLP6974Uw56AYPHfpigz16WOnVSKD9CyEu
/oOBuMxiUHVd1eb97R5FYCWSxpPs3j2iXcgRy6gpyoTH84AqIBTmYkfhNEehhWflUD/HouGjhsbt
Fvt+T+erQowKWMo1fVJl15UP88XtyzUUa8jYpGPAtYLQwEEHkp/a4L2jRD92noqfvvqoUiIwV98w
CefJkXaMTPiceBvqKw+Sa4eLKb96OXk4XsHSpBAai1v7Y6igTWR/coYV4xBd+g+alEG9mPdj/GKC
PPggn+XXYwU+NlP2d6BLhzjLMOIy2I2uety/sHNF0MDvjoNfPR6uuRMYwzuu/1MK2Or3IQdP8/Im
Iy6Cmf1pDbbc58+qNetYEPRiTqwzMFhgWPvsjKKzMDUO976f3bz7ob6Whqe5viDi3CNpt4Ap5gmv
8c0u3FM7XPr4tD3mIWdhysVvFELooRbVuZqzpdCVUNaT8haNZB3wDhPZuJncOPW95IHRMw+YO5L1
Fy5IRfMNFkTt5X1pSWqBF253o7DHvyo8QnbK5tZ/Qix1d0GHu4y1wVB3xPEgctMVBRyKRFNcHfx+
YP9HMZ56rtE4P/dtGFofUfaeI40ywgzpwpeEMKw17iKCtv7b9tx8XKzAI7ocKdU7jsGlIIGm6XSj
HpHI4/Za7yL0bKir7V81wQpumy66CZ97zua7ggG/rxAvjJ7Gp5UgFzkACJnojPx/3XyYhxQ8HNKk
lF1I4Q5ssl3B6DeCKpMCkDMe1walw70HgoiajWzdisuubKSpNivFY1fRQbfmCcr/jN9ivOGy/6d7
/+51CLbJQVgfKJVywF5jrBR5vz2H7sqsdayVWSxa+eNsSOaB1Igz25LvWxhrF2hZWo5Z00OqfrE9
bO8f7oPkGN8qvbdSH89u5bhZafVS3RHVd+dxu6FTh26lsDGhuPX24Wc5dAU+HCZI5BN2U2j6gWOW
th+DK9a/00HslTqFhPq5/xdCmFlKo1zn0EDZ1MEh/J9VkPCyxVIspbApcdfp+eXeVLIWA83EyqUP
xuA7rCLGBA53kmI6kvfSPXBdiKwPh4Gs4ytjLeGgm2czIotz9D5RPz3FHUzs5+7HzVIdzd6oNmE/
lN5XLMxuLn+b7vLbmnxAoyILxnkLneip7Jb3nVOgjnG2Oo9teoZMBjTHs/+W5jvJfxNVfISXOboN
Uqpnq+ONP2arD+/cOgKUXcxIVbBm42CvlN3UCT5pcE24QUTQWfwbHzQ6lTYFoWcWNHlskQj5YfCx
n7yQwNlJzMK8b7HOizaaH7imqVODK0InUFucabeK/ZdasRdipEixB2crdFZ7PmmLYRtG94sqZc5h
DGurTHAjIB1dfvbgfvw44/oL03nvumraa/BvAkk2sND3aburJGbh9HQMC0rFlgh9DWq7j72iykyF
cDGaaWl9SGNxQbVhDyk2FphH87anD/jjyNJWnYxguj0saJsgnuvcNUOwpyKzB1tlh21USEYIwMJI
VLjqchmYKQjz1okTZj9bMPhIaxXkDgx2GSCAtnxB64npBYzbgv2ufX9+zI7nCFB40pu0ada1VW0d
7t/dRXMTnnbS4h6ALt9ItM64OgeXN4OyZVfSoIX5IthWd+mkYtr9FrxvXwhqs4DAOAFWkS+D6UNS
7EuWM1ObXoWkDIHzI7pe5f6exJKMyQ5XR6MfkL68BmDvBnMuIsdY39mb5Y7GW0jYNzQlaRNRY2FR
dujzwYWdDr1tg54vHowNZc9+AKKWz0CrE9pz1cNweq+GBJvuSZ6yiEr2BAPlE8qkWIUuy62VJJzZ
8k67/kGoQLM4ti3kKHMsaMVS2OvkuLmS5kOKOWJgu5sW//bh0OLvckIkOib72mfNKpvdyWpLtRbZ
YsQ7ALskn9oNfSsJJBo49yJgCPFLAfhl4DvVJ21kuCmZFpgoiI5T8z3LKTvQSSzDG13DwOvqQQrd
baaQtJKP7OhTSif8M/9H43dCUv4Kf/qKmHVKgAWdiCTYJ0jLI9YphLfa+BdCtycGp1TDMXT99tO+
WUJz4NBTuZznlotRBdM8CqdUY6sCf4ebl0nhrYYusCP5eXvJqfpSgqAcKRu3mjGCRZALqI3btOq4
XXK3JIbYpin+EfXB+yk9W/CjC65zVSq8ZvSNSXvkASuuMTGj1hiFYYO9EuiMqDUwLa19w3SqymTk
ZbjWHXx3NikLCMHImiKVi72TK9vKrXOrMP3BJej7EL7cMlIofhwYQ4d8sfRikwzT+1qnMO94lRrx
kkfbNC8td4+/AQx8QTGg4C6rGuijzBd2LEeAjxRAxQlK/KXuJ+aWrx25P+xNUfcnG2p1EE4Mt2QB
/1wEolHqhNol+8On4BPyuZQx+ixbu4uFaF/9g0DAMSCFbVlyrg6dMdbg5ku8ped2+WF5mSMafA+P
LRqwKzMAg4BAQ/8fMyy73SzujeqxIgYgb2H+Fo6dlVTzCEY3NFGY+X7wBxJyVSb1V2t5IdU3K0iG
IOh2dERZtfPY4JRCFPJKBCkrW5NiDZNA3l3rxFyF5h4zUPS7QpbBsCnGTYt/28XQOhG/qqsKi/YU
6muUs/stamvBu47BLzu3aaqcL+OhyyqAGmz9Mb/YJ/B2n64sXMkAIT6dXwbCW3Y6oOZpOVy/syBT
ZV1dCzYOo12vbRrKfTqOmHtiCE5vsls3+50GGGmWD0tR3xSXYOfd+X2lBNxZTmkYDvfravPNbQ0h
0baPDxkjBA0F3nBnIyWmzpvnToO3/+g0aFQ/5hLOVo6UPJ1wGWbRAsESl9yOKaQFC3Ah5Kw9ckmy
bMsdgBrAX5grOcJlh8QKBkFqUVXMzDx+ifgTGfwcrI0Lt1RZo8rbNOGfDBTgawJYlbBSsW/B9nx+
5g/2Pj4UDuh8blwZKt7/5mlqdf9pLK/WE7RBp09ZsQFII/5KMl42bgpm6a5TLLhfuAKBq9Y10kCJ
SpVbKGy/ONLd4EBYTl7fxPSopOjtGKR4mfFPh8EjVbP2tkzda3QuKN0ZKX369SmETfi1AoVVWzKS
MK9N9MZeXK76WChuqE5yl6Ucj3a5DXWHN1zhHrT/sQtdV74qzqkBUQWydjU1Dd8KKRKHlR7kFgtP
A9GE9Puuc33avcF7CCfqYDy6C0Ebct9ONe0wn26aOCBmM9cFTTAsroBYIm3tbCxTIxYNRMs/UXR3
phfOuUEeHXiPmBYUyM8rChhe093ACWMmL5dJNhBpVd1f/ynQK2v6VRqmKq1i07joft196BqOm9N/
IapEpHDTksl7h7Le+wWKWZBRxTzCn4wM6IdEcLCeWNC30rbGuQHj3SO6rPaMSVVNKPT9YNOjnog/
KV4Dcx1TQa+DugjgGKRgoal/4i/W7Nhhg7QK6Ay/nnvH5Vka/qqg8JWD6pAOq6ov09tYn1Q//qFT
IttMSacp6mggfKmLkIaBBhSa1VQxkT+SQPz71c8cnsPSAc1mdUZ5WgGSAtzO7YHJg0hN6vXqwnyy
esZvY14XEPIILmvTzeeRqxEGXFlvFS3QCrA7X3Z/AgtmrkpDr30fI6O6UiMindGRwfD+VjhfQoH4
0e9LDFPcX6WYqqrHYiLZrKKXXce+q1V64ruhhuAMyN7ueg3JWhSB8XQyZOUb7VtfVXdBM+zj/RvQ
jRXIfMrQi99UKmf2OH9llp2nxx1SCZg9Clo4SQce8usD1KY1bk2euQCNmCjTj2qEwLZk6aBytV4o
B25YgY4oVXcTXVEueubE90qevWuNoaUukZr5S5T0JhyRHdLxhBDMU2pH+acV+S5IXjqi9J8KlR3b
bKtCToGYx7AXyNba64fnYACXGtceJrIl5TNZdBueQ6VU7qo/1MlsXpX1SR6BNiuFFbFOd9zKoEBo
gxpVApCFdiLejmkthpGGZP6cG6awCC4RgvEOJ//eCf1mcRyeolGWIep8lfbLYlenjrWJZyRXetd/
pBgmzr6p0RIHiWd8fVsZ/H4tTP0sXOT4YGs79n295l+s+BOXY/7gFASb63ktipfURdIOg5eEX4qu
CrwGRlTYfmcNFiEEOZ9icc3MoPgoKKZZ8HdSBoTyS3SCCqEdix+gYYa2vjXXNFFMTyBeqY4365up
Sz/fvhbeyWj/SyhZsvq4gX0gYofD3DGl/pzvOTssTpNB5Ogexj1XB1KXZFrP9NXyBC2O3jtCQz7k
xTfNX2/sKvvAXiorwVv5uJTjCB4b0uLgQJfsgge5WZuCAMFdTDEa6Qxj83hp9rtZI3oSmkTENNjI
Y4Kcx/40HDYYNAXSU/yCNlhv7tYr6WzjsGZNEZ2xjaPWVPJRdO0W9z59QjEE1b42Feg5D8bqJE14
zwNN2FthrJd1Ozmiy5c3BKHkVQDlfMwB/Z+urcQosHgknpIiNn7hmnPkMglCYEv/3GjM5qGY3mH7
G1Uvj/FV37+kGDnUTf2cZklCOB5CKwk2IpF+hKwpwShLor8cBigKydlCNihkypybUbL8nb/MguC7
8Wrlfeo/YDyuwEYA/SgdXzfu0eI6QfRZ95JdyWW/EK7SEAswAQQ45HQ/+F+7JvM+Yn/qmJ/zCW7l
HLvRjn+TAeH7q8PzZUgHi+a4uKXE2GqYoW3/9HGbrsvy2qbXLtU2mSjBp5op9b1udWQI2Eam3sRi
p0hVl91Az3XYcBq7gwA06xIchTFbccz7SVr/vRtvfMBF8xgQ+1QIdnVmRxL7wcCyHPrkShZWdT0W
nJDMHGX87oaLlRaM49we1FekDlDHG+X59MLg5wRMg2alv8184R5pAXkS6yu51peylxD+bJMhawme
M7qgCzkYQxRLBqm9BGwy2DsVwjSwc5R1FSA0htcyYw/xjUIxJ6NzezGAv4RPE1u8Pa/WOJxfzv8h
xe0rJkT3ilLjY+1kmiiTmwwOs4CS4WUvzTM723pl24LD6EIezJYEkba+1L813pja7SfI+T8f6D3p
5o4/TZ6lcZncik2/HgsXEzF4UQqcZR36X0jIqk+jfuL20svw0ha9I3FA75P1CvjscoqN5LIJXDP7
qVZayZs0xxrlofzO4NtpZiDwyQYjtvaeZvzHrQI64GiE/N8iyhSe7EDwn3c1sFpnxOwf/qHajOex
LC4mSjWw4ZmMsLqoC3TWV621Efd227E5Svg/Hk1yzNNOoosggTyTb+AVkQB5NM92SqP/WezhBPLL
vJ3rfgGrd8lQo52rG4iyoraES59Zieywywx1hhLpooFT9dV69/sp+XkTzVuYhFlvLC4ob41x00wP
CnI0zFMTrD3/r0KK+j8KEFI6EWpHUBpLcn9bGby3W78tjdOoWWycB5GhmVIoWUGuHWTiyb4VMS2Y
VNDyPPz2T5iudTzvAjcJ2EMweL3LolQSQ7f4c7zHhRSm/dHs0+afKYe/Y1aU/aAKh21nRpv71o7R
AiRmDtfCMAjLMwHRa6/wuvmWOaYcEB175vW2Tew12o9ESFO7NZvSSPMl6LKCxCFxLISUCwtXolBj
0mdZmbRILr278MXjP7lS2m3gtTW5BVX+1H+cmkTZ2Ve6rAWJqwtwlUvhjfYOehYN1tw2B7tQIcKI
bCB+7v8RCl5Pb979CHv7TgxAe6BVy7vPfMFIm9C2ELUKSDhgTwvu4vvxA7/ugGb5dJjt3WgoNAJB
xBuRayXckWPfMBO4y0byfzHzKzr2EE/t2zN0SMPoe4wwx1zguGbluS0f/PrTtxtlShwMy799C8Q2
3woPl9iBstdz/6bwkGenJLsxgKYaVBmBWTeAuZ4v4riaUFn6C7abK/8S47qUKizJAp0PT4a64yQZ
YvhGBSb66zBCis2Hl2kI/2+x/FYX+suFCLYUfTYqHCiMVE/ZbyFXKghE6r1DEulkHTCcF0rgOcZQ
NEOwy8LTOio8mO68NB9ilIdfi9PbUXf3rnVsysmhosneN39r+IL6J5u1VSzm7LWBVkKBqGiJMm/6
ofBzd9RnlxHX9bNBetEBL9q6CUHD2iHdi4AdimXvdO7BUOTvekHhfH5Rw+E2Jaz+O86SZwuaNwFj
Ht6MIpTyIvU1njbS6/2Tp+s6q7nJY8usuMYnPxNVNW1taIgND8KJGtpMk9HAkr0hmkjZMLJQdmsm
ZOi2qdjF7xUIpqsU7/kV4UKcpQeOCJF+EWWk2C/PtwYnYIV0sSmKiexj/FJzYfZhg6xVqx2xlD6C
ZFOfI74CbGKSppx93ilyNctCjWQgXWB5Qx5tE/TgIMj91iYXPIsRmdbfdcs17oqoACXmmkBHVuF3
msoStWl01r/PUq3WMN/RwSgv2ktFRQNpLrQs2tPIHIva8mtM3nknqZXlADWrjcN4m1sDxcnKZoTX
Z6aQUIxdFIj5XnR2/yhU8P7VHgIaEcBMoR1K5c07L53Mh+l4VjVTKEmE26M+GmzQ6NMEz+N+3lni
0ckUZie2Lqtfg8u11P2BMxyeC7OdU42ykS9enphvU62ujgi8e1A4Ze1OJ2kwWSqGzVKUk1GC660R
LL26INmRotXBHopC+T/pjJtOq5mIT3cRNu+DUY/iqDzvdJtHBgC8oH5LWe/7MH/gcYIoIo6Ts20U
KQh8NBZPu5zQBawM2dRI9+sCkg3MS3uZ9ymVT899wQG/djaT1KH9rA+h7H/EcD6f/IyjtrdAkV5m
X39knA1+hCzn8VVKZxsipg7E6a09Ln/dU728+TIgssEKRv7Xccu0xWDaCfO+arszVLQ6t0WLDZxg
Rsl+1u+9LG9E5dngKtOwwPzeKqBy/mDzL8umxk/wC2S2m/Nt3MsYo7jurNnuhqRgEqpZRUOFQ6jW
FGaGR5GdtzX1azQMCEyoXr16xP82fYTPV/xBOoSsSBDDHNxpz6ifkZ496IUQ+qyjF2oIaJ76Q1am
BfY/pPcfjdvtr0xQnBkSy+bgRD0Qbc7pXxup97LFnUUm+DCbBiJqIgHAZmTxybs3BkqUAC4alzI4
u31YFfS8TXS6eCYd+oC+4At/kwwlobG2KmmtHgb+qm/7DeTXOAxSmsCtavqP64vOGpnowQnW76+0
tW8Oviw5Ib1fcjxOpMdZVJ8EwljAH03ER07doqV13tIndtEqKWbpVJkiIi6Qe5DpmNUNfEnq5wER
fKFRC3oNgNPO3PO+tTw4qisHiN9phF57re4gZszJ+tlD5LWURhfdAZ0Dese9NipAii35jTXsIiD9
bKKDBtkAXM8BpVGGcU6+/52pliCWPdJZx3PBxCC4pRYWunNzeE38H+L0f68xNLV6w5RMYlyIvGP8
5YkfWk3nJQG7LsjVTzsu5h5XPmkATk9gN3CUcar0WF2zo5VETx4+zEfmCLiQdkGjUAKRK+dzdznL
xcPgPTaz7GcwWDJRVNGclFmZTGFA8tchFwvlMziJYb/C4Dez9Te8FoeleBA3qVu3eMt2mtFY2XXw
yjhQkR+LwMirpF1tTmVvgiXROuB7ioz3deoesn4iOujJnh7kxCA4sfiJ8gD+4XVw9jow+Rkl8oct
zWASHXTQ81RhdZLtaHZs7DPLua5imaQZROcJFfSJtYvohVMhBDcZbQOO/Jtd94hvTFllJ1X/1AZY
nbLptHlBkmHUkzyAXPE2thGa7p/gPmLpW1LWBPfP1OUyM4de+4cE2Q8TacG3VlLIGKC/fMKdOAn8
ulcYub8+M6UeRXxtGGr0uOwRuZPUGy+W/tqz4r4yTgGuXhmPj+6f4FHhMR63Wh2tPVBOIxBrYs8e
IQWn6CUIAzFJx4krX2CWQRwQsHO6oYad4RPMSHKt0npEBF7YJs95ika8c/MEO2gvw/3gqCl6RQzP
YaKSD5T+RnkCxnDv8qq+bmRgcZyhmLEoAqbAxsECb7xBwu62nEH0nmsgt8drpxB6dPZX/pvYeZ1y
BHunwmCUj7L0sDCgRBAUXLnB2d+8kgmw2v276LlU6+FU4LdVvlYjRxxBaHLib+vVpsndmWRfJaVO
Oq1FJhTKAa1XQ9eAVGFHmIxPftr94L94BRlwM13BtGdJJQ3sYo+VTfB6J4rJVHC5J+CahllKw20G
mnjK5xJQgzA7H4GibxM3jft3/chweIv5NUxExD4gijyF599ed0K6/fFUDuPNeDzMRf3nKbeU7BYf
FoZvWzV2jk/XyzMHRGIVfHBFpnZ5587J/j3kVbWR717B7eOpR6h5KbV2h6MglpjleEu4ReI2qo51
EiSt0ItWgpnnap1yfnqcJwK5kpLQYwdzj27jIaGaFF/aUsxeN9UmHQ22y7HbF8EziN4jsbglQk9l
lEfoFL4/QRexLrS/RcK1oFx6eaZniL2ASayNeGMYc+gvWdaz5Xbe+TwBZxqEohfcZHWJixp1J8wk
MhWUxjMaHNfll4K2lrRVXbEnLsbIdstl/vFD5qUSx8sSVhZ0vpPkF8jkD/LMTNYZETP+22c1zrxk
EZmDF815JqkmVn3J0Xnvbo5XT64Sr0k639LKrhFCRJnSB40mJX+66SEt3+7cFkrFtYZutBY79DhN
3gwx23RXkCP3NYB8xMb/FypL5bXZ6n1EdZE0wBDqx8ak5lYHfBLLwoQm58lhXRVh3JVwwXBgsIly
95EZ/U1Mg0bdI3RqHeAa3FrfyWmuew/QXmOMNPTrtzybgP3X+NtcO5JCiOfuMG3ANXKtv4qvmdyC
JsMABtGZZiP/BGtUx0K+gSvnLuLNeKfrDYLtD1MJRuitY2/iAus5dHLOIP+NpCkXB3wBIXvFHehj
7bbIbacZsK+R2O/E1ShvIcAw7in1rgOFwKCgsC8AmMMQwkkMxz4l9M5A1Km/WlDhCwdU5WftbwCz
E6CRu6xSvAbqUEuvB+o2bq5xua81URZNr8vZp79ItZIWsl0WtApxWGIXwWHIvqx7tcmbJwQ2ifw9
zZQXMB+Cpv5Am1Je48giH9wzu/GvoV6gNyRcsmoaOllMIK7lfgbjdBBn3Rc4x0t4R6XWwBIQFKQS
0l8mN4oEqDWX/2Lae/oa34JxPzxT/W8yBtC4Kb/YZYKcDnolVdQOmsG7RausOGK1+/t832Y4e0qy
sOFxjalrJqE+iLn7T2oZLH0HOrt2/ZUDiOuNY04Nrp4qvZHisEAOEfAVcE+atYLM+6rjQDDHOQ4G
qHwXYB9b+8tY4DKyIyQ57hlPKBNydX/zawLk4sACTZQYqRPtcIWo01h6M+KXB6iVQGdpPgF40CTw
mW3J/VMDYr8pnuGa7OxStcP9URDXC3v30OHwT3H2M0+tOEQ2hO6AHegHNPx9jkpsdlqPvO+57NN6
nbW7SvIWYwDdG6RSXFdAPnkkA1X1TXDkpdSvHPiJi3A3TV9e7vVZ9Dth1I7/R6HedXuBPENfTc3S
PH73VRbkhvhmJsQ6JJvYkc5B61L9tDBM5V8A8n73Jm1sMRg+TQSW2zpqpJ6Ve2+st32v60EMbTpQ
F99Sn3QdrQix4V2TTB6zou6R+4SEslY/s+MlYaSTBcWDl42tk4FUnDpnam2MQFXagEpoGenfkuk5
lUCrj0ASZwvXqqXGltFesWpNjPa9M1DjLTrM9L068hSpfWpBsqruuu1Wvt9LKA38dJMQkYuS5/qn
Bi5KJDrWF9VAWVr9jyjn8AHYAwvTFllGoccnc7sxjaA7Y7OFKnP+HKoAxQMzwwYFXfz6gr4KIA4I
+ixguZw60IY/vkrzvCgu5I0T6dIMSQIFOZWPLGvIU/iI5jBbMd0dYBhdl3bHG1BAu5Qiw5DcMs4j
AvBHMp6HOLtbvW6c3firKXvk29hXsi0a3bgM1OG7zcoUvAK7lJzKdVtD8mp1tQy188ZmJ/6pvQ9l
Al3eMYTSFg/cNL4t4AwpA83gLEMiG3Dug4zxa2zDjIEJfzgPk+1S/oUEoCTTivLsdllTUj2Ipujp
qQrOWVHY10WgsTMrjDXux9MdofulSI+HKZUa3nCu22jN507sTX+aohU7U1HrfhJgQheP7JF7EFJt
meSXkrEf5IeJENdFP9fvxTUs4Gms+Y1yJ1J3vGvE5ww65u+IHpPk7Mf7IVPlVR604Q/l+2nw6zgE
xewSghQD8uBq3JbF9ODcp/z+D4/TXytBGwHGPDcPo53VXPt1yDFj50mGetI1cRT4uj17zL51p1LK
jXWAWPe//uSufNzGcsvf9Ohyctnc7R0FS0Zbe3iBSI4YiHhdde6CL0F0t9t5Q19JcBYxOAXUidfh
eDpOSfJeIu0hU2bwITFjhE+EENr0b9D4Yk7mzAGxvle2UPSAnvRx3dGnrpwXmfKfdnYzawKk4Aaq
SYB6CibHrBPOYlU/C/oa8JT8QDnh9NF2xSwozHi9Tn9q/f7H5LU21l3KjKv2THXmrVaLYelq4z1X
gl1sMNquSP2qwF5NEuvDXygYohfnX9Mq1kUk6RdOQXYJIVuP8DrX05t0/I1tz8Thr5RBzKORBd9R
gD3n4EzRaFABklSYpcJA5p5AdapYpIqE2PG2jto70u1hXqdSnayXJH8OD66CVDgphfIk0CntV5nZ
FqKysVGzg4iVc2kOvvPFFZAjcu4w2Ab+qoRi3uUA7JX47nooKCo2EyLGUl73z674gk9NaPN2arJL
UakFN15b1Rn7Jw1bx2CL++wRnfQ0ncXYNpwqXuzOAS6eDNfsAAdF+XXAAfGVb4xrM1OsnSrgKrqs
fy8BANnrMbxYxj3pRzqVI5VKEOqsMd1RSe5J+sYE4O76IKNzbhV40AWA2BAWIVcAvr1rUL9rs3pL
K+jfjOSKUm5BU0j7phEHZPznx2BG084RQDpzBWTIBOsIM5qMBdbVs2hSdb34hY0N4Ke1lxePn2tc
E4L7GNIMw/SelghT4yiaBJAg8nEHGDe6WOl5dM3pD4TIgW26OQ4HvGEaGBnJITtKw5PDILAlGLhy
n94qPCJCoFAvvPCwu0quHIWVfp/FdPd9u/KAvWzXwfiWPHPeE1JMAFFu12WUfF5yjXsCjVZ8amNA
0jzJChbb+ijP79PzaUdj0oAWe9Wjcpe9ZxlNElTOYXNNQ8wrbIs3ZT0/CDgybFmTWTqcKysJdjyc
cqyJ6qIx6y9xFgkHhNE6Msqvhhp4cI+zATUDWqn9BAilPiaQtTm7zz9kYRPgnfBY2dMAU3/LOSiC
Ya9wCO0xnJt1bcUvhDl1/IBwQ1NVY80b9zcrfsL/F6BvB0bj4G/cp9SUAxgCcF3MX2wRhxuX+xnE
GIGRtYyQwO8RzeQ6TBV0SO31DnRHnW1EHNhip7zlbg1X/j+aq83Zxf3VJvZV+Ss/Vu04eiPJCVim
Wist50tHVhGuWDnUiXiDzB66wmyCfqGDyZYk0hcxBxMLE7cHXMePWv+7QyDNSegTTsKcdhC1tAlk
ZWl6b9KTNvBj07rHJi5cAF8GwoLKhWDsmVYQf6suPHHwnrVKkwhY5O6TDZaejdRDH9S41DIWmqEc
vBYUFQo6xYmwLu01FMIe0S41JxFmNJ2/BnyOkdEN435sI/qIavyRZlNo16jXYq7jrHNN8YrzkFt+
yf+N2/ghPwRlSoc1B5yJSjoJ+zczH4HP+1IKC8LwyvQbWTR7gPZpp8w+868i6/IakW+hHtEzr1KL
N4fOCOIhCNn4t7httD9ijB811txiegjK3yc5I5K6YhSI6oZ9gWzF8MMq/Lae2iQ1Vr1nWOZmntDr
MAAg53I6qUdSVoB1whlJiG72M+VLHogMwuzfzd2qRh4sYRCzxCgx8SOCnu00zsuoU+BLohJ33BGL
8BARtYMNC7dBIaVFUifbm2ZRx/shPhQQAwGX5NrB2PCDgLBOFwFP6y3EreESi41GHyVqPLUd+nFq
uts9S2BRGlJLDYQoDocWbuqDoFOYDWQrGSpn/7rxGPA4fSJHCJx8bCPwfz9FmUgG0iJapw8r1+sa
MOCNNDep/ndv/B3NLz+iXDJ7B4ATa34lTAoEOnuRNKMGS/thvq5VAT3EI+CvVRx6xBhIJ+tgJmA5
0dZbNfjwwXRlnYLeZMDLdtZIDcFy4jPZwEVXiUVlSEMIxVTNKeWxMYRwthBmj6A2go27gr+u6bA1
kLugAaEQUgZr4Y0BZUYi4Fb5607kz9WAIDUODgOFzBIrHhO97yt+e0blhLN3v7ZNPJ1UCZMHHT7c
ctpoFmMTZv8kcUbZMFt98Wck4jAn42CArp4C2Tv7ErZGbxghwIKvyB1sY0W0hDAhlfnVCGlo3qET
gP+G4IPi8ehPsuR90714lk1eAEmVt/5ueYsjzi6DK6MaKT1Gt+d6zZMNVcP5OtHmJLxRiXx3ey5J
YwPkWnktPrXIUbMNJVD3Bm5zkRTRE4CJtNfO0/v9PwO0T9Ytook8AQCYy/NbwlX8E0lXL4xGSiln
aLzDrVrn9nwXy3eUk1zjtWNPORHc/4LkecRQaYIZ//mnxC0jmcYo8XnweAPa4k3u2kTXRFFisa1p
T1sduCv8CbOFTEpkYa4XluVTNNrYclxF/iotVziKNwC9hOyA+rnD5oYmenJQsauZVJDNmvvchRa2
M4wnrr4am0+Lam5/8hZF+reSVn7zY30zG9Yb9TabwiGt6RtZYrbKy+zp2JeAaX3zZ26B7nnfeRAj
qTcmxRjX0FEPsiGiBkV4RjKTuUZwV1Xvo1zHzmJItYcWC8d/72D4vBsLyQ8u/HJQ+MA4bYVcDFLq
dl0tBTqOcWKyAwUcv/EtK4Acj7GMT4LK/Nlf5tr9c0ht+o4Byry/nbDuahGfl8Wh7l4zS3NYs8WV
e+6nnxXXoKh76pBilByP6+0ioP0l/KiWHjkyeF0nOeBQ8pPC5oy1PUdbw3Q0fZo5DIP590NSEf2Z
NGK0DbW8cGXwO//SmnjxV5zyb5UGXABrQj5CLIw8DUXho/MSHL22Kn4px0SpksWb/FWrZKZNK6yU
MiVqtPlVx18YbwRrTm5Q8BVFEN3SBv0mnHsRrSOygGuoJy+unlERAOVNteJfmuJ5TS3o/KRfG6jK
mInimInVIPEyFEypDW10HhbZtJLc+CZ6djrbvaS1iLsplDfHr15ckXGN/XK+bcpubhMhpHdZFTQy
1jLGNNM44oUp8p5EDKC5KsbyKsCKDIwhqdK3+OnGOCpSkb39dtEi9yUrD96zdqPg2b60d1EN/o5Y
ysZDX5KFlUlZ2Rxiax59bIuDe9OdCL4QjmYcsZ3GZF6Ha12ipKr2/JWYKiYndcPzUtgslgNZKwOK
q9++TVcV/1TSn1jgDM5Tjo4OngIAPRXRsAeQ9EHaKxj5nFehzf41QYCRtQKypHZDSesS5+3zX+jg
UuOWd76MPpwWfVNIlik9PMwbAPWoKiJC6bzA1f9Y2I0EGhcavoRvyb4nvbz6pAijVRF7VChHF4MB
37Rzm59vhlpl2Ki0N40HuLvH3O4kMPmzLcczbCzOEPz/KYFstTFstPpNbTgbxCzcFlmT40+quK5n
m6KnTbU0hqp5itgeQRPRqYguoyIx6l9LoMcQNPKrdwBlL47vCKfEqJYUCa4nJh6Lri+hT989pInA
nB43+m0tcpt6UxdtIlyUiZux2Z3KCa8yGG2YIezOjJ2IypHk8US27tLPstiUf9lUZc0AjO0MzFQC
2SYSVS9yEQAmYILSHE1oHIGmR7690hdMx7acmCrRXbcSBU5Lmn9od48MOo1vZo4IrNshJJA1YqVw
tf5zucLGxYr23l4icBI4JlXtllUCd08qvIs94oUg+Lb1aPy6o3z+LohW0ZUhS8MMxgedqs7pXv1E
9X+6sohX3xwivR9JLvB7LSVs8GFdR3Hp5MJQWjk9oDicEM6gTXSOcU1eY9v1x4RiFDNjj1GDowpb
Tsq3Uty2B5aITnofbub9mCUk1wZDQhmocvXFWg1yXzAqcBb1lNfg1yacBUleXbimrkcNtOBwXhPH
hKVmwoK1bFf3D+SjSEKcX8B0GHOYFqPFMrGII5soI90PCMnbpNr2+/MjLyVYfBgczzUnse8rw1yp
MLky3aMDNCNh/EFtwTTpfUmj2eBYBggCbjoUAM/X4rJUl6mDVRVtlcaA4X8VSNkrW/4l5monqPv0
FbNYc517sQxoRQ8Zq0Kl/JrZLTmmAm11gNuGmv/5i7dzWD+mnkiDgEIm/vTEdE/vlgFOi9Nona3Y
KjL9IfbjToQTHbeB3jPboyFyxN+tW7mE8M2oYDsQvuvSSysrTWugOBQtCJQ/GhR+p9tOSHh0nR//
bT9MNJgSU7zzy0E7rgpMLI2aMIf4iQL6VKVHPyWtsf+FSbd6u2ch243XUdYukwgRQVN0TNBFGjjx
w5MvARKFzAVD+tNNBEJa2XbToyzSCXmV548yNyS6QxKYtYe2Vue7Jq8+bcyTksvo2/YRLWK6KtMG
68VC4YCbBCgh/N4rZ3rtzTEVYycGvvfvG6ppDIHelPVNg8r9tXaZaZ62hTDH8tHx7/tmOiQes1E8
NcCVCJM/i5hc3Dq/4o/2zspKnc7e2qKFxZDhK/QJtzsDqak7DX65kWcx9WGBghXqGo+j4mP52oym
C45yfoE1WY+uFyYA/ecqYgbf1IaAF9raC9CtUeymm6aivVStFqqnLGnREuZr0cDr9n9gOBjNx/+7
mKKkEBwEOcmFaqPJivpI7yBd7zBP6p+XFzxBCdkNOz2xiX9yHBKFC7t0/goGCrute0hYut+4pLSJ
elWfTPHnK6wSs5k8tdIyHVqA4WEeATYkoga3r8aDDV1aGi65rzLTo3PjZQ2X//6mn4UXY8g9y8q4
IM0DbwMNcX13voGDR4miNAwP1LMiI7NAB3E9IJKm/bm0/WtUNuYCuf91eoTPkXBEJ6whzwzS6xFz
CBbH6N+iV84f5gLRDC2BKBu21NJfLseC1J3dhZW/dm3oYqyX/Z1z1j36CDcisFjYZpvV22X2oaEd
oa33Rw4FbUaFd4MVjTjSi4ysI5JGP864i4syWtjq9Hb6sfLCQjTkMjzRyrg6iD1E4uY03XGHzRjP
K1aQG4SyNVh/ukQUs6nuffS5ZHsgmS15FIElpjJXlpNujDGuMC95UQj1OLBDIYxBZyOyxnqWGp+p
wgWMT+RMVFFpgM3zEP3vC2THK7Ah4Gh6cVAmi2aeESIHBsFP0y5GDdnnan6FxQbjk+/YWOhRZLnF
5+i3tvdUuEoCc9wgw5XuyCyZ0eiWplB0g8HpHOOHj3t13nNrF+oDnLiSOGMkGE2+O+7yNMKLPDC/
QUlEVHqltI1emGgHMpvFlhIyBQAXBLouU/fsvXFVAiIoXwnnAl5vEgTx+jelln04W6KDG/5nmokK
5eusDQ6hkVxgdv26mk+yaClp9D5OQwd/vVNgUMsCo9oqC4utX149TMK0inS7mKejV3ayts+Zrohe
gmTeiDYjk9iKMmD6BRepQR+PAbTdZDjfLvf6WHUHQBwHdFTwpKtbv+GGWJcl8QyUGzWWzsFKxNBH
X2KSTB/NkmdyGtj3Y37w6BcRhjFAPi1So9HqSaW+dHxIMXdIvO0LRgRbLxutg1+6hXwpClDvNPWX
VxRYs9xaHsA7doSBIeuExnOrfQ++DLZLbtvY0PzN5nHQ8stIHPS5d7CZsAHbEF9wZFEi+yQLoyVE
K034P4qVOFmLJjla+MWdr1ZZ8XPXnfd2BPPNx6sDIwVfRzuBmmPTA302vw0FZ+drEfRCZf6Ttb7o
fomVzMHotC3whaEJyET5KpMkW2FRdQ/qJYAFqVNRrMV+5ZD4CyLcKbp/V8KzbrvIa3j2+2+kaLDk
fiiSeuU/4+jclym8wbS1TVOxL7SlxkBtcoun3s7kA+bZyn82NcKlCeJjGLNauPIfydBM5S6I3jv0
Wm2nG0U5/kpZ9EDJFhcno/SMgBVGfAqH+JZEr0mESVaZ00cM7s0r2zFSleS8HhbMyNClXAYgGeb+
8ifJHPjuJjkBPQyumNOHFh/hxpwXRfuUFcovl6/Qg31r3WcAgvl3yzmzRwkfi6y3lRVBY2z4vl7x
3btif2DmrDCffy+XG2M7H/7drUPePQHcVJloYDm9286SvDBF6Md+0N1ZKvgn3DrBl8N/kCoCd/Og
JyGk+nmeyI4uN18F+FxgQR1F+fLOSNRJjy1mAiCFj6RKBLHUohsxp35tUcR0bFYjol6AyWpztkVl
svi1h5kqQHpI+oW3vkkR76uviEw5lVSPqyOhCxFICe3e0ZYHTOTC44Mx5mAar41ysvevIZmEN2P0
Ny0eN+AHXgo3OoIdqpY+vCARzMCj7m+kK9BESK7RQGPF1ATvO/OLsRE8HwQddSlFWTQC6W4AUpaL
nIvRyCzHL7PsHBNmXYP/oYm2a97jtbtXJml0M6aSiBdKpfhIY27MS/6zAXgvPBknrMrknHQqH+23
9XQq1Q38QL+O4WCrWJkICNq3lb8zAj68jV4b7Tr4p09e+BssEzLLyxz/IE0KrJP75R4LeFzXAksX
wvHoR6tfLeUnpUdWHrAW4ouurvdbH2tbONWyaTaSDkL2jhSuvpPZ4bgH8sUfneldb8t75zxZg3AO
scEzmrFuMCxVvnJm+OeKE+K20KmU5ljWlxqSydBGj+e+CtW9n3AIxgIm5dCnrB/3JX2UK1M6JHT3
lHGj2g2Vh0oupHfpTcYsfBqpo2PDvZvbsfkVT2u7gthM4/s0WonuVISnPWzi0W2eVe438YjLry6F
TGIPlUwcKGaOjuC6WOeLoHJd7X8xncsgJxb44IgtPWe6hzSBKLt00Fm5bsvXUY7ja+IYAjBMb2MA
6Y/oV3fUpgBZsvkkciPd9ilQfu2OzFHNXoB6lW2vcwhCRFO7F1knRPo5KPdEylW2lPPDbQx/61TQ
YPXQaDXwOb06ZU/Zz5T/ZxJ8HHnDtDNHqFHvu1gLEqcaHoV/8xfcGr9M3FChCLKb3ftShhp2mRPi
20jveq3LVS8sg8ZvIfQtb9cUMHmYENKiqdLL6bmdj/GfHrRH3q0l4qlqQcJYdxsAX/QdSRrFxlKH
2ffaVRll+N/bAUODwIJwkEPoUEZdsJGlbrseC3n+6MPGgOCg6mlPK326jtWnFj3cc85saRHDFyNm
h0C4P1NxlppWQ2iOfIW+Jk4mDS2O0oY3o60A0E3OzBFEtgPVE1rXXu4LL5i+WlftjlowdaYnI2w/
Gaif8rvAvaVwr5jqVHfgo/SIzR4b4sH4f3YpRzIDztPXGMxqX85CPFFWLKl0PdbEFIqCR5lvVj88
xcMguPvYCsoyJkJkzQeLqbgxbeT2ySPPWJD0LnTZbSqX+vrE59elxHJaYgymgtLNN7i+Y3pIo+BY
plnkf1meFICwsa3oJuqkKOi6qulGGz40XY5GU4Ur0ZfjnrwsbXLSOowOafJifEwswWSJnpKYhL5x
QPT5Ua4I9M2TMIwWo+jpqVneG7XgUDE5+0VrEhGtS8tHr9vsF8dRylh9y+6W3TBrx1lXe3hN4Agh
HdCZoQ9/17EOrNcZsUuPiZVwlPEm0swbikd+1bmc+ZYm6E/JEDZljI5foVcWoCh75p5L35ogAYna
MNIy3KgfFe7gcGvc8yPsJFoGtUNBmt/3Nlh0pkL5yy7UyMYSWKmItcWNp9hptU02XKqtx1RvLSx+
MJ4UZOJExd+qQrGKQHdSbaMfK+RBnNge13gNj6eR2xEwmdAXIyRBtqgZLeyxaFOJ5TLfMbEL3A3L
+K4di3lMHlvc328NLhKDmfEZIXGFgH0e65tsQN3+0kC68gW0rTT57WYsmQgG+WqVm+dT9rsLOlyL
JfBpktf64ko0FkMBuzD1zkx0/bqImj6QHEOLBJm+oWa6f4Ij0cGjKM3TevI2xMre01pf9Q8nP6fO
uVQoFOWU9+KlxoEXPv1f7K/oLvrfiiUaKD7y5bCysI84pZk8v8hNk8r9GmNX3GkPxXkhyAoiXMTb
IfbSeQ6eltDb4rfcovER08o5xRbxsS9NUWTKsrzYQ+Dg6Bv+9G45wJmBGiku2q5I/jsiJ8HBvAp3
n8/dcwQS3l5tcaRHLBkMnfE7eEQYoHCAJVVsRwLgMgTCjI1gRVcteaTQ7SQdg/qTn+Sw3paOqWZW
f4mvEmVSHH4OZYT/duR9B9PMqAx+5M4/bfHlEbaP8oGTa/Uk76C5/7JyW5f59GTL2auqOIL4m6DU
J0151B8oDw61JpuL/xmNhPSUeOFOud9zYKne4mfSRogy0HvPyxz9DSVmuz++a2PKpNRDb2O8xiZK
5+/kuZjB+FAwhWy823VZ7urphPR8FIgSxuVgRFcaL/q6X8I2TQOkafxlc+FfHmHfuOa8g50M5qrd
31GrGggHsZcMLRUEbLhvxoN877GlLJzXd0S4mqOXIfEGFzthC4Jm0nov1lS2RHmLc25dRXF4nlGZ
agHvVBsHmwoQ+3VvkdRAjKJnVZZpx7G8P+VqQvoqssYKmSg+xVy6FkidBVWPdrTnJTYIwItgKBJ+
XV3qdDzbZxU/3dGRvKFSrbCdM4yrKzZ24c/9YbL6882E1l7UJKyasXk/HH73cTacMtOZKBatMCzY
sB2LVp6f/IN4smJ/7jE1y3xKjidGljJTs572rgVvzpKtXUXUVlUcqxBfwIytGv09AOadPVQ2xaz5
HIlXyTmZv29TPwbSPitLdrbMlzH2vnTmP/fY918e8zD82yNzg/zJE9ep5pd4uuUjOBwxZrmMUQ5z
gfXynfpm5RXYanjiFAx2lxtu+blL+VRBtjFSMA+K6eXbNwt4TWU+zJNQrfbzrZgSLx0VK6T+MnY3
rmDG2XchjwPVZgoDaNaEzdn0h+E3SWU5Mzg9/x0XZnmkLu1h6NM+Fg9P4OjOTL7yfqgfIO/NidX/
Lc4Ti2tTST9q+4yC9SI2eCWnx3pnW89G0eu9F7lh6o+zH37zD0aGO/QdLgNHY33VIDbrZG9WWdJT
8TzWy8vLsGq/Qsu3eyitEUys1CmNd4fK0rSfIQYGBjpQj2IV9vC+stm3Lwe06Fy5G28k75q/DGUi
roDyterWW615bnRvulbp0JsYwTswnGA8MKXc7/mOUmUZ78b2kKwkbUvLzpvARUla3yweFpB8xBqK
mBddlJdM1PDB+4/q08sxgUo7v78wkYVqq2G9zeNVVG3SaOgIwN4kNrXCUZ6moNfj3WlFuWrSgC5U
hImcPRYfqv1Xc9ymZxUF3CaSmO0OehIiylgm/OsxutuuNGNeWQUrk9NUiVfYK9Gm8qbi5clgi5e1
8fFBjqzJ2UUyx512+yYkOXTvNdDNwl9pTUcTFpMZRZD4bDAuf4EhadGnjdV5noh9Q0yttS/1z+Gc
jt0Pz1DJWQ3Nws4Xjy2CrQoaV+kwP6GLb/xvANfHfF0zmbDvFwOKLwaNwbC1Y3JIyPqGy5noNpbN
aCYIDsWANoOZvMapjgwV2LTO8WqQ/Ne5wdzakIOgijv9RRgVoIrPkNYyFNDWt3TMuFRONdSm2HOR
zvl9WYEYoSxW1aVY6fFbOFHkZgphwkcWm1Spmm5oLu7M9JxXZCqTLagUy14/sz3UzjLKS+/6B0Xr
6k6UQltzt5SM9JyDiCG+DI6I8AgJ0gM66VZgIOr3UStCIma47uKKY/TO7O4kI80ZuljkkVq2FwfP
zKFSgXwt+7u5avtbQYAdRD7c9HpFOlTD/uq0ORQ4EWgkT58SttwAFM17PLj92eVf4D7dZotAHuyC
6ZeKfnVENsCz1QAzS9WtvwP9TH1UIZ/RbbmRZiNGgVviINHScySStC3oGuAbasCp9JE1p5AsQBgk
8Uu11HfCJF0/rjCpD1Rh6aU2QFRrzgK92D39pc9EREKCY9I18448av6VB++rpdTMBuVWs9cMNeAm
uFu0kX1j75YCGlM2jLajr6hDKC6cDEmiuweFaCk+w9vn+PQBLtdsS+wAmzwdLdZPYbfheDw/L3+S
RyVKNBoyaRYYak/nTctsGpWegfVCjbq/ERyw2VTFGVRzTM9GyBeFmYgVN1xJ3DLvs10LRgxqwo8q
wRcdgOVRbEwXjmGOIxq9H7ZvSXcEJQjvoEsoXXrzmcIj+BUvr0akzQ6nBQIL4Sqb5VP3758/3GS2
DO999CcWOaFmNbbHgl7Hses83QwLZVdunRslKVFd4RVJXe0XImGLMz4vZ03sQ7kYlsz3bo1HNr+C
FYJdHtp99cLbRnuyvh8xsvDCdnvu7O1IJa7S44SpcbYqTMvFhFx9wzK77dILS5rBzKNGRNvn/pfG
1chP+NsTaMrr5TqW4oVPr1vkvC2gAwycPCxTljN//cRicz/DF44O50NcjXYjqfq7s8cwaDYm4eUI
rUIHKi1s0q/9klmnvHEE5Gf3DPUksBv7WomqCI2Oh53yUalCHd2/EKQU6pGhAUNT8/Bt57WrGZXh
Qc4V0QkOBTb2u0FZjj1MMb46lhUGyEYrTqH/ERGIuma+SQ5Ofh3guxgB6ZB8KCHI40lkxTV+O9of
4Ch4d3emC1gPx/7BhY0arL3dUHdSvKEK44gE7p5XJOeDmy8UAZOKWMiCOwV6LecLHHFD+mDEUqJD
o4xhvN3Otl23Y+MEDnx12VGJitdQZ+lerTGih8HNJ9B3veG92LV7J65biTomaTNkryf0aIr1WZrS
z0euqVt3P5gP+bKNTA7/N0lnWxziUvNPHlDJAEQWhtGHGJuKZU7Vos91F1hGaTVXwUgyoFcDO0to
JxTceVMhnPTnzKJJ4PUdT3A8dc26FQ9Yd7QGZ1ZshoWxrwMNEVQYjx5Cklm6623lE4E/jPzGYo9o
aTpLx9CPvrMdxfssINUabsbb3n0+8gmM/5zNozbkKY1nd/ADA+Xxdxsw6nnMv9HBLZa9Mijnn2/s
SFhtgvG1E/z5n3m95HDu1LNXt4w4OXf6fwU0UaOaWLTvSbHIa4MJSIUrluqNVFj3944cNtG4z5XS
YC3eCCFpeaBs5h4p0SFLJAK+0tgNUQHlMaB4wBoN28huhuOWpATjM1BOQ12NTHukY4ge21ONg61/
Obb8W8kwI8XqVfra+0jogtcGxc7IQYX2GfxRAR5NLUCtdwP1vhNmhvW7SPJTSrNywgRYOiJ1Wrbi
QBwqbALVpe8gtbyKAbW1378KSUYoAIWNg+eMDyO1WuKc6Vbe1OLmgWcontKfj1D5m/kbV2YLwXah
ltK/N9PxGsvZKS7UdnyNOlijXc/3MX0gdEak0Wgh679yaJ4vdjiWFWTbInn+lwHB+5BHQ5xqZt+d
3A+bwmuMLqGWkEJ7h6EBnc0ZlyUtlOXgEiCmb/GhYSjSmpsQfAwQmTNRwRIgEKUqL/6uhMxoXCdW
2WmSN6hmh4C8D94qdAVST6gf5kLzYcyxFghTaoMxEJSd/qAZyY7T+3o6huTv8FeKEeRpEp6N9LGB
vycykzfZJD/v8d0z66xs3tHrWlwbbgtlODZRZD5QsKcEwbkRpdQAZMcI2vTjbVsZrS9DiyLMgny9
31ENfBe6BdqIvULHy7WGtwgEE7QwVaXXnaOFvWGpR1A6brMkz0YxpbtoMn6HvMqYpnY0rp1+vrhI
1u2VMNqItumlL7jB+vVboiTICVNhEA8ej2CwCdppwc0/721wNf0975rxaxck6Cy2VB25C5YY0fLa
6LiE6ZbMbaoFTzKb5cI/YK/gFgi9VAx1UYjK3u/yA2MUb/hKmo3q77AxUP4JpP0TUpGC/3vtJP4b
ASZWPlDUpcMqLPlvt8FNVfUUHIK9MhCR7ynk7fLcAhB3oYIm+o81ctrVA3KOE08t+yn+V1+lIh8R
37DnSjTUTcldGf25lCwfPVi7iSQkxdCvvjSVo2nqzmDClG1EUnrsvMU47tr6TCWR0iNpusWpAdjp
g61jPjS3xhIQUOxPxJsqXjq/muiJ4EJh2jvqNAIk/pJkjLAqreXMbAjo+D2OIUNGZnlREE78zD6j
jD4X+mJE2QOw26QsPUDDH8m6PdaYPeelH91h1+9pqwXn9fhfrJQD1Z5pg9baPLzJfLdOOTpN1eRV
Eps0cHku/4Xbv3A/Wx1LA0WqwpLWwUqL9738KhBqHiIJGD+eVrme6S2oA3P6Km0aXIWuQT+3ToQO
oNemIw7I8+qXtJ00oZMrTa+xZlo7OC07Nifs2YvpZVfmKd08ezaNYOFqwdsz7hGjlJ08crgvjoQ6
M4OKfgHcvv0dDW3qaV2yGKWfwwU/lrQGkFkthSWuujOkXfOclP+KR0b1oc1vukq5CFOOI2Va0w+7
WjMVsMmw2EpdhgTCjEfCghlPVxOc8wzGxkTcX/1MT4GDOSgjwUS/gG3oT4nIPilMt00vyTXIsfLH
cNzBXhwsXRgnjIfMYt9mAGN2cxESxxnvKnZAvvihWBruXN6qR6+PAg0mJo4kqcjSbz2pY0sfrV+J
9rLoNdEFgaTqDKNfKxmf/aBjho2NckyobRH/UUdrGUQxq6OqGs6ZVoDRLl9v034OX0rh30hb+h5R
4aU/CVdKGEKdxvSJMenubqcvbBYlpGUrXAHFuoGtpXFDmvKOeUjesyCiUv+THtMsSJn8XFxZ1BuR
Jl9gT7fUA8/E5tA7L6xjK20UEgCVvdWzqGNzQL8k5glRbaCouGpd1ijLZUtWY0CcVdm5HtOBvuGW
E7zUu6hNmBTglkPiifSC+L+4OEFENUKMSY30neZo7IiZS7VyN5pdB8i589v1qgJx6WD6baZ5u4jR
YRJw7HSYYTSfKWuZ2KtRa5TY1rSswUu+z4KRrxsGc0p0ifVuYYw9odrTtstl++7sD2XwLamBl9Vt
+mJ/aggAB7GBBxQ+hguKscvRo79gIA1ezgUNbA7CJRzABN+KMWys7OcrFAiWuHiAAnzvB2+banNI
TTsRLnMM+onAswbEnrDka/ttKdXYsUMAWYqFO3yZKywleV8TUYdCB1FzSW0DaSf7SSOUlaIcT4nb
kBVGLzSr+3zDq+laoP++ZReyqmMO+sUeVTN+UBQulgLURIzsd1Sjamrge3nmMgj8k1JOoObcDacy
tgqSbHxudRvpJEJlcdWsyrPV+rOV3mUv3aWRsbvKZrGI0ejNc5xdjRFmamieqWqcN3RjAsJDw6+p
M4+rKJnmQMXuB331tB0KRTlsWmnKbmtwqX5UPHX0DWoGVUz4EJGLRBJci/gaTQZ8HY6JDiTWrQPv
CCWrSA+s40mW1Jaa/QsLJkbKxzPdCwQtwQM3VX5mxF0sGWRpaAYF+aOXBUQgqu+hbE7bdx67cHgo
UJZlO9ZCop5Dv86aFNQTUg5+xVbF5Dnyikk2ys7/tH6zaEqwoWELWVCCWV0ptjB64pbxd7R3zeFp
0VMeHtdeJIoExjSm9bguMLZRur7rrWOndRXF1R2wkLu50CgKi4ujV4AlJppKgk1CLMBic9XSwwWn
93bkH8qX1dRjv4wpHRTh0MdM23q822zpNymCJHS9HtMdAq+biT8rc3u8QTCSYDmlShw5IeBQHCK4
UMKLx4bwMAkkRAMoYXXivZ7EKxdtaJ0HPxvilsi2I6kZdewQkBZ6NdLY1NwT7KraWKoUcc7o87wO
VMSFPvjrka4l8pKIJcqMWhB02v/gwof5bJcih8uBcUT4CzH5ySh8A35ru81s++7YI4Q2mRbRLDP5
cwYPZGe4hNBoJbvbqxrQ2y5R2dkrykQ6Ef9VRDg4I36+YUAfgaBHOrd3Ixv/cDmm5y5JKd2nmWYc
groMGhTg1nxe3dMvcTjaifvWcobDZy4LYKLTPHDEuibDXnV0jpl+ueHWd09Nd0o1BTqiX+HNE9Pe
GUY4uMX7/GMVNQNXXf4xTjULYSN/WB/ZQLGc2XoE/LauJrelkk6CbMdSXfuiMxasXZiqzeEMR42a
I2YmVqhX8zEKt94myMbQnMTdkyh6GT70nTjH4mVShBXT9vSY6Gxc8CuU6pMXE4wZThCcyYk6uatl
BlbTNArwb2jlRr+libMWRU3JdF2+uuU280HXPBI4OSQe71bnJLuUqUIOO0oaewF7FRFH+UWC1rtE
Kw8fU+hUbAkuyC2LHYcyPlIvDBiVt6mODVycBD7mNRsDoQQ70ClK6PoAfs+Sp25W4B+yafE+oGju
Q3fAhMC3k10qeZB5T6w2/PVCnUZwUb3DlTAGXEtersGBQ5xpsjEg85PBdYCKQwerq697ll45+nRV
B97RsR1PUCXEZ9ZdydjKxE9nvwJo7fuEM14z5L8VZcX/fCsdUm+j+zyM/aRCA8NrIoYpP86rAW9l
tZVWuL+VbgZ2e5Cp917p/fhHO/TM5oWAGK+NVU/ydQVOW+1NmxA9BnvYpr/BgAzETd5myd72x0Sb
5xzBBQw0UPDD9Yik6KFtEBN33GX6Ku19aVPju9s4lDBFfoVaJytLxRZeT0r5MytMgjrPOSZn56zh
jafShO0qE751va1RJHVPrMc51eWIIuDAw1nHWi5vlucBX/ZyvSEPV9vngYRcDckoMMTJkIXGfNWh
uJmg0l5boFu2vUGDWbvMAO4drCza60qXGIQHVz3b5nfxTt0G3Ydn0t5HMPmXpOAfr6JiYj+yGpvv
3uvI6PM7UCwu/y2qYCRYE9RwOWTOU01FKT8H/hGKoA7FKBuZk9tr/Y7K+l9fafJiCmYDis1KT5qo
ZtF5mEW6HBO3L6M6wwUieyLRgjsIm51sGe2sjRRkVlt+xe58vIkj5Pzb3rPR9tdhuSCeuJX1H1ED
t09zx+Dt+78G/nrRtfmZfGa3QMry1OcrZrS2AnGKCzdgnWsCEhEEGRsvM161nyvGppzYDIZSANwU
tPKIxWUd9X5C0Re/QtvQ08Pd0G9FG1p8aVcR4Aa3pNfB6LwZbawLGYf+8ae+q8XYxUqC7HObXBP7
puTZBBfXVqYob49WrHcTempeFx96kbTjW7IvkUbD3thBYJDLZxAux9OmEc1HwbxAiVWMhgGtmawY
gxbh+C8zLRCclY4g/Ony+t2czy+UREKPaj06PQ6eYoOWPXXQeAPMh3j0+t8GujhKrGKuHXxIMktt
QjOq0kx3mbFyFacl2J09j5HqR1CanL4p+ZhVE9fqkoNt6bMemlbFDE9gcmBwkHEjQ0RnG2UEOx1r
fwU6erCTaODb5GHEpMksK5k1mB/Y4LSVYKtphW/ONzw8SACzjaBVN7sTNs1QT+Yjv+r4VhLXbYsY
1JRmX4h/gzuUQL12SsUUiw54/KgKFo4g+RQgsuyNREzkDOv4SxokE6u16xkOKgI+pxcpj6lLnv1Q
4PVvAQfhAHa+mZ8g3ccT7MF1SbwST2wE4HfOzhA70ygGcsn6GL42PEQszV4n8zsjwCSC7SKe5qdB
DMRnCgGKkh3pgpXjhUfDiFgTfUUWAYoK5Pw6m/50A4vkq0Le5RsFEpy2B7ayEnI0OmQ1pPuMO1WG
exNx2oxzRj2lFY50sibxO/bxXGmn/gjMpqjCvFYVQbUcNGQlcg6A5zys5VJxk9wbJ44Okez692m7
eTRKGy1ahJq8o4aNWZnPZ3onzetG4elK8RqDW/F2r+R/0/crOQ9NDhZQwB7R1B1QE8VLirBoP+Rk
kioja3kkwEuE+jGrCtjd6HcvuGRQdrkVXQgcLah7A+YXrnJ0zunUxtpk0T3YYN64NMQgfaM3E/ss
gJaKgjLqZjmxb8kPBLT377KWC6u3CdPEl6lERpwqUR8plA8drfbpE6TVPYsAVpB1NNcRoA5NDXcV
vVb2CUgIMmiUvyENZ5I864GiDaKm561SXUbsmExi9thq5p+a9dC76X1Sp1SdcVf6dzDwU0NMBQzJ
yzhrDn/iRpIDYMDILNRIGmrKpCeHsSSrn1O9aNQrscDeRRFzMQEiIJQOtyfKj2urZWaM0cEqv2cU
bbCQhPq038d9wksXInxEMN9kXxDBGdjsoHBtn+qI7Fphpwj8Cmho+xNKC4TRq1mwlnL4s44wUCwv
DrkyBWW8Z1sVhBjlVd13INpYvfN425r7b764de6DgPVDOtDR4vVSa49YSfjAtiwVXjs0KlPc2h9n
NBMy7EYO8Ok6iMMFg7Lx4cPfDe+EQX3q4AuC2MfJpX+skHv4g9hmMQyEqg6eME54cocFkXPIz0C8
3w+6vNjcUqHSafs4xMzkhi67a5gXgc6GmZQKnFagHzA+/MQCqOYVsfu10DbNcXSL81J7f4uo5IHl
nr2yHZQz9EM0aRj0ifBgfgXLhhKXsMis59b8B9cxKQ0hehSN7B/GPJboP8Ja9S+imXb9UaGTAB53
0+MFe8d/kNxJ7aEEYUWlX5jTsTjrT2KbhwAWdkd+7F7MAFl1uewmqeA9zgGpqSZZowYsrtj77rIG
sgRZOiyaWGopPMrooDCWhjd3zukGhX66sTmQ3NVRHzBzPYkX0rNXopK/yeZskWDoJE4/g2hgNxZc
OzP5UCfvGxwn73YOip95OWbHDAUkYUzZMKsiMnfb7XyKEV68jgS2SxkmF0Z3dOlh33F0v62rZze9
mdyK9nRobg1SwG7ipXoO6IbC9Yd9xnbe4QZLt8ZluVzQGYMuW3EGRFzaZbvknYLlEv8eveQPLpd7
W3vIUR3FcNKdafDsunwehWecZQVpLiPjsG7MZzYSQr3i+SCrhkzCI9jNruvKtgwH/z23pmbixtBV
upnJ27DpWA3dn35aU9r8Lhxfdm2Yy8CwZEOn/f7EFyN9kWVH3NUrRPfyz6iJ3bxHJ89l6jwyaD2I
a7GHxYguLRDjGmf6Stk4attKx0p/3kYymrhZZfl1efCqRFeSlV7HhrkKzeoS8OSAr6QXbpq5ypRT
Ul4i4J2hLSyIy7+FT05cEfUexMYoy/lALwlTZszeSuLxCHw/9FVDhTmDhMjiAQM9XDgGm8tWilgw
ke1EcM9VMtkbEfZVotiitpZGii6PxXFaSY7xff8YvNs2qKbBfsMwZgFOlN+w3ci2Bv4WC6FIR5EO
bKq4V1IAlNcEpDhkvnbyiD2ewKovhdwkefVMLlFh99PCiar7hyEvg2bfQSI9/N4wr0CqUGELe/B/
rig1gNde6PJbCrOw3Q1BfdoikGohbwbX4yedvZhtYrTqBa09BnAkVCKS260LzV2xsdt6TqHobbhi
iTEv7POd99ItVpYPaJGUjCtAwu5VJbyAO2S86fdgZVNn7C8cWnEi2bqoXovSt0t89E9LMgz+pOCr
hgcZazHNl0KX/DE1e9RxKhpb+hkp3l8fHROqMtrIUGTx770cOHMIl9gdhvMjcNtA/o74Ch/Mfpzb
vlo+OvCzJSnZlJxsVL8cGPNhXHYADG9ebE7Z12vA+5wJ3YpC+mnUAGragwlTBpoBSbIAFKzPzDXj
WmiEpMUfHDgVmBNi5+1dQ2v6eHQZcwjCwBuUkQoPPIdP1uC2YgThB+USDWJZJs85+tHtosLUwqNT
1qcqaZ+n4dQu6GFS0toCZq/gZUvWUuup8OUJORYuyZ8axeT8PER5mjDuq7KgVLnKSiH6GakFkUib
uKPQ6JhmCpFm+EcjEvFUWfWb0diE+7ChYARnS3EPXPSA0iCgjdhP4wfFHLBUExfL4QbzjX7TtAM4
tLr8EYKiJAmifDGhjBF86dVlu7Ig8/exZlXTVAI7Qjz5tyCK8pisLbrRA2bfrz6z2e+ny2xo1cBY
QeDmJAUCtI/1Cy2yqJEMgfcgFOuqjer7VnWUF3+5GvDzwMba2l9jgZwxGYOGkrRU36EdahBYqLTU
4jMLAZgvGQeBDKCeuIYsUtOqYT4Yrb6xKod0oQbYoSV5Dp39klxG2HqWZq0ZU01e2Z0jjcFP6Kev
EoRjrmhr8eM3eJVTi2D4dPDmpusIdhHh9HlLLKFwzabbnmzMT8xJSew4aLvFDy/N6+pVZ83AyE1U
YAFl+PleYZQdalFy75oN3WDQmaXExKCD/trcZAr4uuRTg75CtlBtB0mtGZut/0BSTo4PnmMEv7Qi
vkYxk2J55qKUaakbjI0R+bptrN350ndIkLdKZLo59Vly/O+/zaVyh41ahFdYYHtXDiMhn+k38PvD
pf26ZWoKKDDmtKDw1DZXBYJoWnvkZosv0O9ODWT5i0Ye4ZuFF76rKzg8P2LDjScHTbtDn06k+Xtf
Ds2BmzoQct9Uj0aj2kNxx6uKQgMGOcyc/BczhXLNlwZ7KFY04dlXgFOsuioWr2mnaSWOe3y7pUyK
Loxa1RYOVvzz2CMe3c4Co0jQSIRt6BNerpsHcqEVFGoJ2BPsWpu86DTKXdttE1o93onVR2k6mChD
lzrWU/2NyZXwXW46h+/GA+2ebZQqy/izcOVGvCFbycaoLiBrChIbN7qwRBPRB3wMFh0GDJCVHhNF
pZL2y2bB1w6jBPovpy0nSLm3l/bGpY4gu1OgMdYXqGB7muYQWp02yP89Do4NvfW2o9KV0E+wgQ/S
niJ+djo58qhJB37ypMgMsFZ3e8CoMoSkxuMGh2LDnHKKgAIitDM+hYmolU7KY4Ky71SwZfTLgimh
zhKhUXcMytJKQy1mLRIKU/ZL5RExtyMp5dyR0csfdHcO/ea+BZ5XC2ZdTnai8fBGoJ3wFvOHVQ6M
ZtFSMtpw89ubPEfH6dkH9k9/ULs9GUBECAoAmvfyqObwt4pYr59oQdkbA6brkH+Ax7bG5GXT78PE
o1kU52UKbN5/FW6L3qR8kKpLo87k9kt2pn7ioJPKGVrVq9B2L7xzHI1ozF4hLvYFrL6vWaPMoWHb
t+HhP+5uNihtThGr7o/XZhQug3KyAwGdpb8JSVFULV+l1hOD99Z08hdKlFhs1p5XPMBNiVLZZUIE
AB93QlaBquzs1lhTwahsXJUSUjsQBkwfnZpcjJ9jq3+W9nUkOA4edfj7rF2jU729pCHFXVZYgvgH
fv/C9/k8uviUR2ld4d7y6/h5PZWJx7Fn6zY6DGGCH1zfBGI1iyv3OfCA5ZmibmyGZz5VsO4Sf1t3
+9MMhLw8vqNWFw0wM13RLFIwsQXgdgxND/MO4Psdl2H5sqSB2BBfjr2TUPIsGj2F76lnskVWkkZZ
UDK6WwJaxt/3jRbLH+plRARd+jyY7SLVURjh2nCs18ap0xsHUAQy7OEj0Sc9ZbHtBWUZlnEAZIG3
abcuP8VLs0SJA8Lvdij4N78cEdQkzHCmUyQIMuaZ0zID5G1QmgtR+Aek+Qm1aw92VyPyclJPC3Kg
KdVu+t2xfS0XoNefzFaSzDqNh9ouh9sGaGEViLfPMaHgZOiLn0d+1ZHR7lQ+hDe2szITq6RrmBrm
/hKmSOKEQjt1X+6Km4OVTGmm6wVHsxFiP+lBY6V37V8n8MOzpbJVwreoOEqENX3CwMsGhGTGliN/
yGQ98RquP6bkOgmoaW8kS/yl7I84haFqRKJkMLzFMH0a230vU47kXb0sRU4EvXudHsijTdll2JqN
G07cbQXSNR/PPne2awShQblYQia5vZWb0Ts7WugO01yJtxe+t/JGvXGAL/i65YoyAoFyHahxLgaf
7bcpqg5MVba4mr9B0LiyJI5lrWHOLJcBahECxEAKr+OIANNLaYX8J6lNIoAcOBkUAhrhXW0GvFlh
2wS+VP4obxAaeWFnQoLIYRV86attHLIBOMmlMmczUqLOLjR+lpvn3O3mjK93NuHrO1GX6m8P5j9n
E5WFUBkFKUHUZOJado763gx1Td8/xVeGuwPb+V4wCTtba5LY0qcv2Xwe9pU6yfHN7hywRxwy/Dn3
va1QPfUcw/I0eyFW6ZD0UBoIUZ3BPdowDrfFFHUB0K5Tbl+pE+/Bbi+P38ccrnY+8YZ6VuGIgM75
LXl+1+TJCJzP7aalm4L5nMDukfzpgpTQa4OLNUbUbXiS/Mps2wkUtoAgoHKKfIYaUy9M1BoybpBZ
dwPjDVAj4H5/q60jP+ho6KoMAe6uX7XnsM1IMBng4YnvRxuQOWjk2eQmRw00jQGdx8JNLtOv4TYs
7cmDDoH9cu+iX/F4Y3Vipp7HwBPuOS3Pw3nxuKoZWeFGAmMWrsG/mw7vApQkA+cAdSYa15bXCpAv
Q2tgBklHjbgxkPQhF7xf2pWRC9oqgjTh4lhXjcRMtYbBN5H27gczKJyqzKSlwGKECIWSPMd4reRD
auZnJtxL7iriy1uQ9RKzMmJmQd7XO2MwRQvpVvshL6TWT5sEYlkmy40hkIr3kuYVBuakGShNjL3a
IFtV/DWfD3Dd9j1DUQJrfWkLOu2/irFm+aYjfkNT+sItEadsZEl7Fn3rcqr/SGtDuU/1u59I5v4N
bwaG9aw/hNq10iEHsR0zhZIGxQdIEVyyKtEUz8WaqSB1fpiPXP3sj4btr7/pniQznJxwh5HlQY6c
qup0nnCsyg4CYLnh3NRzUv65Fcj44hGo/apq6zy/crMaWwkpoy2BJFRK8bwf9F+fq8OR3DCDgFuV
ZOA41In9PfMXSd8T6zeZ3eUQgtuLMsWJuXmS4T5Bixb+juiTAKMUW7jX8Mhn9k/3JwYmvbGU0giq
Fg4arqCiXsnYdwcpSu5k3VAw6xLUhxKio9a8/3uZGohxgGVo26IX2Cs9M71fGzlDxJbBiJvg2jFh
4J0rpWBjbQWhRJxhr09eoAvG0iljkgavdx5ceg60RwDvonm9zpAPVPadUMPDg3K5R9k7p77tNFiz
rQy2/ZxEiLsKQfaWbMPP5QqzeUqvYcbjI+UAyo11u8yZDXd/gacO/m+IFuCsK2tUoSHVxumqN17C
MZzmLlFNk5Q5jsxud6Oe4m59wSpT4aRInprwUJs05IjsPNFWMWUAxp+7hioO2gOo5Tj/OAUnhC+x
M6nX/bujGuMU3Pmh+iZuBaHZYz40UyGinSEf7lgApyxchFpymFTuJJJYBxDywjLaKV5vidCw7dss
AHD8ikc4hzntQh0RQMkYlIK62zfW+IxqwBMT9DcrNXr2N540AMhv0BK2D/zaAgPmgUACA0DlRCmS
4tUHMaWIqJOpHJ950oGu12P/UeXfwVcVXHE/yvZ/DRGxV0vdy8nEaWgN65iYtK6qs+Pb5b+IqNJ7
cFoZjFcJEep4TdwSZ1Nfe8tJZbPVTX0hGWS+fWD2sVoRB+iQ6Dk0vucZw2hoWvosrUOCPsAVJlii
zEDWxHtiM7IxPLQ+pqImJQOhO+E+i12AyyP0tVzY8k3/4wIztTREspnsymLPakS3z6kCV8o3UClM
tGjQe3JpucJ0FImal9ArWkXb9qBpiE2SKXNcpOApns8i++VYaAuBfCqFOBtZ0R++F1Qmx4yL3zQf
2jwZ4npS0OSE6vnlisrG/FNFbElSy4n1EazNXkyt8fnm1kjj0MsNzstHNYaT/pfdLVZihoQLiaIW
2AWGIFa2joahthjRpzLqK2TfznXGYeHII2QKziPM6SJwlTCGUJi0d2DRA49pzNeeLJYPDJ6T15X4
N1AT8YmdvOvN2e57PFjJ8Q68VeM+OmvNclRcMVhsGgng/qYc0WOUTGxhZ1Sgjdq8QHho7QOcEGsr
0YCvT2WBzijPU0b5e24DxvM13GYNh36BknqgSuPVCfgQEbjipIsgBhN/UyV7AXlTKNarNVpHpPdj
QQ5xOM6qb/3kto+TYNtXZw3iEd3bS+WMfwb0aHy/hDJyipyDCTRV/bz+RK4c7N6a6eOyUPPia7l/
mf7LDnlAAfuiSi1StWyxEzGWXn2riNsxrzwdXZ8tN4T3XpMwCxf96krDJ2gjwW7YepUqddUu+bkm
7uxwjGlBJn7EOy/YNIQQP6kKiUHW3+04ah6sbUIu/6xAYS3w7LCo4yzsMh06bxzi2KBGhXVoC47J
H+XI/7HkqSCrhSbiCAv41BEzPTdSCzxenFXAOa675xnOohOeqZrnXrAvxnbal2Zqv2EYzebI988v
u1lo/AI4L7JJWIfCU4ZyMwU6e3e/p2cXN6wmUWke04QqWt74zA3x4FSCggZWZLbnvUhC1k+bJH7t
tsXKSR1n3EiF2SRpI/37py3H1xI68Vk+Ys6cSrKgXwy5jn/PEHqyg0BqbtfpkrKj6d1tEIongUfn
ThZkTy4Z4P+EOJR4gDxt1/DGn03Af6A3Swuz3pb9euN6LgIyoIKgrdFSVEZuGRmLfNHiP2/rPk3H
OyczHQOmsjBMzugQiz4woKaOw3QVuWtO+8eC9z9KYO2j54hJwUx/xIDRkYjO9b0bMyURWFSX003t
hQAgyPtIXupuG6LBPJc9M8Lh2I/zmG4vXt+V1Sfg+C4f3dbtv6giStwfaX+rIQctVo5S3CYgvUA0
xDc0Hjow7RXSYzx3UwcyiDFq4mFxcKbl+cRJidd+Zhyggm/wYm5cQxjFUQf1sCX7pmHgEzziqFf6
Auth4YL9Fjr+qONT700IeOGOaGUDLeq5dfXmZQXh6vFgdGsdKKMqyWIoER0KefROXmjj3eVvData
2Av9qniETxZqGZsQyqhozAmrhJUkZIwbFS221E0f2r0xhA/05hsfkt6n04vDP+7Bx1dNcnrJTxcu
PwpSr4Y2K5y/OJN3a2ns6ReT3cXGODvjnRkb5Nag4ml3V9SIalzwT6ay/hDY3S7XHwOmrqhesVgW
Niv1Lnjvq8x0q6YkKjycBTyPO5JhAA8n5Nuqo8LPEiCzx2FAa3T69bPRxoi3MI8CJ0EumiFjSMbc
kX8fDtVw6QkZF98ANPCaoYdxtVVfwSuEbKZ8DU1sTg9/zNckIktz+CdEYl1JHykNrB65rvWazJQ3
VOUC29rx+4p+Hr3GTajsql7AtBmtJO1+GO1k5so+sCzCRFkKekAPQLd0hPxa/C0oDLswbnGnevMZ
YAub9qHAa3wATNW6Z15SlMZhmXzdrbY73yWxasNTD0w88z+1q/TeWwXuTEMtG+ZCUBWY8YWcCShj
vdatLn/uQqVnbILBVBbEN1pOblKM/7kopGN7AtT/ikWZx4CJaU5f8h0JtCIDtFiOKZaHhJndtuiH
KXa2l8xNH6DtRloDW2WObp1585AuYa7rB398qAqPI7ulmcWF1b37kycDkDHkOidUZT4ctKO2C/uu
mhhJ50wTWVzVdFeVSlCE7vT1x8Cd1L01+D1V9RSXtvS5s7/oRWUyNw+9s80BbJZdeUuMetZpaWU0
3n3uRmJfHR3cMLdeKOIY1HOb5b3b36wrlad2PgT4lNB9oKUtoZ5bVbLSUwKpF/Mugg7UAdRF2jjR
Nap22TJMD9YDJ7kqs/2WbJepd+ZCyLRzp4XBq46yfE/5mfHJxtNEONekVRymLvobwgmyjZIM0ElX
rVAz9N+v95Meww1eUk5Dl4bxeulyaLD9Ps4+t2Mq1cmDiGGwvioYaO5qvGnQ8oXfhPmrDXLC7KKI
icnGiiVY53VKEBvcUlGi2xxXlytcYqsopacJEsi+Rq35SptjhscTdHUg9/00aKW8ADxT8tgDGMZS
4OmHWz3/BJngYcHwAYNGruk7blKRT/HNaKy9JzQVeXp1FeRA2BxS1zKQ7SjDh7LNO4QYv8bAPIJH
s6d8WNIror7Gaegg8WTvHFV5p5FgLRUJ9jgu0a4G3SJSOTpeGyao+hCHRRCv+1h3DbHUeNjKMSWL
K/CIHTgbKI4ZnqyYeknVfCglcVYDJsALKL+nBRSzHGau3wNXIehhMLUP0AV/9VLf+nwolbRJYgP8
EQqZFMy8dyEAw6coCdgwYjqQw4vjZOLOUednLCFf8gtM0RNMZvrvou/swoTBPrUjJj13o3wuQqPV
GvgmP0qwm+JfwOvgFc40bps4gyOFseZQOAzgEW43+2BEMH1p3ZXNrT/2CxpnCM4Sqdpn3BJXRRJK
PajV0z55X/dnJzXttruIWRTEaT8WMg5cLeJ0Nd/p+lozV3TKi9sfPKuQ6a0JzGPmG3MHOZpG1o1B
t+c/kNtVqXkU/2Xav4QjKWDQLad4mfAUwNwWq1kc9KKaP+kWq/XLZb1RQ+3gJaT4KV0V+Y+bijgl
lWP6cZa0y9rgYFPNlSBsgTIS8go0bzrdicPfxzBm0qMU2TAQgeGB35ZJa5z6dPpgcLMHCsjYFoSy
QEGFHgs3rypCf/FVkrnDTU0sPkiYnsKbuQwjEJN4N9VsgR39iRfhtUp2sxyRaJs+k7I5fBaNNW+J
fXJrRBrL5MC3ZzxJD1/o12okEPr8a6zxs9/R8/GW+nTIdtJqf335pgn3v78EqVexHaDDhhrHndkz
+vNHFrTaj3xQDp4mRr864uuCsnjfJhBR/kmw2evTgDw3sMqmRD8TQ3x09/fRvW8y5RatQX/dg7QO
xyDWHWIc9YqwuFdwP7AKvBbkxwEHVQ0oYGbaRp2PMnuXca6vCaAUPjkAskI8pW9xrrwCF5s4O8S5
tfdniQ3KO1dXcUKha+ILNZ+3eKTv/dlpaYqvhd+hHqVd/wgmnWcvJnVYm2crhCCnp6mIToTdcDQf
6w+tF5gQrWc7o8VNqXBchRfE0gwcJV6hTgFmTCzu44hEs4ICN9ORodMNQhtKKt9Rilfe1HHO8cgj
dD3zGAGjhmUmOBiHl7MvaaOx3brZKtuq1uTSd+w6tiHUXVBPVKrr38sZyJiONVgyHqjKcV7j07tB
fND6mHfSdB7IfdznodBm6k3jGNkMnkbKD2mrTR6k0iMpq+5Y1uvnPZeBrhhBv+m4ZSjoORJ/Rutv
Y53KUI6eHQ8SKnu3whndlXMj3Cxcf9c32HBgHeP/Z3oht3EQPnRWWIcUuGjHDCf+zzsUqOCnycjl
C8gw4pTRCH1W12gkqe2DZM55dlpJiJ3Zycos5N5RtuNy0FxAOyvLIIn5gVKkF6JSKLk/DwpPwX7U
wNt4l3P/5bZ9xRSbOhx8fTSsyZiwhR9bDvKuJQE/F17HXE/MLSWaXy2n1K5VbOAcWQLicmDPa2a4
K+c81ceBUZS3PVsZGQOnA2vJTzjm2uLGINrfL/VVAD15wqZSxHtb71J8n1v40b/R0X+bhNm4G3Ud
TKVp8F4DfaY4KWjur78JHsqhQMps871LTBq9J1wdQHft9EzLhIWUjnuADIvVnduODQk7GJZVr9mC
z+pjtQtnEvd5gz3dSu8Wk761XReBE4i7MG+Kqw9gy9q29EWW1wi94ArqaA0a4cqaUw/scLXPiOnv
GNHWT17Uy/OGYDcVcU5OsVllY3OzghL+7P9K7yyCrAx1ICqHXrU7rHoI65JSMSReeJwblZgqRpsr
rVpI5aOJaiM+OxJe5QlCKol1CLBEvJ1ushDtR3EXB8JCSGK5qCZjMXbUrgV/gACRFe1XD5H+KCPB
60aaS78WjKPChYWjDliTj5kzpu+ru/HNN94uqWkk3NdT8lgz2DEnKtDwev2xPHIG4Op3Pzlwhc1m
8XZ90EM/F/5U5mgMCcFLw38NalUtRtEy6SCNv10gilrs5S6BtNKR0qMQ/MCjLF8R+JtYjxge5bcQ
8ZgqSEWqfeqnDEDiTTKop/kJp8XZrh3DGwB+BDEQRp9rlj6x0faFgkbdXRy0L9i4HzoGLA802pgr
PwphrYrx5WkpTAOT/QLWTRSpt19/P7KmzvUyFIdi8gJrEah9rgGBcUY3shoLFht7MF+GT2Uwb/gw
4NRhB4jRrxQCqjv69G4lc7sLd69zqzUNXvK1uwPt0MZoy5hH4GqLDKU5k7whGRo3brnVzqZW8GEK
ZoS0NV4/9ywOcN8IE0vvwjFFadEHMkqXP8n47vAfMKxJNGXv3sHL6GWRAimcuME8vJdOwtujBTdY
+R3gMCzGX0wiOSu47dfwnPiaRsXJw8GonQ5BeBMYsok3JOwVmHzRfs06AOFDi8tBUs1Di13lFi8v
dPwSiI+8YqOVmSaB+2Pr1J1mDPyWvoFEAfYKalWG0JhSk83UsDHP35dQFzmf9LEzI0P++hRBCaDY
tmUuXBRgJ9Ye8VjG4Z4jsdVqAo9d3FIaZb7bvM5C5zLOzJ5irfVP1X7PaHkrdFMluxwMU/1tazny
ayrikkVX/0djQbBb56G6KcUD7JzbSOXfm/vsDQ7xSGFNec6Of3VeDVajsXGwCDCgPwSh4zycDNzz
7alJeRUGGhyup2TMqn+h9xJkiPKWtA5f3N0YkkDaQTM2R1Gvy3sY4pq22PIbKlV7wrlgTulLAxPO
VcU6mDbLWu06oqnkqhP2QevD0PJDl5/DqHa7UsN9IZM/wKG8h3Ok1xzw0V5qXSJ98Ec6PDmRDTpa
rBWK/JHEao1FBN8M75zZ0wST4dhkXJ2Z5OycckgWYgK9WGiSOHIfvxU/dpVfk8ZoSqrCcL+jXfJ3
LgMRbSS5pPxXjKcR2a5x8qT2VbrI6KYavZHpTJF3Usb5PjsTaZo8fofzMLbRf979HqKgrKxnqYm+
X+oySAEF0bN5MCPcQ7izEj8/AKf19N65HrKRZ9dO6YTwSPqCEkdJamhpkIgoUCpI7CshwK8EEimd
fYJY1o+3nQsmwV2S7/tJba4ZcIScGI9Y7wL5LEqN74yn3JzxiGVAdO9fKIReeIMt5QdUdM9GRsB+
uBSBRzu+H1h3QsT0n07JlPfRc9Wr45JrsRwiDYxpK/tN7WLXt4vxx4Tw2/ZcLx+MUDev39AY7H7a
+/XnEqoSPpK9KmMZ/+0NkdQ24KuafMz+ewqFr+G+FPtbhUFaQiKS++gqZeu9SvBLQZLaCxLB00t6
DRN2xLE6opduo4s5gm7noCRL+I8t4Kua3Bd0QjevYlVRM3sUI6VaVf1WLPFRIGIzzQ0Xumvpc292
4ZuwWixkTyZpKwJEesI4HEdhSKHxfBF4iZxCrmDjRAAJtQaSXh+o/co2fQ4vxe0C9boU7kMBs8SX
BJdtBhUpUzlSmpV7I1h/rm84KLornuLZ/Zc13yH+1wdIylt4fapmoSi9+Edgbegzi9VIwOoOIeii
fkjBRrSVv6wnT+llRY0x+0b6XjQ/UYhtAoumx/luwmk8dd2mIo16MggolzcEG0HridYzbsFthXoC
FgsJ+nFnPQYSkzY9TE7OFBkm36XfDOkM770DdnyQiHCudjbEvL/xIEkMq3QVhFql6o9Zm72DNeqa
dJv3DbsTBrryiJpU7fVdpHSRLmSNOjdPf8kAbJbtX4q09uefKgzDJAOwj2s6s6IKdh7NIDGO5thM
u1sUxo30zWkwfguJUYGG6WQ6S33ucVg2MnDl1coGBPGRFJWTz5CBeNgkrTTv5+WdESMtdAR+yVv2
oXXkz4FO5+uCtO2wcxi0nVyVzyxbshk9NrDrInisRQtFmzqiDxo+eZkcDpX6eyEyfb/Z2Nu5gO9d
kamttyfYKm5yKwbGip/LZsD3U2BXRdF8vI3SREwLDBnb+7Wl++4GxK9xd0moJKFbAPJU2q+ow48X
nL/7dsNm6LMI12o1nVW2FyyuUS1ouew3F0GNS3tF94X9+BsJYYA2/LDIb9NO1Zwjp8mbmFkT+wgx
ySEkGlyruLfaxfcyyW3PiMGtu2oxS2Nl82obKGZUfDYrRLOhTOC3tfq5zMt1EIiW1NOOFpHSUZWU
2n+Qcw/MQWByHj4VkJLnnnCNGgp9fXoMBWjAzy13mqZkbRRDKXWXmHjTOlgb6Z3rEET2sZ3sAE4Y
U08LOMRCKEKACVo2L3h4j08cpM5DVBfeN7avXnOytjGqBTtNQ70UDWPlB6BSnYv2eNAjDT51mKec
gwmqED6hEWhhvqqa3IuPDethb5mleQIhtjRu1HtMHBlAD42XczrCrBf/xmWNqjbN4yvVtFPACsz3
q0C+psu9gr19TNMwUYRsO65k11iME7BR7hprv8k8CEqyWtISmBTsymxmpr8UFa0cdDLnCmV9b2SG
5eIQywYWJijbo1WOd6nlN9x/4mfUWyoPlI50JY2RMoP4I9NrliPFXhL7QDYxWbaKgV35RCMCIXC5
pVBjKTb3GMivaRik2E959pBuCxYnk38X8SCshWaqc9nW5v2+Ocp467xToF2gp95gS/NecZEghIuR
Ipd5BBhKZCuG9Yo7TFXtHVRU1rMPC2EZfznPKjMyHcUfZ0HkKDosit9H25yRCF/3sf1Wq35F+Men
n3HOcIWdKWdwV4ogyio1HClfSaG+ZoaEttbkPkpviUWnHETymldejkFMMQrc2w8TjyhCiO4ZELEa
21JIx4EBRxWOf8y4g/DTHkHdOuDhEzUx+y2Hbc2yNAnAh/EvG7FQwTCuJLXyEaKL14wVZYNsurG/
XLPNMJluR2Z9zR0lChOM3PI3UJnPYbquE17JGvHj7z6lEqQChrsizElanG39FAoEUdO+iMVSYz4S
aJgItqhwdFuSVwgMU3nlBnO0mAMRxoVslcsuj5gVqowggzuXv0RnJqg9dnDjGnqTHv4wNrv3IpPr
xmMrmz9KVm4B4H3OhQwW4t2m1zRpHZl2EWDhCejW2+V6mFBlxvRFu9G0Af45qOTpXFwrhr7ah9dK
l8Tydzh9Hlm7y0Okkh12E2xOjY6sTUZRA5hMiipQQgYUgKjqXD66G/XMIU24nuGuL8k9gSYrtBC2
VeajCifqPUEVO1kRXUCeZc1YP293CXSybBonb8IBilVITPguoRrD0ILqTzXCRxClt/iSadl+Mf/N
jEP8yO9HkHzoMbnbwg9BNvtujuE/bV8J+nZUbMfvktAk2Mu3jMwmErZTBW0TdW4Vi6fgiBytCWCG
gw7Y0SqkdEWd0IBhUMqPcqBETGJCIaDQxnHVpgHRvZtUeYAmsFtbGjvLw3bI+/eeX3bRqeiPPEAT
UcJv8XFL0p3b3XYUQQEQ4myIGhktN7JZmKr4N4/t+3B5z8js7/dEfyxZXO751cbuqhZbUTq7qxhr
Bsw7sKy3+7W1MqDF0AUm0V2pX8K8eMZrLpMmCBBkYrUzPxwVGb0ItCcQAhoSf5Lb6ZgngCqQLAfp
9pFNbUe02wNThm5uMXMpfCuBf9X3quVQ0OewyHGXH+/LERhU2PGnKNJ1DYXt+eUravPVDnPSG0ne
ypHA/zZN9lBnwKQYxwE+uQcm2H7x03pRJYDjOtG+YOSQd+77wzON2s/pNtk7XE0ctMnEn9AE109n
2OS16mPPyfzxcvBUnIRbY3b5VxL6BzB2loJ6RYchS/4G9uLQxecita0YSJjM0cZ3PGXhNJpH0Lir
9fz/+5vrboluCwIXAWAWjDZYa1BdQXaWg5usILhDdmhZG9b205NUmRQEI/pthScstu9DYeCfL4aH
0/oBAwpYg+B/jKbpzv1JR4TDROrgQPUTarOXmvRO6ry7jq7NhSBxrDl3vibG7feMEOgzJjpFYg8K
5TfLVMEbEk+3pFguxu/LHofQRzoTMH1TFMB2iJBtGoPHwr3R+zMa0b6LdiI7o5Mh7HzI3XXeQdmc
ux+S1XtTINMw4bk5ZeRoidXD6q+mh8eBpsjFRr7vmYIQM0mLD6ixnQ1LX6Tjqs8OvA9XzPc4/z+c
ggQxddiF/eCsIKsz+LTZyTZu4oQRvTFbxa4eBH0itlcSs8x4GtCOCKTVzhJEIhSvfNQ60ekMoTYY
TFbJVSRPC+v7KO12ryotv8pFYG/1BI8TSRrc5MnndpSNPjsW01WLdO3GQsAWCGfJ5fzr2umWVEVU
vAQIgIHux2t/3Mwsh7gaf+ScDXYQnO2rjkZUHFN1Fn1X/CDA9zgVu8ek/h1oZy5hDbK9DC89wljD
zzUB25DtbOQPnt86PwgAmacph5SYCJZBWIKIweTamEaxQZmXnyEeUfnVDVMHZgC1ppDNUH6cs14a
P+NK+nGvoSgNza88aGg8mvVTHo8HfiGYSK+qr8oEs1Fgx50iAflg5VNQnTJbJviGewYkn3qe/M89
6gIdejaCPXAlTIPlnaXkRMva1Vt9XSsZ/1b9JRttdEEYit/EJx0a7eyNjrLxwGsiXycCTfkre25U
TM+KBU2mfvYYgBuE+BWxg51cx8o8/hdagE7ENuXkiO+AK/G9sHhjLQwVPNu5XrJ9RBb5kpMW2D6g
/SKldCe5zFFPirC8mAwVujjGLGSW42b9mpe9btGv0KjUc8B2NSPdgmxu2EM8m1YrUOZhRmtUoEus
Tj3+DlV63G9mtjlbzcGE9Wp2Xq4d0rEWWpovj0h5sI7xgfvy5/Yh7cXhhyo+hugESUNZQrBX5B6d
6vSy6iUsciChMGtDfI+IlsKFgEF08ROOwlBWPdvchNuiLfsY1FHgpTgafAUFgLSIkh1PMzX4uIUF
nsB3wPO6jvfmqdwEkw0xZhcB0ftry5GMT9uqBlIh5wAzDRhXoM9gR20mXnSuu5vqNWpYa6lA9MkY
wqZSHuJs4vl+6kLrTqWvs5gzDZkYM/NFl//+9Cg6VmzYs38tV/ZS4y6Z7BjJUiZnK9qTrrNItGz1
/RCJtDZxneltd3Bhq8y0hCuK4stXLPkOBZzZN5rMRWIdAItfEGYrTiBuwl4v8bq7IbsZC7o9i/Wn
0p5PKnl+EzAGeM7X+R1/irmLu4D/IiSUAVMuj9Nm2TNO7rlRgpm42ZjzcNrdFT1RC5rU7cv7TXG9
RrI0PHJxMG6BnsN7Pg7ZMnSCw4lCQx+MKzbCXyNJQ4sQVa2Dltyjfc/2wQC320zH51psRYNumaUH
2jvNrO+uZIppG185GcrDuglSlb3sQJ2iNgy1esclKjT/pVhzYzU/9p241zxMgKOCo03U8NRRySgP
PZox0MdRtnaCpAEbW9E9kub8MjdxQ25sKQXvCseIHPEcyOd9ZshvysWtDHZ5h0d+livAE8B4PdWj
1U2Wp2MSYAkTx6PKBy6HmOC6/b9Ui5Ve0KM9mOZoBIMf3OZgLjfvo3vnzWFDKOx2ZUx3zrHNssns
YMzymaIpRvTDyPcHumb/PXOzKIUscvrYM3ZDQVRmcFNAp2d9oKPJ/cSsjTqxXW2rZzShT8JxXnAP
oHYUtFTv5gsLdevHSBk4Ja90W+x8mFE+K+v3XjNKBWHO9IBWbP5BNPxFr/+Lv9tYamxFEsNAOHeA
ovRK9erOyn/8TxKqE8zGfjDsofZlw0mUERzdinA/eA0/G2sVPrjAoFpF19ieBg9PvgP8FSL5fwx4
VD2poea5fmV3hm6Vm74x08gnHNXZys8ncxctD06F6XB+utbG8WvGevg1aphmk02sxL1H5XkuLTZj
NoKU2C3RMknCNIdgP22pk7NiQO99EGgwb1KHOdNn45jgkDfwciWk3XUKAlUJs81t5VBPHBH2Qc9b
58yfSiZv8VU7U8J3SIKboJsczITh7B2j0juedaGX3h/DQtGUqXWZaeE1yVmUnXJVc4kpj5TfvCa8
k2FIWeFK0elIAADpe0Ez8FsZPAwIHEMPOMEgCxau2Pjayq3ijWqyks9bLFdufRz4zN3vl2CM/bNF
lieeVR4IsmID/0k74gXALxo92WXCUFaYG2IdG501GD1f9V2zfWOTcyBLy81QsCE2WMEXRysIjoMU
Imwv8YZ3FZMg7+yJIvG4AQsTKluir0Tv69i+noB14znCs7YwRcMlpVE7QL3d3fkmhnH42MI90AP7
5jkD0oWtXnM3nebWHxgZ6dQVw1kyFuqm1cnOp31VFk9Xdx4vBG6Pe+I7qn2vHaC4uyqMPQDoOKPE
YqLWnvsVexoU9UCDOsdOVJMCTV4qVpnSCZw+SgF7Jh9A3WuhGrKrdKrnHcyQx8bklsYFFciIHoiQ
ys/X1K+e6VXjqNhk2ZNIwv4DGBZgxeu54r2zSPSS4JOwWfV4JfpZyX9nTUwPoawmcWEhe+W3igH9
FZFHNz8LJibSNMaCLhnweSq7ad76QecM5DH3EutHYKdzav0CIR+byg+5XOdsxrYTPkMExdZNggUz
8qFvCUXx49jmExSUQy/+Xr+sAqWU/zrousOx52JRYL3GTU/JiDFU1RqayEXancNp6kcr4qjkShH7
VRHw/iBwEm4/TCiVH+oc+iYza3e7gVGgiv0ygj7JYAEEbZ8dV5pwrdqvzZJwG1sDKMawnG6vFg0h
EEeC41jUn+8UtNB9eIYtosWnxoGy/4WIcIJ2k9uehEBfzXDC0M2SaoV+kGB75+QzSgIk9EzmiDJF
qsNQaulb0sjzsd/wAK8gJGi/Yh79nVLpLIxcFa4OCvMTUAdbAWhjfDALV2tnhP6ffiMhtulyNP8y
74r3IOWm0xeaAwYkrq1XYe4p+r+KSFquD6emj6GdgmlKJjOTZ0kBCHW2EEJxaVkxlop5pPL2iOtR
kjaqkavjZq9B1v/0zcM3xCoBKZsMPdGFVxYljqlD4jQjewJyEbWqwdgMVrd9SNhqoNn5lqSm1OZq
BO2TU73R7r6l+31WnWTzNk4rb+Gcs+CcYdzys63zscA1iEaD7t0EWrJHSQdLw9Pw+Mr79U4OiB8m
xGBFOo/6a9E+sKnyGbJujHFznbKnmPLcUMZCCY2uSns34/L6N1vFjMrRDd3xkB/z29mZPHdw5hxO
0mOFJjtQ158WNmeZS6sJI/2HT+kwaFwiOHe/iXt6BTYNYmoXMg0rtzZom4yh2NvsQ0cZvYl8YWwt
GesfUiU1HTgUi1KyKKcPi0bRKKHJE1SFEsu1G4PgKxExXCM6cam5fJDcjvrfIaZC8/ORF4T+7l3b
vgArlNyTKi0ai77sTekswE/UEN8gLcGA7aEjZ40G+opgyX8U/T3Ygz5BUkadWHIk6aKe7CxU7XMT
3ohd9jt9EvOCIfczEGPYhCGOVwHYhepo/f5XYQzQf69+yHE3SPqlnj3Abrsqvfr/T+3Uh77rkhNt
p2eSGv3B+OzHn7PiwRg9V80aNjQpR9CVI3cciD1pQDqBokvSLF0L+fm5GrI1HMEh0sOPiKCGABBp
jpcDYYO2IgbR4lG405z8ggJ1/43y2G33jw2GDBvm7oOZ6JpHSyxKO2EuH6FAd64CkcvgtwwYBTS9
/jzMcoTMeJmjZwmLHqF/bxepcPf3msgKCD1HzoBHgNG6mPKnzvhrnpYVLIfg4fw7KXYrg9rUzMii
wJHmIsYcSasi913DSzfPYRVw5YpehGNHIbzZHBLRSdhZeR1Hn3LiWmnv1Dg9SC4fj6zaVu6BchAp
trgzTIn0RQdpxfRS5MpOK36Vi/+8EKVIJo7ge60DwcZa8MmcD/qm55LOfkas1cTbk22y3HzqJtMF
G8LA/wnd3SD8IbJDimMokxrcoAA0Dwx3xWkaJHhx+/NA4dosAwcicmh1ljRAXDhgKGjaMV/XCXTm
60bF1UfJXwVG4sAfXNUWzRK5a3CNnEH1OxVQs1mEZc9alVKVmfkQ+ArnWTiW8cb4Jj3h4eBBO6t8
HYiMzWK6LyNkwPDzc0RyePVEUMe+H/ENQHa/fGRijk8mZUcBzT9J2L+4ncjmBMi3ZEyJAZL0+8zw
X1SafO+ci4NDPUxKP74HFCTf0sXawXFgLO6EHE25OG6170CPVSw+PgADhj5OitRcKmn71BdvF7pw
03UoweFIY5fVa5s5vmW/ZyGgc6DIu347CQwR5YFwbkVdXXQAvKLgeyepB2xO2hizEnr8gqzPTdDq
D/UjpuIGVzg3udOV401rslb6nSpBthZWyzBSjN3lX9P+JaEqEdlYZ8K2RLmGEI3kqPWCqbAeNXpC
seZoeo2En0h8NjiLCOzJ6B084P8Gzn4WxBPP7iEI1IrrvI6lkBGRLNtjzbELZDdy4ZYoZIV6CSQP
/vu5MnP8uSSqTpLF+ig462h/K2nmgn/19XqbOKy9XJ7pmezgZN/o/MPNgNLogW01jcxCCM6BjN3d
5ECtBfVqFyJJ0Bb+IFn4XL4+4rUoABXAThVhF5WMQYIT/Zw9Gw2HcWHOCWqvZgCM0roVNI/2hZl2
0IVLceVU+qMtaHezrzuesrE2iMg8XD6MpvPOeQDcUrQbE70kdCexw86nhCEOisUh7F6XnPPIDEHj
MmLzBlI2hHujOYVLDSf8f6/3y7U3f9g9sdZon+YG5RqctARR+OlVu5QEKHMo7GOWSKOUMFkNJW+0
8UFwcSoBvfis6Er4uu+J7SgQQVKhmAFsOmhuzlX7kgOSsjHAoYMWjR9eJOLksJX92JAVQYr53I2R
+Spr0WvTTAdxsBLx7CAnsyLvxQh0hV2+b2YCiSiYkyqNvsr0ut8OUt69OTBaJFRT6UXn1/qEnWg4
4n9rPm05HMKJz/wCbIaUQ91bURezKUDN0xo48RCCg4BwsNhYbeUV/MEYqswrQW4+ErdWoU2ePF71
G2vj5OI3Pl2CA5i3UyCi5xdQt+XTH5p908yvtTMhB2Cr/JSvPlqjfbcNRDHApmP0wVUfq6KqQGdS
HR7yPQvJ26Z5yAy+vK/r/eFBM03irdqwCtW5kC6Y+BjR01RHrluSJk2WjxFvQqc3keHfbXLCxPtb
IalAQbTPyahedtakHar85ABwpzNOb/B01MAy8L9VQYIEDGtMj1145XEiVMM2En2tSWMtVM+sTZgq
dfJbJzx+7iwR08Y72z7/+P2JtT1glWPqzF50dk/U4JtKb+CX7txncdQxV6sUfDen23/4JYucsxkA
z7Y6SdGnQQ5XKayd5igiWGcIQy6uGSPXIGufGLPBa2DRkBLT+5IJP2f/Nup1QBd+XUO9fNeaq3/s
pL0mT6R8Ce5vxlAOLYxI7Ut/RE+G/QChDO11BxwgomBQIYBT93wfLaJvOsevc0yA7Uoyb2SylWRc
Zo3Ja2ess42LuW+FIsNrA6t5fNtbSsCJSVuLOuJXlBDQqNA70nZ8i1w/LxAq+KAXA+xKue4EMXWt
viCPmMNwRXsg3EECoBxsfZrVqHt9870ci1w40qphl/FR5pLY8B8chW7OjZxicVg5uTR/YQek1Ndg
UYdBRb9uYBXXEfAekWD4e5rBzroLU2b2vXwlhxX0ImKcyIw3XR685edfbZW1fnipNBZ198RsFHke
/b21PBVkTBW5hFF/UM37ln6Xx1jaq3OOY+IrJ8HFk/6OpUJtRNa7FQeosG5zqNFLa8jWqQTZWymG
Wvcs24PcQEpeoBGX0XzWYUZK09ljZFCBkdvzWCEFWSi8O6SEPFgy9Ji0D+wHt+gLaOHF+Snvbq0T
W1vwZSPSIKjHd7BTZHRA4It02m5D4UMlNyuP3bAgtSrsyQ+vX/Z7PGWEn93ibi86iXzWyHWX4pS8
3K70rpq1lM4e0SXPdQCN0NgXrcFm4wLF/sIeJtvTZzjl1NAulWYZ2nyU45roxrdiTloc8mp+wdeu
HS9ZRjRqwVlGxN8C9Z91rFQRZKCHISkRmEQWSVTZwTXKh4xdTuSKF53+Y4YlTNMk0nREcJxOc6+i
VkY55vp5dADR+WyMCKaRYpSFwNCf60WhGTTDelAt4bzeOJ3LybUBotkXsv4ReSLqjQ00RIxavKFo
2hdjFYju3/jbSpx/hglrU8dt/zCE91Whomrxh8F1GZyyjZondAnAZl+DOfs5CH1pJ/iCa78IPAqN
0yOipn/Wn/GZR6aLAle4huB+gFlPkUj09ov/niytIrziw4EOQHjz+f199nta/vP/tnHUpedk9EPr
ipqWeM4FuBMCjv0q1yg3KFnleCuLoH2xXP7butnrCIyEE0OvEn8/QLDLCZxsBnedRH/0eMqAX1dP
hKDWGdD+Jo2R09y9BokgBbWgQsM17WoLLNq1fOF5GCsXZkLlrAk3ErYeC23jX8aBXsvZ0y2YQIJQ
rXC0HR9Xi0RTHQJrLFTig3neJ+vLLdROqm+Z+K6blFnWuYHJxvp+Ke/RQDRorRFhkl3xes0wunO1
SGZOdi81qceCGEGLMdHnPx2Fwt//vuRiBL75lPC9gLRaEKnHmran9y0afZ1ro3KswcTMgsWr+NIz
02J+AAfWB5FRPqYc7qJlzkOAh53PcCmhGzfFD3Y27BeROhX88gZvv2PsvJCn+5qHThOV2U7Mu4rw
RedWeVTjeAUT7tVrZnKZ4YuZhTUO+6dwNByoeuPEr7bYh3BL2IPMJ7sxQAE4RcDw2SdH1nFmkYgt
3vd4eSgwEjk6NZhq4XTKy8l/lNnOGN7h720tNJu7bQqmqA3grQ4UciOBg36vD/NABLqwmJQK3QUT
WiUqvRNSlyJz/roBobP9scfTqO2wHyjxhlBBv+unqABqgWxPAnNV4dBZXqDl5yxMKWGiKLdnlmhq
pdC0ImZ/ZSBicHgNjUtp4rbp8sp7fQcF0erYgxDGXZCRUQNIMe4A7Y/FDzsXupU0d1jkeErNHzaH
v+h6pHRyFAKA2CqNcU1mreUvmsN4O3J/Nmg18bCN0IPrTDKSt9aSsgjDRj6t73JNOMcRoyoq1hlc
Tyw09zm/8RLc2iloEkWIQNGNhMga5bRF9M6+EtWM+fH2kdnP9dOAGROTkKxeYgP/Edt2eGUSv/a6
V89Zn+M1DCeQurUu+Tka4XhyNxCutma2l0IJbwtpyqPZd/hUIPE+nGIieZyt5MYD+Br3zQX4pWX+
2+hgInWMLHZXElu8FANsLUlTwJERicpOPQ1boQN9qzg/v/akLcPawC5bg/Q56OFeizdDWfHNtW2m
MV2Z/GJaLxivptmbbtNNfYmuJikWqgCgtG9qIZcqp1DdO71uQGn4Q/jJWDrmzgTnx4zJyr9Vzaef
GxifauLvRXJo0jTqkUmbSiWtWiBzQOf640DYbZZ9m5pBCxPeyjyHOAPFxSu0x1B7vlv2Rdg24eYx
Bw8AV/vnqeNgkNI1SiztE+e1qtq/FfW51DIxpqZ6IkXjEUAvtv3aK76WQxY3u2zIbzKX/CZztu75
3Sp6ekhQDFF67J7aOF6B9/tkS2TUT/YLTYhGmkLkXS3aYCuWJqFYlDBxQHEyd1zxCjhwGAdc7Tk0
Wad5khbyNDJElFc5EJkSWKdW8eFJ2ez6SjYnv9HCPMi8oZ5ieArt6xPv/uf3lKC5TIvB0kqNiRCK
Ud1G3Nplh22u8uSMQTi2kU2asT7gGPf+YeekOtQsUgQNGvxzF4rpnIv1OPA1jGi0h9qKNyS1eOt+
g/np5wWAg5spaUkTaVF5buHQGo6KP1fvF7Jv96emotfauAseaXxd7mw9tj8B2Sefska0UalOkuRS
B9tDJHC9XopUTW1cZzTI8RFFvZIUjTADakDWyZ1nc7RbyTdGNV5R9csE26iMZd6N/6GV5VjLFH73
/lcYdYI7pJLfGAcpG4M1RSFsAjRBSvMjZSCpxyQelewi/fQdk37RYY+MzAMRloqOfuzsxqXJtZ2N
LCpw3ucgTFn7WPwSroYByRB6Uhz7aPRVOls7uJ9daCG2+4Lg0aj3NIG/OH3wlGIGWEQzVSSlOsdT
WJh4ibuMhvXl3AwFr60/j71dth2iyQIp7SBuncMxGG+blxlzt5vV5Ce62cUmYKnjDTG8J22E9ITe
m6FIHtDguMpPXxLsjPGTgZQInLxivUa567UK1b0C/9njgJ6qjX5yHqc2U+gM61AExs7UvhsFsH7U
FQLN7Jnxmd8E94dBlnAvVvCsG8L5IgLJY9845sO/BH04604HlIBAbNHjQMTDDzLmBqv/A5ogOLP0
y/GxMiXqyS3s1xE8O5kG943CqYuZYXYkoeG7hvc7NfHp0QZcmRZMwYCIttGPqVGhtmdqG+v2EYqp
53zjmqwB2si9/twWbDZBDuiZmpPFezs/QMvbPefz08h+xqMlbh6qnKe3mXUKlClIAfDsTpG5ODS4
OdAfBXQJHFSrf5q2m4tFIOguH9hMQ/kZNc0UXqik6pK/E46uBuCjhdQrdsaJgcIHsqD55Fwv+PCD
6QcdcIlH7yHTBIkVUoVMSmzE7uTYzYBmlrl51rQNBXD89bxfHoG7S0LfzUz/bwqh5d4uc4W42KIn
NQVFjIKzbp1dF35LbSV/1K3vKAIj4QrNwoY6jir07QSBp0juZW7IU8W42mAz3n/PNC9Sdh+cvEIW
9WB0hoTIiOudeLuHivtdHWteJ0/NpiqJ3Ti1jsLOnO6AhGy3EUWS7uUmNNj8qf+AuVJ2ZvdjK1nu
NOuj0L2jnZYezrOFraeK4BwQDcjMsMAZIS4DTgXNmGszOPgzQKnwyHrTGSQvTzLo8pe9mFPBCIyk
Xs6doR9OJdBAcSp/SImgOLA5LOFhGihLk9z7g1wpDZor6sGey9aKipSImCnWrb1ZVtapqnS3WmtP
XKcIJaUJHHo1oXCFTKbAQaXHqp5rHDIGjJc2C+7aNzXHmGon1eqWGNWBSCMYPAdAJVzGF5/bg0Dx
/ChwVGek2U8rAFSlIsMyNHCyjevNq4PO2vpClbw/rlfv2EDMNCjCKrB84hsO20Q0aj3cOcQAk0Bv
82qMVungzkk4P0hnlUm3KlwHSz6ndxPvrw23T8+pQ4EMraiOgVrFN2PxipK2ZmCs5jBQ3Pgnugvk
4rITWMvNQYTzm8cqW4f+pRfoUbCpAsorOt7ocEY34kf9jpO7qTZQjS5zPQUH0IE3lMl3X05AANZM
kfEUhbx9TR8HjGbxcSsbJzj9UNmljTPWQ/00LihbGBGENc00lbD8MMbo3UYLdNRELkLwEIYQ9yjT
sh64wFGf06NeSs/1dk0zZDMFVaCb1abu4dNi3WNEVypVUSwQsmWkfJmGX9E6OKBYStv0tkQx93x6
DnZVTL21mVlmLbpWOcUSfRHNyyrhxJ327Laqi6TmHdSY9M2mLTI/XY4EWGx+NTE1kg+6hS7oh8gR
yB9R9/LnbirmYXNp/Bn25clnjqjIbT5YguhWh6H9aVsuLP7ju9q9eXCtYayVDq9Gy5VmnSclfXE8
wcU7H8VPoEYVPPloDcR6F/CIasA+5RNBzMMwO5zZuyI4QaGAaVJeN9J8IJh4DuDToYQcHHrZiRmv
i1ljCEVicociBk5w6yz3bZZkse0vE+IM28B+S/xsLyHhH5GHxp/DIM1eGF4c9W58iSk/royLVya2
O8qMakli/ilZehHXU5MPLsOm3WZTvR+frCScaSkAOOjSbRt2yQffi2ksQukuN6jJWyjniQqbe4XK
/8wJjnF6h7HQlDNvatF95Ou7x0oynVAW4qnfFWPcezAOmodaV/Q0LpsCSOppSONoxsTJok58qzFc
9m0iD5+QjAXibQLIXwyUoA5vo0S7Ucxs8Sc2OMc1mt6N2K8LD6FMCiQkNwuqtEXarWQIgRdXLnwe
pHvkNzL3iy9V7dc+pf75Rga+ZVElTtOMduOjW1G17AAM8M77RkjVPphR/hCVT8RozZ7Ua1IFDthX
3CVIsb6khTrmldOvGTx13aftR9t4HFTIddWtoGzwMoED4nMEMYw8fTMn5mUdcwjc905k04QgAn5M
th+XH+FktMtdLQN0e09wlMdVDuy79tqbIQ2aCgpm1IG09ggOcFL55sH25x7CJn1F7i9U7PSKDFxv
Dlbx+rEDYRJ0ZQKZ3JhCxUj0UNQHTqeIzniM4BbAjJzhZqhNMonV/uEMAQ+zRtrMusiVzUcd/WOF
GZtNGAd4CM0Is/cy7sA3xvhr4EsR2K2WD8kK+wvCTmFGOsLmfbzUofZeLbujjW2TOqj3xW6shmGL
Y/dKSbTqQYNL4i0kyJXGipIPaITNMRSGGyVwifQ+7dC1jFWTZzlulgXQaedfnEZF5s2slSCSJjiP
7Uh9Hg5Za0y1slXeLWkg5g/6YVnpZKjqhbnv/FwvtZr//0LajN7dIPdyB1cuyJPRwGwLgznWBQ==

`pragma protect end_protected

   
endmodule
module AXI4S_INITIATOR_MIPIRX
  #(
    parameter g_DATAWIDTH = 10,
    parameter g_NUM_OF_PIXELS = 4
    )
   (
    // Input Ports
    input					   CLOCK_I,
    input					   RESET_n_I,
    input [g_NUM_OF_PIXELS * g_DATAWIDTH - 1 : 0]  DATA_I,
    input					   DATA_VALID_I,
    input					   EOF_I,
    input					   FRAME_VALID_I,
    // Output Ports
    output [g_NUM_OF_PIXELS * g_DATAWIDTH - 1 : 0] TDATA_O,
    output [g_DATAWIDTH/8 - 1 : 0]		   TSTRB_O,
    output [g_DATAWIDTH/8 - 1 : 0]		   TKEEP_O,
    output					   TVALID_O,
    output					   TLAST_O,
    output [3 : 0]				   TUSER_O  
    );

   reg						   eof_dly1;
   reg						   frame_valid_dly1;
   reg						   data_valid_dly1;
   reg [g_NUM_OF_PIXELS * g_DATAWIDTH - 1 : 0]	   data_dly1;
   wire						   tvalid_fe;
   
   assign TDATA_O		=	data_dly1;
   assign TSTRB_O    	= {(g_DATAWIDTH/8){1'b1}};
   assign TKEEP_O    	=   {(g_DATAWIDTH/8){1'b1}};
   assign TVALID_O		=	data_valid_dly1;
   assign TLAST_O		=	tvalid_fe;
   assign TUSER_O[0]		=	eof_dly1;
   assign TUSER_O[3] 	=   frame_valid_dly1;
   assign TUSER_O[2 : 1] =   2'b0;
   
   assign tvalid_fe = (data_valid_dly1 & (!DATA_VALID_I));
   
   always @(posedge CLOCK_I or negedge RESET_n_I)
     if(!RESET_n_I)
       begin
          eof_dly1			<= 0;
	  frame_valid_dly1	<= 0;
	  data_valid_dly1		<= 0;
	  data_dly1			<= {(g_NUM_OF_PIXELS *g_DATAWIDTH){1'b0}};
       end
     else
       begin
	  eof_dly1			<= EOF_I;
	  frame_valid_dly1	<= FRAME_VALID_I;
	  data_valid_dly1		<= DATA_VALID_I;
	  data_dly1			<= DATA_I;
       end 
endmodule

// --*************************************************************************************************
// -- File Name                           : axi4lite_adapter_mipi_csi_rx.v
// -- Targeted device                     : Microsemi-SoC
// -- Author                              : India Solutions Team
// --
// -- COPYRIGHT 2021 BY MICROSEMI
// -- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS FROM MICROSEMI
// -- CORP. IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM MICROSEMI FOR USE OF THIS
// -- FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND NO BACK-UP OF THE FILE SHOULD BE MADE.
// --
// --*************************************************************************************************

module axi4lite_adapter_mipi_csi_rx  
  (
   // Clock and Reset interface----------------------------------------------------
   input wire 	     aclk, // clock
   input wire 	     aresetn, // This active-low reset
   //write address channel
   input wire 	     awvalid, // AXI4-Lite write address valid. This signal indicates that valid write address and control information are available.
   output reg 	     awready, // AXI4-Lite write address ready. This signal indicates that the target is ready to accept an address and associated control signals.
   input wire [31:0] awaddr, // AXI4-Lite write address.
   //write data channel
   input wire [31:0] wdata, // AXI4-Lite write data.
   input wire 	     wvalid, // AXI4-Lite write valid.
   output reg 	     wready, // AXI4-Lite Write ready.
  //write response channel
   output  [1:0]  bresp, // AXI4-Lite write response.
   output reg 	     bvalid, // AXI4-Lite write response valid.
   input wire 	     bready, // AXI4-Lite response ready.
  //read address channel
   input wire [31:0] araddr, // AXI4-Lite read address. The read address gives the address of the first transfer in a read burst transaction.  
   input wire 	     arvalid, // AXI4-Lite read address valid. This signal indicates that the channel is signaling valid read address and control information. 
   output reg 	     arready, // AXI4-Lite response ready. This signal indicates that the slave is ready to accept an address and associated control signals.
  //read data and response channel
   input wire 	     rready, 
   output  [31:0] rdata, // AXI4-Lite read data.
   output wire [1:0] rresp, // AXI4-Lite read response.
   output reg 	     rvalid, // AXI4-Lite read valid. This signal indicates that the channel is signaling the required read data.
   //Memory interface
   output    	     mem_wr_valid,
   output  [31:0] mem_wr_addr,
   output  [31:0] mem_wr_data,
   output [31:0]     mem_rd_addr,
   input [31:0]	     mem_rd_data
   );      

   reg [31:0] 	     awaddr_reg;
   reg [31:0] 	     araddr_reg;            
   wire 	     raddr_phs_cmp;   

   //------------------------------------------------------------------------------------
   // AXI4 Lite Write Address channel
   //------------------------------------------------------------------------------------   

   ////////////////////////////////////////////////
   // AWREADY generation
   ////////////////////////////////////////////////
   always@(posedge aclk  or negedge aresetn)
     begin
	if(!aresetn)
     	  awready  <= 1'b1;
	else if (bvalid && bready)
          awready  <= 1'b1;
	else if(awvalid && awready)
          awready  <= 1'b0;
     end
   

   ////////////////////////////////////////////////
   // Storing the valid AWADDR 
   ////////////////////////////////////////////////
   always@(posedge aclk or negedge aresetn)
     begin
	if(!aresetn)
          awaddr_reg  <= 'd0;
	else if(awvalid && awready)
          awaddr_reg  <= awaddr;
     end


   //------------------------------------------------------------------------------------
   // AXI4 Lite Write Data channel
   //------------------------------------------------------------------------------------   

   ////////////////////////////////////////////////
   // Generating WREADY
   ////////////////////////////////////////////////
   always@(posedge aclk or negedge aresetn)
     begin
	if(!aresetn)
          wready  <= 1'd0;
	else if (wvalid && wready)
          wready  <= 1'd0;
	else if(awvalid && awready)
          wready  <= 1'd1;
     end


   ////////////////////////////////////////////////
   // Writing the memory with valid data 
   ////////////////////////////////////////////////   
   assign mem_wr_addr = awaddr_reg;
   assign mem_wr_data = wdata;
   assign mem_wr_valid = (wvalid == 1'b1 && wready == 1'b1);


   //------------------------------------------------------------------------------------
   // AXI4 Lite Write Response channel
   //------------------------------------------------------------------------------------   

   ////////////////////////////////////////////////
   // Generating BVALID
   ////////////////////////////////////////////////   
   always@(posedge aclk or negedge aresetn)
     begin
	if(!aresetn)
          bvalid  <= 1'd0;
	else if(bvalid == 1'b1 && bready == 1'b1)
          bvalid  <= 1'd0;
	else if(wvalid == 1'b1 && wready == 1'b1 )
          bvalid  <= 1'b1;
     end

   assign bresp = 'd0; //Giving OK response for all strobe and protection conditions
   
   //------------------------------------------------------------------------------------
   // AXI4 Lite Read Address channel
   //------------------------------------------------------------------------------------   

   ////////////////////////////////////////////////
   // Generating ARREADY
   ////////////////////////////////////////////////      
   always@(posedge aclk or negedge aresetn)
     begin
	if(!aresetn)
          arready  <= 1'd1;
	else if(rvalid && rready)
          arready  <= 1'd1;
	else if(raddr_phs_cmp)
          arready  <= 1'b0;
     end

   assign raddr_phs_cmp = (arvalid && arready); 

   ////////////////////////////////////////////////
   // Registering valid read address
   ////////////////////////////////////////////////         
   always@(posedge aclk or negedge aresetn)
     if(!aresetn)
       araddr_reg <= 'd0;
     else if(arvalid && arready)
       araddr_reg <= araddr; 

   assign mem_rd_addr = araddr_reg; 
   
   //------------------------------------------------------------------------------------
   // AXI4 Lite Read Data channel
   //------------------------------------------------------------------------------------   

   ////////////////////////////////////////////////
   // RVALID generation
   ////////////////////////////////////////////////         
   always@(posedge aclk or negedge aresetn)
     if(!aresetn)
       rvalid <= 'b0;   
     else if(arvalid && arready) 
       rvalid <= 'b1;
     else if(rvalid && rready) //hold rvalid high till rready is asserted
       rvalid <= 'b0;   

   assign rdata = mem_rd_data; //connect the the mem data directly to axi4 lite bus
   assign rresp = 2'h0; //return read OK response
      
endmodule

// --*************************************************************************************************
// -- File Name                           : write_reg_mipi_csi_rx.v
// -- Targeted device                     : Microsemi-SoC
// -- Author                              : India Solutions Team
// --
// -- COPYRIGHT 2021 BY MICROSEMI
// -- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS FROM MICROSEMI
// -- CORP. IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM MICROSEMI FOR USE OF THIS
// -- FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND NO BACK-UP OF THE FILE SHOULD BE MADE.
// --
// --*************************************************************************************************


module write_reg_mipi_csi_rx #(
	parameter CTRL_REG              = 'h4,
	parameter GLBL_INT_EN           = 'h24,
	parameter INT_STATUS            = 'h28,
	parameter INT_EN                = 'h2C
	//parameter g_CORE_EN_DIS         = 1
	)
	(
		       aclk,
		       aresetn,

		       mem_wr_valid,
		       mem_wr_addr,
		       mem_wr_data,

		       ctrl_reg,
		       glbl_int_en,
		       int_en,
		       int_status_clr
		       );
   
//`include "memory_map_mipi.v"

   // Clock and Reset interface----------------------------------------------------
   input 	     aclk; // clock
   input 	     aresetn; // This active-low reset

   //Memory interface
   input 	           mem_wr_valid;
   input [31:0]      mem_wr_addr;
   input [31:0]      mem_wr_data;

   output reg [1:0] ctrl_reg;
   output reg glbl_int_en;
   output reg [7:0]      int_en;
   output reg [7:0]  int_status_clr;
   
   ////////////////////////////////////////////////
   // Write registers
   ////////////////////////////////////////////////
   always@(posedge aclk  or negedge aresetn)
   begin
     if(!aresetn) 
	 begin
	   ctrl_reg <= 'b01;
	   //ctrl_reg <= {1'b0,g_CORE_EN_DIS[0]};
	   glbl_int_en <= 'h0;
	   int_en <= 'h0;
     end
     else if (mem_wr_valid) 
	 begin
       case (mem_wr_addr[7:0])
	 
	 CTRL_REG:
	   ctrl_reg <= mem_wr_data[1:0];

	 GLBL_INT_EN:
	   //glbl_int_en <= mem_wr_data[0:0];
	   glbl_int_en <= mem_wr_data[0];

	 INT_EN:
	   int_en <= mem_wr_data[7:0];

	 default:
	 begin
		ctrl_reg <= ctrl_reg;
	//    ctrl_reg[1] <= 'h0;	    
	//    ctrl_reg[0] <= 'h1;	    
	 end
       endcase // case (mem_wr_addr)
	 end
     else
	 begin
		ctrl_reg <= ctrl_reg;
		//ctrl_reg <= {ctrl_reg[1],g_CORE_EN_DIS};
	//    ctrl_reg[1] <= 'h0;	    
	//    ctrl_reg[0] <= 'h1;	    
	 end
   end
   


   ////////////////////////////////////////////////
   // Updating status register
   ////////////////////////////////////////////////
   always@(posedge aclk or negedge aresetn)
     if (!aresetn)
       int_status_clr <= 'h0;
     else begin
	if (mem_wr_valid && mem_wr_addr[7:0] == INT_STATUS)
	  int_status_clr <= mem_wr_data[7:0];
	else
	  int_status_clr <= 'h0;
     end


   
   // ////////////////////////////////////////////////
   // // Registering the write pulse to W1CREG1 4 stages
   // ////////////////////////////////////////////////
   // always@(posedge aclk or negedge aresetn)
   //   if (!aresetn) begin 
   // 	w1creg1_dly[0] <= 'h0;
   // 	w1creg1_dly[1] <= 'h0;
   // 	w1creg1_dly[2] <= 'h0;
   // 	w1creg1_dly[3] <= 'h0;
   //   end
   //   else begin
   // 	if (mem_wr_valid && mem_wr_addr == W1CREG1)
   // 	  w1creg1_dly[0] <= mem_wr_data;
   // 	else
   // 	  w1creg1_dly[0] <= 'h0;
   // 	w1creg1_dly[1] <= w1creg1_dly[0];
   // 	w1creg1_dly[2] <= w1creg1_dly[1];
   // 	w1creg1_dly[3] <= w1creg1_dly[2];
   //   end

   // ///////////////////////////////////////////////////
   // // Stretching the W1CREG1 write pulse to 4 clocks
   // //////////////////////////////////////////////////
   // assign w1creg1 = w1creg1_dly[0] | w1creg1_dly[1] | w1creg1_dly[2] | w1creg1_dly[3] ;
   

   
endmodule

// --*************************************************************************************************
// -- File Name                           : read_reg_mipi_csi_rx.v
// -- Targeted device                     : Microsemi-SoC
// -- Author                              : India Solutions Team
// --
// -- COPYRIGHT 2021 BY MICROSEMI
// -- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS FROM MICROSEMI
// -- CORP. IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM MICROSEMI FOR USE OF THIS
// -- FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND NO BACK-UP OF THE FILE SHOULD BE MADE.
// --
// --*************************************************************************************************

module read_reg_mipi_csi_rx #(
	parameter IP_VER                = 'h0,
	parameter CTRL_REG              = 'h4,
	parameter LANE_CONFIG           = 'h8,
	parameter DATA_WIDTH            = 'hC,
	parameter NO_OF_PIXELS          = 'h10,
	parameter NO_OF_VC              = 'h14,
	parameter INPUT_DATA_INVERT     = 'h18,
	parameter FIFO_SIZE             = 'h1C,
	parameter FRAME_RESOLUTION      = 'h20,
	parameter GLBL_INT_EN           = 'h24,
	parameter INT_STATUS            = 'h28,
	parameter INT_EN                = 'h2C,
	parameter MIPI_CLK_STATUS       = 'h30,
	parameter WORD_COUNT            = 'h58,
	parameter MIPI_CAM_DATA_TYPE    = 'h5C,
	parameter MIPI_CAM_LANES_CONFIG = 'h60
	)(
		 aclk,
		 aresetn,

		 mem_rd_addr,
		 mem_rd_data,

		      ip_ver,
		      ctrl_reg,
		      lane_config,
		      data_width,
		      no_of_pixels,
		      no_of_vc,
		      input_data_invert,
		      fifo_size,
		      frame_resolution,
		      glbl_int_en,
		      int_status,
		      int_en,
		      mipi_clk_status,
		      mipi_cam_lanes_config,
		      mipi_cam_data_type,
		      word_count	      
		 );
   
//`include "memory_map_mipi.v"   
		 
   // Clock and Reset interface----------------------------------------------------
   input 		  aclk; // clock
   input 		  aresetn; // This active-low reset
   
   //Memory interface
   input [31:0] 	  mem_rd_addr;
   output reg [31:0] 	  mem_rd_data;

   input [31:0] ip_ver;
   input [1:0] 	      ctrl_reg;   
   input [7:0] lane_config;
   input [7:0]  data_width;
   input [2:0] no_of_pixels;
   input [7:0] 	  no_of_vc;
   input  input_data_invert;
   input [3:0] 	       fifo_size;
   input [31:0]  frame_resolution;
   input [7:0]        int_status;
   input         glbl_int_en;   
   input [7:0]        int_en;   
   input    mipi_clk_status;
   input [3:0]   mipi_cam_lanes_config;
   input [7:0] mipi_cam_data_type;
   input [15:0] 	word_count;
   

   ////////////////////////////////////////////////
   // Read registers based on input address
   ////////////////////////////////////////////////
   always@(mem_rd_addr[7:0])
       case (mem_rd_addr[7:0])
	 
	 IP_VER:
	   mem_rd_data <= ip_ver;

	 CTRL_REG:
	   mem_rd_data <= ctrl_reg;

	 LANE_CONFIG:
	   mem_rd_data <= lane_config;

	 DATA_WIDTH:
	   mem_rd_data <= data_width;

	 NO_OF_PIXELS:
	   mem_rd_data <= no_of_pixels;

	 NO_OF_VC:
	   mem_rd_data <= no_of_vc;

	 INPUT_DATA_INVERT:
	   mem_rd_data <= input_data_invert;

	 FIFO_SIZE:
	   mem_rd_data <= fifo_size;

	 FRAME_RESOLUTION:
	   mem_rd_data <= frame_resolution;

	 INT_STATUS:
	   mem_rd_data <= int_status;

	 GLBL_INT_EN:
	   mem_rd_data <= glbl_int_en;
	 
	 INT_EN:
	   mem_rd_data <= int_en;
	 
	 MIPI_CLK_STATUS:
	   mem_rd_data <= mipi_clk_status;

	 MIPI_CAM_LANES_CONFIG:
	   mem_rd_data <= mipi_cam_lanes_config;

	 MIPI_CAM_DATA_TYPE:
	   mem_rd_data <= mipi_cam_data_type;

	 WORD_COUNT:
	   mem_rd_data <= word_count;
	 
	 
	 default:
	   mem_rd_data <= 32'h0;

       endcase // case (mem_rd_addr)
      
endmodule

//=================================================================================================
//-- File Name                           : interrupt_controller_mipi_csi_rx.v
//-- Targeted device                     : Microsemi-SoC
//-- Author                              : India Solutions Team
//--
//-- COPYRIGHT 2019 BY MICROSEMI
//-- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS FROM MICROSEMI
//-- CORP. IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM MICROSEMI FOR USE OF THIS
//-- FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND NO BACK-UP OF THE FILE SHOULD BE MADE.
//--
//=================================================================================================

module interrupt_controller_mipi_csi_rx 
  (
   rstn_i,
   sys_clk_i,

   interrupt_event_i,
   interrupt_en_i,
   interrupt_clear_i,
   global_interrupt_en_i,

   status_reg_o,
   interrupt_o,
   interrupt_overflow_o
   );

//`include "memory_map_mipi.v"

   
    // inputs 
    input 				 rstn_i;
    input 				 sys_clk_i;

    // input
    input [7:0] 	 interrupt_event_i;
    input [7:0] 	 interrupt_en_i;
    input [7:0] 	 interrupt_clear_i;
    input 				 global_interrupt_en_i;

    // output
    output reg [7:0] status_reg_o;
    
   output 				 interrupt_o;
   output reg [7:0]  interrupt_overflow_o;

   reg [7:0] 	 interrupt_event_dly [2:0];
   wire [7:0] 	 interrupt_event_rising_edge;
   reg [7:0] 	 event_status;   
   reg [4:0] 			 diff_cnt [7:0];
   wire [7:0] 	 diff_cnt_interrupt;   
   integer 				 i;
   genvar 				 j;
   
   ///////////////////////////////////////////////////
     //2 stage synchronizer for interrupt events
   ///////////////////////////////////////////////////   
   always@ (posedge sys_clk_i , negedge rstn_i )
     if (!rstn_i) begin
	interrupt_event_dly[0] <= 'h0;
	interrupt_event_dly[1] <= 'h0;
	interrupt_event_dly[2] <= 'h0;	
     end
     else begin
	interrupt_event_dly[0] <= interrupt_event_i;
	interrupt_event_dly[1] <= interrupt_event_dly[0];
	interrupt_event_dly[2] <= interrupt_event_dly[1];		
     end


   ///////////////////////////////////////////////////
   //Rising edge detector for interrupt event
   ///////////////////////////////////////////////////   
   for (j=0;j<8; j=j+1)     
     assign interrupt_event_rising_edge[j] = interrupt_event_dly[1][j] & !interrupt_event_dly[2][j];
   
   
   ///////////////////////////////////////////////////
   //status register based on the interrupt clear
   //command received from the processor
   ///////////////////////////////////////////////////   
   always@ (posedge sys_clk_i , negedge rstn_i )
     if (!rstn_i) 
       status_reg_o <= 'h0;
     else begin
	for (i=0;i<8; i=i+1) begin
	   if (interrupt_clear_i[i] && diff_cnt[i] == 'h1 && interrupt_event_rising_edge[i])
	     status_reg_o[i] <= 1'b1;
	   else if (interrupt_clear_i[i] && diff_cnt[i] == 'h1 && !event_status[i])
	     status_reg_o[i] <= 1'b0;	 	   
	   else if(interrupt_event_rising_edge[i] && interrupt_en_i[i] && global_interrupt_en_i)
	     status_reg_o[i] <= 1'b1;
	end
     end

   ///////////////////////////////////////////////////
   //Intermediate status register
   ///////////////////////////////////////////////////   
   always@ (posedge sys_clk_i , negedge rstn_i )
     if (!rstn_i) 
       event_status <= 'h0;
     else
       for (i=0;i<8; i=i+1)
	 if (interrupt_en_i[i] && global_interrupt_en_i)
	   event_status[i] <= interrupt_event_rising_edge[i];
   


   ///////////////////////////////////////////////////
   //Intermediate status register
   ///////////////////////////////////////////////////   
   always@ (posedge sys_clk_i , negedge rstn_i )
     for (i=0;i<8; i=i+1)     
       if (!rstn_i)
	 diff_cnt[i] <= 'h0;
       else if (interrupt_clear_i[i] && (diff_cnt[i] != 'h0) && !event_status[i]) 
	 diff_cnt[i] <= diff_cnt[i] - 1;
       else if (!interrupt_clear_i[i] && event_status[i])
	 diff_cnt[i] <= diff_cnt[i] + 1;


   ///////////////////////////////////////////////////
   //counter difference for each interrupt
   ///////////////////////////////////////////////////   
  
   for (j=0;j<8; j=j+1)     
     assign diff_cnt_interrupt[j] = |diff_cnt[j];

   ///////////////////////////////////////////////////
   //Generating interrupt based on the counter
   ///////////////////////////////////////////////////   
   assign interrupt_o = |diff_cnt_interrupt;


   ///////////////////////////////////////////////////
   //Interrupt overflow error signal generation
   //when the diff count becomes max i.e. 5'b1_1111
   //This overflow flag doesn't auto reset
   ///////////////////////////////////////////////////
   always@ (posedge sys_clk_i , negedge rstn_i )
     if (!rstn_i)
       interrupt_overflow_o <= 'h0;
     else    
       for (i=0;i<8; i=i+1)
	 if (!interrupt_overflow_o[i] && diff_cnt[i] == 5'h1f)
	   interrupt_overflow_o[i] <= 1'b1;
   


endmodule // interrupt_controller_mipi_csi_rx


