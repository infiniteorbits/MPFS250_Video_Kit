//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Sun Apr 28 14:50:46 2024
// Version: 2023.2 2023.2.0.8
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// FIC_CONVERTER
module FIC_CONVERTER(
    // Inputs
    ACLK,
    ARESETN,
    AXI4L_H264_SLAVE2_ARREADY,
    AXI4L_H264_SLAVE2_AWREADY,
    AXI4L_H264_SLAVE2_BID,
    AXI4L_H264_SLAVE2_BRESP,
    AXI4L_H264_SLAVE2_BUSER,
    AXI4L_H264_SLAVE2_BVALID,
    AXI4L_H264_SLAVE2_RDATA,
    AXI4L_H264_SLAVE2_RID,
    AXI4L_H264_SLAVE2_RLAST,
    AXI4L_H264_SLAVE2_RRESP,
    AXI4L_H264_SLAVE2_RUSER,
    AXI4L_H264_SLAVE2_RVALID,
    AXI4L_H264_SLAVE2_WREADY,
    AXI4L_IE_SLAVE3_ARREADY,
    AXI4L_IE_SLAVE3_AWREADY,
    AXI4L_IE_SLAVE3_BID,
    AXI4L_IE_SLAVE3_BRESP,
    AXI4L_IE_SLAVE3_BUSER,
    AXI4L_IE_SLAVE3_BVALID,
    AXI4L_IE_SLAVE3_RDATA,
    AXI4L_IE_SLAVE3_RID,
    AXI4L_IE_SLAVE3_RLAST,
    AXI4L_IE_SLAVE3_RRESP,
    AXI4L_IE_SLAVE3_RUSER,
    AXI4L_IE_SLAVE3_RVALID,
    AXI4L_IE_SLAVE3_WREADY,
    AXI4L_MASTER0_ARADDR,
    AXI4L_MASTER0_ARBURST,
    AXI4L_MASTER0_ARCACHE,
    AXI4L_MASTER0_ARID,
    AXI4L_MASTER0_ARLEN,
    AXI4L_MASTER0_ARLOCK,
    AXI4L_MASTER0_ARPROT,
    AXI4L_MASTER0_ARQOS,
    AXI4L_MASTER0_ARREGION,
    AXI4L_MASTER0_ARSIZE,
    AXI4L_MASTER0_ARUSER,
    AXI4L_MASTER0_ARVALID,
    AXI4L_MASTER0_AWADDR,
    AXI4L_MASTER0_AWBURST,
    AXI4L_MASTER0_AWCACHE,
    AXI4L_MASTER0_AWID,
    AXI4L_MASTER0_AWLEN,
    AXI4L_MASTER0_AWLOCK,
    AXI4L_MASTER0_AWPROT,
    AXI4L_MASTER0_AWQOS,
    AXI4L_MASTER0_AWREGION,
    AXI4L_MASTER0_AWSIZE,
    AXI4L_MASTER0_AWUSER,
    AXI4L_MASTER0_AWVALID,
    AXI4L_MASTER0_BREADY,
    AXI4L_MASTER0_RREADY,
    AXI4L_MASTER0_WDATA,
    AXI4L_MASTER0_WLAST,
    AXI4L_MASTER0_WSTRB,
    AXI4L_MASTER0_WUSER,
    AXI4L_MASTER0_WVALID,
    AXI4L_MIPI_SLAVE1_ARREADY,
    AXI4L_MIPI_SLAVE1_AWREADY,
    AXI4L_MIPI_SLAVE1_BID,
    AXI4L_MIPI_SLAVE1_BRESP,
    AXI4L_MIPI_SLAVE1_BUSER,
    AXI4L_MIPI_SLAVE1_BVALID,
    AXI4L_MIPI_SLAVE1_RDATA,
    AXI4L_MIPI_SLAVE1_RID,
    AXI4L_MIPI_SLAVE1_RLAST,
    AXI4L_MIPI_SLAVE1_RRESP,
    AXI4L_MIPI_SLAVE1_RUSER,
    AXI4L_MIPI_SLAVE1_RVALID,
    AXI4L_MIPI_SLAVE1_WREADY,
    AXI4L_OSD_SLAVE5_ARREADY,
    AXI4L_OSD_SLAVE5_AWREADY,
    AXI4L_OSD_SLAVE5_BID,
    AXI4L_OSD_SLAVE5_BRESP,
    AXI4L_OSD_SLAVE5_BUSER,
    AXI4L_OSD_SLAVE5_BVALID,
    AXI4L_OSD_SLAVE5_RDATA,
    AXI4L_OSD_SLAVE5_RID,
    AXI4L_OSD_SLAVE5_RLAST,
    AXI4L_OSD_SLAVE5_RRESP,
    AXI4L_OSD_SLAVE5_RUSER,
    AXI4L_OSD_SLAVE5_RVALID,
    AXI4L_OSD_SLAVE5_WREADY,
    AXI4L_SCALER_SLAVE4_ARREADY,
    AXI4L_SCALER_SLAVE4_AWREADY,
    AXI4L_SCALER_SLAVE4_BID,
    AXI4L_SCALER_SLAVE4_BRESP,
    AXI4L_SCALER_SLAVE4_BUSER,
    AXI4L_SCALER_SLAVE4_BVALID,
    AXI4L_SCALER_SLAVE4_RDATA,
    AXI4L_SCALER_SLAVE4_RID,
    AXI4L_SCALER_SLAVE4_RLAST,
    AXI4L_SCALER_SLAVE4_RRESP,
    AXI4L_SCALER_SLAVE4_RUSER,
    AXI4L_SCALER_SLAVE4_RVALID,
    AXI4L_SCALER_SLAVE4_WREADY,
    AXI4L_VDMA_SLAVE0_ARREADY,
    AXI4L_VDMA_SLAVE0_AWREADY,
    AXI4L_VDMA_SLAVE0_BID,
    AXI4L_VDMA_SLAVE0_BRESP,
    AXI4L_VDMA_SLAVE0_BUSER,
    AXI4L_VDMA_SLAVE0_BVALID,
    AXI4L_VDMA_SLAVE0_RDATA,
    AXI4L_VDMA_SLAVE0_RID,
    AXI4L_VDMA_SLAVE0_RLAST,
    AXI4L_VDMA_SLAVE0_RRESP,
    AXI4L_VDMA_SLAVE0_RUSER,
    AXI4L_VDMA_SLAVE0_RVALID,
    AXI4L_VDMA_SLAVE0_WREADY,
    // Outputs
    AXI4L_H264_SLAVE2_ARADDR,
    AXI4L_H264_SLAVE2_ARBURST,
    AXI4L_H264_SLAVE2_ARCACHE,
    AXI4L_H264_SLAVE2_ARID,
    AXI4L_H264_SLAVE2_ARLEN,
    AXI4L_H264_SLAVE2_ARLOCK,
    AXI4L_H264_SLAVE2_ARPROT,
    AXI4L_H264_SLAVE2_ARQOS,
    AXI4L_H264_SLAVE2_ARREGION,
    AXI4L_H264_SLAVE2_ARSIZE,
    AXI4L_H264_SLAVE2_ARUSER,
    AXI4L_H264_SLAVE2_ARVALID,
    AXI4L_H264_SLAVE2_AWADDR,
    AXI4L_H264_SLAVE2_AWBURST,
    AXI4L_H264_SLAVE2_AWCACHE,
    AXI4L_H264_SLAVE2_AWID,
    AXI4L_H264_SLAVE2_AWLEN,
    AXI4L_H264_SLAVE2_AWLOCK,
    AXI4L_H264_SLAVE2_AWPROT,
    AXI4L_H264_SLAVE2_AWQOS,
    AXI4L_H264_SLAVE2_AWREGION,
    AXI4L_H264_SLAVE2_AWSIZE,
    AXI4L_H264_SLAVE2_AWUSER,
    AXI4L_H264_SLAVE2_AWVALID,
    AXI4L_H264_SLAVE2_BREADY,
    AXI4L_H264_SLAVE2_RREADY,
    AXI4L_H264_SLAVE2_WDATA,
    AXI4L_H264_SLAVE2_WLAST,
    AXI4L_H264_SLAVE2_WSTRB,
    AXI4L_H264_SLAVE2_WUSER,
    AXI4L_H264_SLAVE2_WVALID,
    AXI4L_IE_SLAVE3_ARADDR,
    AXI4L_IE_SLAVE3_ARBURST,
    AXI4L_IE_SLAVE3_ARCACHE,
    AXI4L_IE_SLAVE3_ARID,
    AXI4L_IE_SLAVE3_ARLEN,
    AXI4L_IE_SLAVE3_ARLOCK,
    AXI4L_IE_SLAVE3_ARPROT,
    AXI4L_IE_SLAVE3_ARQOS,
    AXI4L_IE_SLAVE3_ARREGION,
    AXI4L_IE_SLAVE3_ARSIZE,
    AXI4L_IE_SLAVE3_ARUSER,
    AXI4L_IE_SLAVE3_ARVALID,
    AXI4L_IE_SLAVE3_AWADDR,
    AXI4L_IE_SLAVE3_AWBURST,
    AXI4L_IE_SLAVE3_AWCACHE,
    AXI4L_IE_SLAVE3_AWID,
    AXI4L_IE_SLAVE3_AWLEN,
    AXI4L_IE_SLAVE3_AWLOCK,
    AXI4L_IE_SLAVE3_AWPROT,
    AXI4L_IE_SLAVE3_AWQOS,
    AXI4L_IE_SLAVE3_AWREGION,
    AXI4L_IE_SLAVE3_AWSIZE,
    AXI4L_IE_SLAVE3_AWUSER,
    AXI4L_IE_SLAVE3_AWVALID,
    AXI4L_IE_SLAVE3_BREADY,
    AXI4L_IE_SLAVE3_RREADY,
    AXI4L_IE_SLAVE3_WDATA,
    AXI4L_IE_SLAVE3_WLAST,
    AXI4L_IE_SLAVE3_WSTRB,
    AXI4L_IE_SLAVE3_WUSER,
    AXI4L_IE_SLAVE3_WVALID,
    AXI4L_MASTER0_ARREADY,
    AXI4L_MASTER0_AWREADY,
    AXI4L_MASTER0_BID,
    AXI4L_MASTER0_BRESP,
    AXI4L_MASTER0_BUSER,
    AXI4L_MASTER0_BVALID,
    AXI4L_MASTER0_RDATA,
    AXI4L_MASTER0_RID,
    AXI4L_MASTER0_RLAST,
    AXI4L_MASTER0_RRESP,
    AXI4L_MASTER0_RUSER,
    AXI4L_MASTER0_RVALID,
    AXI4L_MASTER0_WREADY,
    AXI4L_MIPI_SLAVE1_ARADDR,
    AXI4L_MIPI_SLAVE1_ARBURST,
    AXI4L_MIPI_SLAVE1_ARCACHE,
    AXI4L_MIPI_SLAVE1_ARID,
    AXI4L_MIPI_SLAVE1_ARLEN,
    AXI4L_MIPI_SLAVE1_ARLOCK,
    AXI4L_MIPI_SLAVE1_ARPROT,
    AXI4L_MIPI_SLAVE1_ARQOS,
    AXI4L_MIPI_SLAVE1_ARREGION,
    AXI4L_MIPI_SLAVE1_ARSIZE,
    AXI4L_MIPI_SLAVE1_ARUSER,
    AXI4L_MIPI_SLAVE1_ARVALID,
    AXI4L_MIPI_SLAVE1_AWADDR,
    AXI4L_MIPI_SLAVE1_AWBURST,
    AXI4L_MIPI_SLAVE1_AWCACHE,
    AXI4L_MIPI_SLAVE1_AWID,
    AXI4L_MIPI_SLAVE1_AWLEN,
    AXI4L_MIPI_SLAVE1_AWLOCK,
    AXI4L_MIPI_SLAVE1_AWPROT,
    AXI4L_MIPI_SLAVE1_AWQOS,
    AXI4L_MIPI_SLAVE1_AWREGION,
    AXI4L_MIPI_SLAVE1_AWSIZE,
    AXI4L_MIPI_SLAVE1_AWUSER,
    AXI4L_MIPI_SLAVE1_AWVALID,
    AXI4L_MIPI_SLAVE1_BREADY,
    AXI4L_MIPI_SLAVE1_RREADY,
    AXI4L_MIPI_SLAVE1_WDATA,
    AXI4L_MIPI_SLAVE1_WLAST,
    AXI4L_MIPI_SLAVE1_WSTRB,
    AXI4L_MIPI_SLAVE1_WUSER,
    AXI4L_MIPI_SLAVE1_WVALID,
    AXI4L_OSD_SLAVE5_ARADDR,
    AXI4L_OSD_SLAVE5_ARBURST,
    AXI4L_OSD_SLAVE5_ARCACHE,
    AXI4L_OSD_SLAVE5_ARID,
    AXI4L_OSD_SLAVE5_ARLEN,
    AXI4L_OSD_SLAVE5_ARLOCK,
    AXI4L_OSD_SLAVE5_ARPROT,
    AXI4L_OSD_SLAVE5_ARQOS,
    AXI4L_OSD_SLAVE5_ARREGION,
    AXI4L_OSD_SLAVE5_ARSIZE,
    AXI4L_OSD_SLAVE5_ARUSER,
    AXI4L_OSD_SLAVE5_ARVALID,
    AXI4L_OSD_SLAVE5_AWADDR,
    AXI4L_OSD_SLAVE5_AWBURST,
    AXI4L_OSD_SLAVE5_AWCACHE,
    AXI4L_OSD_SLAVE5_AWID,
    AXI4L_OSD_SLAVE5_AWLEN,
    AXI4L_OSD_SLAVE5_AWLOCK,
    AXI4L_OSD_SLAVE5_AWPROT,
    AXI4L_OSD_SLAVE5_AWQOS,
    AXI4L_OSD_SLAVE5_AWREGION,
    AXI4L_OSD_SLAVE5_AWSIZE,
    AXI4L_OSD_SLAVE5_AWUSER,
    AXI4L_OSD_SLAVE5_AWVALID,
    AXI4L_OSD_SLAVE5_BREADY,
    AXI4L_OSD_SLAVE5_RREADY,
    AXI4L_OSD_SLAVE5_WDATA,
    AXI4L_OSD_SLAVE5_WLAST,
    AXI4L_OSD_SLAVE5_WSTRB,
    AXI4L_OSD_SLAVE5_WUSER,
    AXI4L_OSD_SLAVE5_WVALID,
    AXI4L_SCALER_SLAVE4_ARADDR,
    AXI4L_SCALER_SLAVE4_ARBURST,
    AXI4L_SCALER_SLAVE4_ARCACHE,
    AXI4L_SCALER_SLAVE4_ARID,
    AXI4L_SCALER_SLAVE4_ARLEN,
    AXI4L_SCALER_SLAVE4_ARLOCK,
    AXI4L_SCALER_SLAVE4_ARPROT,
    AXI4L_SCALER_SLAVE4_ARQOS,
    AXI4L_SCALER_SLAVE4_ARREGION,
    AXI4L_SCALER_SLAVE4_ARSIZE,
    AXI4L_SCALER_SLAVE4_ARUSER,
    AXI4L_SCALER_SLAVE4_ARVALID,
    AXI4L_SCALER_SLAVE4_AWADDR,
    AXI4L_SCALER_SLAVE4_AWBURST,
    AXI4L_SCALER_SLAVE4_AWCACHE,
    AXI4L_SCALER_SLAVE4_AWID,
    AXI4L_SCALER_SLAVE4_AWLEN,
    AXI4L_SCALER_SLAVE4_AWLOCK,
    AXI4L_SCALER_SLAVE4_AWPROT,
    AXI4L_SCALER_SLAVE4_AWQOS,
    AXI4L_SCALER_SLAVE4_AWREGION,
    AXI4L_SCALER_SLAVE4_AWSIZE,
    AXI4L_SCALER_SLAVE4_AWUSER,
    AXI4L_SCALER_SLAVE4_AWVALID,
    AXI4L_SCALER_SLAVE4_BREADY,
    AXI4L_SCALER_SLAVE4_RREADY,
    AXI4L_SCALER_SLAVE4_WDATA,
    AXI4L_SCALER_SLAVE4_WLAST,
    AXI4L_SCALER_SLAVE4_WSTRB,
    AXI4L_SCALER_SLAVE4_WUSER,
    AXI4L_SCALER_SLAVE4_WVALID,
    AXI4L_VDMA_SLAVE0_ARADDR,
    AXI4L_VDMA_SLAVE0_ARBURST,
    AXI4L_VDMA_SLAVE0_ARCACHE,
    AXI4L_VDMA_SLAVE0_ARID,
    AXI4L_VDMA_SLAVE0_ARLEN,
    AXI4L_VDMA_SLAVE0_ARLOCK,
    AXI4L_VDMA_SLAVE0_ARPROT,
    AXI4L_VDMA_SLAVE0_ARQOS,
    AXI4L_VDMA_SLAVE0_ARREGION,
    AXI4L_VDMA_SLAVE0_ARSIZE,
    AXI4L_VDMA_SLAVE0_ARUSER,
    AXI4L_VDMA_SLAVE0_ARVALID,
    AXI4L_VDMA_SLAVE0_AWADDR,
    AXI4L_VDMA_SLAVE0_AWBURST,
    AXI4L_VDMA_SLAVE0_AWCACHE,
    AXI4L_VDMA_SLAVE0_AWID,
    AXI4L_VDMA_SLAVE0_AWLEN,
    AXI4L_VDMA_SLAVE0_AWLOCK,
    AXI4L_VDMA_SLAVE0_AWPROT,
    AXI4L_VDMA_SLAVE0_AWQOS,
    AXI4L_VDMA_SLAVE0_AWREGION,
    AXI4L_VDMA_SLAVE0_AWSIZE,
    AXI4L_VDMA_SLAVE0_AWUSER,
    AXI4L_VDMA_SLAVE0_AWVALID,
    AXI4L_VDMA_SLAVE0_BREADY,
    AXI4L_VDMA_SLAVE0_RREADY,
    AXI4L_VDMA_SLAVE0_WDATA,
    AXI4L_VDMA_SLAVE0_WLAST,
    AXI4L_VDMA_SLAVE0_WSTRB,
    AXI4L_VDMA_SLAVE0_WUSER,
    AXI4L_VDMA_SLAVE0_WVALID
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input         ACLK;
input         ARESETN;
input         AXI4L_H264_SLAVE2_ARREADY;
input         AXI4L_H264_SLAVE2_AWREADY;
input  [8:0]  AXI4L_H264_SLAVE2_BID;
input  [1:0]  AXI4L_H264_SLAVE2_BRESP;
input  [0:0]  AXI4L_H264_SLAVE2_BUSER;
input         AXI4L_H264_SLAVE2_BVALID;
input  [31:0] AXI4L_H264_SLAVE2_RDATA;
input  [8:0]  AXI4L_H264_SLAVE2_RID;
input         AXI4L_H264_SLAVE2_RLAST;
input  [1:0]  AXI4L_H264_SLAVE2_RRESP;
input  [0:0]  AXI4L_H264_SLAVE2_RUSER;
input         AXI4L_H264_SLAVE2_RVALID;
input         AXI4L_H264_SLAVE2_WREADY;
input         AXI4L_IE_SLAVE3_ARREADY;
input         AXI4L_IE_SLAVE3_AWREADY;
input  [8:0]  AXI4L_IE_SLAVE3_BID;
input  [1:0]  AXI4L_IE_SLAVE3_BRESP;
input  [0:0]  AXI4L_IE_SLAVE3_BUSER;
input         AXI4L_IE_SLAVE3_BVALID;
input  [31:0] AXI4L_IE_SLAVE3_RDATA;
input  [8:0]  AXI4L_IE_SLAVE3_RID;
input         AXI4L_IE_SLAVE3_RLAST;
input  [1:0]  AXI4L_IE_SLAVE3_RRESP;
input  [0:0]  AXI4L_IE_SLAVE3_RUSER;
input         AXI4L_IE_SLAVE3_RVALID;
input         AXI4L_IE_SLAVE3_WREADY;
input  [37:0] AXI4L_MASTER0_ARADDR;
input  [1:0]  AXI4L_MASTER0_ARBURST;
input  [3:0]  AXI4L_MASTER0_ARCACHE;
input  [7:0]  AXI4L_MASTER0_ARID;
input  [7:0]  AXI4L_MASTER0_ARLEN;
input  [1:0]  AXI4L_MASTER0_ARLOCK;
input  [2:0]  AXI4L_MASTER0_ARPROT;
input  [3:0]  AXI4L_MASTER0_ARQOS;
input  [3:0]  AXI4L_MASTER0_ARREGION;
input  [2:0]  AXI4L_MASTER0_ARSIZE;
input  [0:0]  AXI4L_MASTER0_ARUSER;
input         AXI4L_MASTER0_ARVALID;
input  [37:0] AXI4L_MASTER0_AWADDR;
input  [1:0]  AXI4L_MASTER0_AWBURST;
input  [3:0]  AXI4L_MASTER0_AWCACHE;
input  [7:0]  AXI4L_MASTER0_AWID;
input  [7:0]  AXI4L_MASTER0_AWLEN;
input  [1:0]  AXI4L_MASTER0_AWLOCK;
input  [2:0]  AXI4L_MASTER0_AWPROT;
input  [3:0]  AXI4L_MASTER0_AWQOS;
input  [3:0]  AXI4L_MASTER0_AWREGION;
input  [2:0]  AXI4L_MASTER0_AWSIZE;
input  [0:0]  AXI4L_MASTER0_AWUSER;
input         AXI4L_MASTER0_AWVALID;
input         AXI4L_MASTER0_BREADY;
input         AXI4L_MASTER0_RREADY;
input  [63:0] AXI4L_MASTER0_WDATA;
input         AXI4L_MASTER0_WLAST;
input  [7:0]  AXI4L_MASTER0_WSTRB;
input  [0:0]  AXI4L_MASTER0_WUSER;
input         AXI4L_MASTER0_WVALID;
input         AXI4L_MIPI_SLAVE1_ARREADY;
input         AXI4L_MIPI_SLAVE1_AWREADY;
input  [8:0]  AXI4L_MIPI_SLAVE1_BID;
input  [1:0]  AXI4L_MIPI_SLAVE1_BRESP;
input  [0:0]  AXI4L_MIPI_SLAVE1_BUSER;
input         AXI4L_MIPI_SLAVE1_BVALID;
input  [31:0] AXI4L_MIPI_SLAVE1_RDATA;
input  [8:0]  AXI4L_MIPI_SLAVE1_RID;
input         AXI4L_MIPI_SLAVE1_RLAST;
input  [1:0]  AXI4L_MIPI_SLAVE1_RRESP;
input  [0:0]  AXI4L_MIPI_SLAVE1_RUSER;
input         AXI4L_MIPI_SLAVE1_RVALID;
input         AXI4L_MIPI_SLAVE1_WREADY;
input         AXI4L_OSD_SLAVE5_ARREADY;
input         AXI4L_OSD_SLAVE5_AWREADY;
input  [8:0]  AXI4L_OSD_SLAVE5_BID;
input  [1:0]  AXI4L_OSD_SLAVE5_BRESP;
input  [0:0]  AXI4L_OSD_SLAVE5_BUSER;
input         AXI4L_OSD_SLAVE5_BVALID;
input  [63:0] AXI4L_OSD_SLAVE5_RDATA;
input  [8:0]  AXI4L_OSD_SLAVE5_RID;
input         AXI4L_OSD_SLAVE5_RLAST;
input  [1:0]  AXI4L_OSD_SLAVE5_RRESP;
input  [0:0]  AXI4L_OSD_SLAVE5_RUSER;
input         AXI4L_OSD_SLAVE5_RVALID;
input         AXI4L_OSD_SLAVE5_WREADY;
input         AXI4L_SCALER_SLAVE4_ARREADY;
input         AXI4L_SCALER_SLAVE4_AWREADY;
input  [8:0]  AXI4L_SCALER_SLAVE4_BID;
input  [1:0]  AXI4L_SCALER_SLAVE4_BRESP;
input  [0:0]  AXI4L_SCALER_SLAVE4_BUSER;
input         AXI4L_SCALER_SLAVE4_BVALID;
input  [63:0] AXI4L_SCALER_SLAVE4_RDATA;
input  [8:0]  AXI4L_SCALER_SLAVE4_RID;
input         AXI4L_SCALER_SLAVE4_RLAST;
input  [1:0]  AXI4L_SCALER_SLAVE4_RRESP;
input  [0:0]  AXI4L_SCALER_SLAVE4_RUSER;
input         AXI4L_SCALER_SLAVE4_RVALID;
input         AXI4L_SCALER_SLAVE4_WREADY;
input         AXI4L_VDMA_SLAVE0_ARREADY;
input         AXI4L_VDMA_SLAVE0_AWREADY;
input  [8:0]  AXI4L_VDMA_SLAVE0_BID;
input  [1:0]  AXI4L_VDMA_SLAVE0_BRESP;
input  [0:0]  AXI4L_VDMA_SLAVE0_BUSER;
input         AXI4L_VDMA_SLAVE0_BVALID;
input  [31:0] AXI4L_VDMA_SLAVE0_RDATA;
input  [8:0]  AXI4L_VDMA_SLAVE0_RID;
input         AXI4L_VDMA_SLAVE0_RLAST;
input  [1:0]  AXI4L_VDMA_SLAVE0_RRESP;
input  [0:0]  AXI4L_VDMA_SLAVE0_RUSER;
input         AXI4L_VDMA_SLAVE0_RVALID;
input         AXI4L_VDMA_SLAVE0_WREADY;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [37:0] AXI4L_H264_SLAVE2_ARADDR;
output [1:0]  AXI4L_H264_SLAVE2_ARBURST;
output [3:0]  AXI4L_H264_SLAVE2_ARCACHE;
output [8:0]  AXI4L_H264_SLAVE2_ARID;
output [7:0]  AXI4L_H264_SLAVE2_ARLEN;
output [1:0]  AXI4L_H264_SLAVE2_ARLOCK;
output [2:0]  AXI4L_H264_SLAVE2_ARPROT;
output [3:0]  AXI4L_H264_SLAVE2_ARQOS;
output [3:0]  AXI4L_H264_SLAVE2_ARREGION;
output [2:0]  AXI4L_H264_SLAVE2_ARSIZE;
output [0:0]  AXI4L_H264_SLAVE2_ARUSER;
output        AXI4L_H264_SLAVE2_ARVALID;
output [37:0] AXI4L_H264_SLAVE2_AWADDR;
output [1:0]  AXI4L_H264_SLAVE2_AWBURST;
output [3:0]  AXI4L_H264_SLAVE2_AWCACHE;
output [8:0]  AXI4L_H264_SLAVE2_AWID;
output [7:0]  AXI4L_H264_SLAVE2_AWLEN;
output [1:0]  AXI4L_H264_SLAVE2_AWLOCK;
output [2:0]  AXI4L_H264_SLAVE2_AWPROT;
output [3:0]  AXI4L_H264_SLAVE2_AWQOS;
output [3:0]  AXI4L_H264_SLAVE2_AWREGION;
output [2:0]  AXI4L_H264_SLAVE2_AWSIZE;
output [0:0]  AXI4L_H264_SLAVE2_AWUSER;
output        AXI4L_H264_SLAVE2_AWVALID;
output        AXI4L_H264_SLAVE2_BREADY;
output        AXI4L_H264_SLAVE2_RREADY;
output [31:0] AXI4L_H264_SLAVE2_WDATA;
output        AXI4L_H264_SLAVE2_WLAST;
output [3:0]  AXI4L_H264_SLAVE2_WSTRB;
output [0:0]  AXI4L_H264_SLAVE2_WUSER;
output        AXI4L_H264_SLAVE2_WVALID;
output [37:0] AXI4L_IE_SLAVE3_ARADDR;
output [1:0]  AXI4L_IE_SLAVE3_ARBURST;
output [3:0]  AXI4L_IE_SLAVE3_ARCACHE;
output [8:0]  AXI4L_IE_SLAVE3_ARID;
output [7:0]  AXI4L_IE_SLAVE3_ARLEN;
output [1:0]  AXI4L_IE_SLAVE3_ARLOCK;
output [2:0]  AXI4L_IE_SLAVE3_ARPROT;
output [3:0]  AXI4L_IE_SLAVE3_ARQOS;
output [3:0]  AXI4L_IE_SLAVE3_ARREGION;
output [2:0]  AXI4L_IE_SLAVE3_ARSIZE;
output [0:0]  AXI4L_IE_SLAVE3_ARUSER;
output        AXI4L_IE_SLAVE3_ARVALID;
output [37:0] AXI4L_IE_SLAVE3_AWADDR;
output [1:0]  AXI4L_IE_SLAVE3_AWBURST;
output [3:0]  AXI4L_IE_SLAVE3_AWCACHE;
output [8:0]  AXI4L_IE_SLAVE3_AWID;
output [7:0]  AXI4L_IE_SLAVE3_AWLEN;
output [1:0]  AXI4L_IE_SLAVE3_AWLOCK;
output [2:0]  AXI4L_IE_SLAVE3_AWPROT;
output [3:0]  AXI4L_IE_SLAVE3_AWQOS;
output [3:0]  AXI4L_IE_SLAVE3_AWREGION;
output [2:0]  AXI4L_IE_SLAVE3_AWSIZE;
output [0:0]  AXI4L_IE_SLAVE3_AWUSER;
output        AXI4L_IE_SLAVE3_AWVALID;
output        AXI4L_IE_SLAVE3_BREADY;
output        AXI4L_IE_SLAVE3_RREADY;
output [31:0] AXI4L_IE_SLAVE3_WDATA;
output        AXI4L_IE_SLAVE3_WLAST;
output [3:0]  AXI4L_IE_SLAVE3_WSTRB;
output [0:0]  AXI4L_IE_SLAVE3_WUSER;
output        AXI4L_IE_SLAVE3_WVALID;
output        AXI4L_MASTER0_ARREADY;
output        AXI4L_MASTER0_AWREADY;
output [7:0]  AXI4L_MASTER0_BID;
output [1:0]  AXI4L_MASTER0_BRESP;
output [0:0]  AXI4L_MASTER0_BUSER;
output        AXI4L_MASTER0_BVALID;
output [63:0] AXI4L_MASTER0_RDATA;
output [7:0]  AXI4L_MASTER0_RID;
output        AXI4L_MASTER0_RLAST;
output [1:0]  AXI4L_MASTER0_RRESP;
output [0:0]  AXI4L_MASTER0_RUSER;
output        AXI4L_MASTER0_RVALID;
output        AXI4L_MASTER0_WREADY;
output [37:0] AXI4L_MIPI_SLAVE1_ARADDR;
output [1:0]  AXI4L_MIPI_SLAVE1_ARBURST;
output [3:0]  AXI4L_MIPI_SLAVE1_ARCACHE;
output [8:0]  AXI4L_MIPI_SLAVE1_ARID;
output [7:0]  AXI4L_MIPI_SLAVE1_ARLEN;
output [1:0]  AXI4L_MIPI_SLAVE1_ARLOCK;
output [2:0]  AXI4L_MIPI_SLAVE1_ARPROT;
output [3:0]  AXI4L_MIPI_SLAVE1_ARQOS;
output [3:0]  AXI4L_MIPI_SLAVE1_ARREGION;
output [2:0]  AXI4L_MIPI_SLAVE1_ARSIZE;
output [0:0]  AXI4L_MIPI_SLAVE1_ARUSER;
output        AXI4L_MIPI_SLAVE1_ARVALID;
output [37:0] AXI4L_MIPI_SLAVE1_AWADDR;
output [1:0]  AXI4L_MIPI_SLAVE1_AWBURST;
output [3:0]  AXI4L_MIPI_SLAVE1_AWCACHE;
output [8:0]  AXI4L_MIPI_SLAVE1_AWID;
output [7:0]  AXI4L_MIPI_SLAVE1_AWLEN;
output [1:0]  AXI4L_MIPI_SLAVE1_AWLOCK;
output [2:0]  AXI4L_MIPI_SLAVE1_AWPROT;
output [3:0]  AXI4L_MIPI_SLAVE1_AWQOS;
output [3:0]  AXI4L_MIPI_SLAVE1_AWREGION;
output [2:0]  AXI4L_MIPI_SLAVE1_AWSIZE;
output [0:0]  AXI4L_MIPI_SLAVE1_AWUSER;
output        AXI4L_MIPI_SLAVE1_AWVALID;
output        AXI4L_MIPI_SLAVE1_BREADY;
output        AXI4L_MIPI_SLAVE1_RREADY;
output [31:0] AXI4L_MIPI_SLAVE1_WDATA;
output        AXI4L_MIPI_SLAVE1_WLAST;
output [3:0]  AXI4L_MIPI_SLAVE1_WSTRB;
output [0:0]  AXI4L_MIPI_SLAVE1_WUSER;
output        AXI4L_MIPI_SLAVE1_WVALID;
output [37:0] AXI4L_OSD_SLAVE5_ARADDR;
output [1:0]  AXI4L_OSD_SLAVE5_ARBURST;
output [3:0]  AXI4L_OSD_SLAVE5_ARCACHE;
output [8:0]  AXI4L_OSD_SLAVE5_ARID;
output [7:0]  AXI4L_OSD_SLAVE5_ARLEN;
output [1:0]  AXI4L_OSD_SLAVE5_ARLOCK;
output [2:0]  AXI4L_OSD_SLAVE5_ARPROT;
output [3:0]  AXI4L_OSD_SLAVE5_ARQOS;
output [3:0]  AXI4L_OSD_SLAVE5_ARREGION;
output [2:0]  AXI4L_OSD_SLAVE5_ARSIZE;
output [0:0]  AXI4L_OSD_SLAVE5_ARUSER;
output        AXI4L_OSD_SLAVE5_ARVALID;
output [37:0] AXI4L_OSD_SLAVE5_AWADDR;
output [1:0]  AXI4L_OSD_SLAVE5_AWBURST;
output [3:0]  AXI4L_OSD_SLAVE5_AWCACHE;
output [8:0]  AXI4L_OSD_SLAVE5_AWID;
output [7:0]  AXI4L_OSD_SLAVE5_AWLEN;
output [1:0]  AXI4L_OSD_SLAVE5_AWLOCK;
output [2:0]  AXI4L_OSD_SLAVE5_AWPROT;
output [3:0]  AXI4L_OSD_SLAVE5_AWQOS;
output [3:0]  AXI4L_OSD_SLAVE5_AWREGION;
output [2:0]  AXI4L_OSD_SLAVE5_AWSIZE;
output [0:0]  AXI4L_OSD_SLAVE5_AWUSER;
output        AXI4L_OSD_SLAVE5_AWVALID;
output        AXI4L_OSD_SLAVE5_BREADY;
output        AXI4L_OSD_SLAVE5_RREADY;
output [63:0] AXI4L_OSD_SLAVE5_WDATA;
output        AXI4L_OSD_SLAVE5_WLAST;
output [7:0]  AXI4L_OSD_SLAVE5_WSTRB;
output [0:0]  AXI4L_OSD_SLAVE5_WUSER;
output        AXI4L_OSD_SLAVE5_WVALID;
output [37:0] AXI4L_SCALER_SLAVE4_ARADDR;
output [1:0]  AXI4L_SCALER_SLAVE4_ARBURST;
output [3:0]  AXI4L_SCALER_SLAVE4_ARCACHE;
output [8:0]  AXI4L_SCALER_SLAVE4_ARID;
output [7:0]  AXI4L_SCALER_SLAVE4_ARLEN;
output [1:0]  AXI4L_SCALER_SLAVE4_ARLOCK;
output [2:0]  AXI4L_SCALER_SLAVE4_ARPROT;
output [3:0]  AXI4L_SCALER_SLAVE4_ARQOS;
output [3:0]  AXI4L_SCALER_SLAVE4_ARREGION;
output [2:0]  AXI4L_SCALER_SLAVE4_ARSIZE;
output [0:0]  AXI4L_SCALER_SLAVE4_ARUSER;
output        AXI4L_SCALER_SLAVE4_ARVALID;
output [37:0] AXI4L_SCALER_SLAVE4_AWADDR;
output [1:0]  AXI4L_SCALER_SLAVE4_AWBURST;
output [3:0]  AXI4L_SCALER_SLAVE4_AWCACHE;
output [8:0]  AXI4L_SCALER_SLAVE4_AWID;
output [7:0]  AXI4L_SCALER_SLAVE4_AWLEN;
output [1:0]  AXI4L_SCALER_SLAVE4_AWLOCK;
output [2:0]  AXI4L_SCALER_SLAVE4_AWPROT;
output [3:0]  AXI4L_SCALER_SLAVE4_AWQOS;
output [3:0]  AXI4L_SCALER_SLAVE4_AWREGION;
output [2:0]  AXI4L_SCALER_SLAVE4_AWSIZE;
output [0:0]  AXI4L_SCALER_SLAVE4_AWUSER;
output        AXI4L_SCALER_SLAVE4_AWVALID;
output        AXI4L_SCALER_SLAVE4_BREADY;
output        AXI4L_SCALER_SLAVE4_RREADY;
output [63:0] AXI4L_SCALER_SLAVE4_WDATA;
output        AXI4L_SCALER_SLAVE4_WLAST;
output [7:0]  AXI4L_SCALER_SLAVE4_WSTRB;
output [0:0]  AXI4L_SCALER_SLAVE4_WUSER;
output        AXI4L_SCALER_SLAVE4_WVALID;
output [37:0] AXI4L_VDMA_SLAVE0_ARADDR;
output [1:0]  AXI4L_VDMA_SLAVE0_ARBURST;
output [3:0]  AXI4L_VDMA_SLAVE0_ARCACHE;
output [8:0]  AXI4L_VDMA_SLAVE0_ARID;
output [7:0]  AXI4L_VDMA_SLAVE0_ARLEN;
output [1:0]  AXI4L_VDMA_SLAVE0_ARLOCK;
output [2:0]  AXI4L_VDMA_SLAVE0_ARPROT;
output [3:0]  AXI4L_VDMA_SLAVE0_ARQOS;
output [3:0]  AXI4L_VDMA_SLAVE0_ARREGION;
output [2:0]  AXI4L_VDMA_SLAVE0_ARSIZE;
output [0:0]  AXI4L_VDMA_SLAVE0_ARUSER;
output        AXI4L_VDMA_SLAVE0_ARVALID;
output [37:0] AXI4L_VDMA_SLAVE0_AWADDR;
output [1:0]  AXI4L_VDMA_SLAVE0_AWBURST;
output [3:0]  AXI4L_VDMA_SLAVE0_AWCACHE;
output [8:0]  AXI4L_VDMA_SLAVE0_AWID;
output [7:0]  AXI4L_VDMA_SLAVE0_AWLEN;
output [1:0]  AXI4L_VDMA_SLAVE0_AWLOCK;
output [2:0]  AXI4L_VDMA_SLAVE0_AWPROT;
output [3:0]  AXI4L_VDMA_SLAVE0_AWQOS;
output [3:0]  AXI4L_VDMA_SLAVE0_AWREGION;
output [2:0]  AXI4L_VDMA_SLAVE0_AWSIZE;
output [0:0]  AXI4L_VDMA_SLAVE0_AWUSER;
output        AXI4L_VDMA_SLAVE0_AWVALID;
output        AXI4L_VDMA_SLAVE0_BREADY;
output        AXI4L_VDMA_SLAVE0_RREADY;
output [31:0] AXI4L_VDMA_SLAVE0_WDATA;
output        AXI4L_VDMA_SLAVE0_WLAST;
output [3:0]  AXI4L_VDMA_SLAVE0_WSTRB;
output [0:0]  AXI4L_VDMA_SLAVE0_WUSER;
output        AXI4L_VDMA_SLAVE0_WVALID;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire          ACLK;
wire          ARESETN;
wire   [37:0] AXI4L_MASTER0_ARADDR;
wire   [1:0]  AXI4L_MASTER0_ARBURST;
wire   [3:0]  AXI4L_MASTER0_ARCACHE;
wire   [7:0]  AXI4L_MASTER0_ARID;
wire   [7:0]  AXI4L_MASTER0_ARLEN;
wire   [1:0]  AXI4L_MASTER0_ARLOCK;
wire   [2:0]  AXI4L_MASTER0_ARPROT;
wire   [3:0]  AXI4L_MASTER0_ARQOS;
wire          AXI4L_ARREADY;
wire   [3:0]  AXI4L_MASTER0_ARREGION;
wire   [2:0]  AXI4L_MASTER0_ARSIZE;
wire   [0:0]  AXI4L_MASTER0_ARUSER;
wire          AXI4L_MASTER0_ARVALID;
wire   [37:0] AXI4L_MASTER0_AWADDR;
wire   [1:0]  AXI4L_MASTER0_AWBURST;
wire   [3:0]  AXI4L_MASTER0_AWCACHE;
wire   [7:0]  AXI4L_MASTER0_AWID;
wire   [7:0]  AXI4L_MASTER0_AWLEN;
wire   [1:0]  AXI4L_MASTER0_AWLOCK;
wire   [2:0]  AXI4L_MASTER0_AWPROT;
wire   [3:0]  AXI4L_MASTER0_AWQOS;
wire          AXI4L_AWREADY;
wire   [3:0]  AXI4L_MASTER0_AWREGION;
wire   [2:0]  AXI4L_MASTER0_AWSIZE;
wire   [0:0]  AXI4L_MASTER0_AWUSER;
wire          AXI4L_MASTER0_AWVALID;
wire   [7:0]  AXI4L_BID;
wire          AXI4L_MASTER0_BREADY;
wire   [1:0]  AXI4L_BRESP;
wire   [0:0]  AXI4L_BUSER;
wire          AXI4L_BVALID;
wire   [63:0] AXI4L_RDATA;
wire   [7:0]  AXI4L_RID;
wire          AXI4L_RLAST;
wire          AXI4L_MASTER0_RREADY;
wire   [1:0]  AXI4L_RRESP;
wire   [0:0]  AXI4L_RUSER;
wire          AXI4L_RVALID;
wire   [63:0] AXI4L_MASTER0_WDATA;
wire          AXI4L_MASTER0_WLAST;
wire          AXI4L_WREADY;
wire   [7:0]  AXI4L_MASTER0_WSTRB;
wire   [0:0]  AXI4L_MASTER0_WUSER;
wire          AXI4L_MASTER0_WVALID;
wire   [37:0] AXI4L_H264_ARADDR;
wire   [1:0]  AXI4L_H264_ARBURST;
wire   [3:0]  AXI4L_H264_ARCACHE;
wire   [8:0]  AXI4L_H264_ARID;
wire   [7:0]  AXI4L_H264_ARLEN;
wire   [1:0]  AXI4L_H264_ARLOCK;
wire   [2:0]  AXI4L_H264_ARPROT;
wire   [3:0]  AXI4L_H264_ARQOS;
wire          AXI4L_H264_SLAVE2_ARREADY;
wire   [3:0]  AXI4L_H264_ARREGION;
wire   [2:0]  AXI4L_H264_ARSIZE;
wire   [0:0]  AXI4L_H264_ARUSER;
wire          AXI4L_H264_ARVALID;
wire   [37:0] AXI4L_H264_AWADDR;
wire   [1:0]  AXI4L_H264_AWBURST;
wire   [3:0]  AXI4L_H264_AWCACHE;
wire   [8:0]  AXI4L_H264_AWID;
wire   [7:0]  AXI4L_H264_AWLEN;
wire   [1:0]  AXI4L_H264_AWLOCK;
wire   [2:0]  AXI4L_H264_AWPROT;
wire   [3:0]  AXI4L_H264_AWQOS;
wire          AXI4L_H264_SLAVE2_AWREADY;
wire   [3:0]  AXI4L_H264_AWREGION;
wire   [2:0]  AXI4L_H264_AWSIZE;
wire   [0:0]  AXI4L_H264_AWUSER;
wire          AXI4L_H264_AWVALID;
wire   [8:0]  AXI4L_H264_SLAVE2_BID;
wire          AXI4L_H264_BREADY;
wire   [1:0]  AXI4L_H264_SLAVE2_BRESP;
wire   [0:0]  AXI4L_H264_SLAVE2_BUSER;
wire          AXI4L_H264_SLAVE2_BVALID;
wire   [31:0] AXI4L_H264_SLAVE2_RDATA;
wire   [8:0]  AXI4L_H264_SLAVE2_RID;
wire          AXI4L_H264_SLAVE2_RLAST;
wire          AXI4L_H264_RREADY;
wire   [1:0]  AXI4L_H264_SLAVE2_RRESP;
wire   [0:0]  AXI4L_H264_SLAVE2_RUSER;
wire          AXI4L_H264_SLAVE2_RVALID;
wire   [31:0] AXI4L_H264_WDATA;
wire          AXI4L_H264_WLAST;
wire          AXI4L_H264_SLAVE2_WREADY;
wire   [3:0]  AXI4L_H264_WSTRB;
wire   [0:0]  AXI4L_H264_WUSER;
wire          AXI4L_H264_WVALID;
wire   [37:0] AXI4L_IE_ARADDR;
wire   [1:0]  AXI4L_IE_ARBURST;
wire   [3:0]  AXI4L_IE_ARCACHE;
wire   [8:0]  AXI4L_IE_ARID;
wire   [7:0]  AXI4L_IE_ARLEN;
wire   [1:0]  AXI4L_IE_ARLOCK;
wire   [2:0]  AXI4L_IE_ARPROT;
wire   [3:0]  AXI4L_IE_ARQOS;
wire          AXI4L_IE_SLAVE3_ARREADY;
wire   [3:0]  AXI4L_IE_ARREGION;
wire   [2:0]  AXI4L_IE_ARSIZE;
wire   [0:0]  AXI4L_IE_ARUSER;
wire          AXI4L_IE_ARVALID;
wire   [37:0] AXI4L_IE_AWADDR;
wire   [1:0]  AXI4L_IE_AWBURST;
wire   [3:0]  AXI4L_IE_AWCACHE;
wire   [8:0]  AXI4L_IE_AWID;
wire   [7:0]  AXI4L_IE_AWLEN;
wire   [1:0]  AXI4L_IE_AWLOCK;
wire   [2:0]  AXI4L_IE_AWPROT;
wire   [3:0]  AXI4L_IE_AWQOS;
wire          AXI4L_IE_SLAVE3_AWREADY;
wire   [3:0]  AXI4L_IE_AWREGION;
wire   [2:0]  AXI4L_IE_AWSIZE;
wire   [0:0]  AXI4L_IE_AWUSER;
wire          AXI4L_IE_AWVALID;
wire   [8:0]  AXI4L_IE_SLAVE3_BID;
wire          AXI4L_IE_BREADY;
wire   [1:0]  AXI4L_IE_SLAVE3_BRESP;
wire   [0:0]  AXI4L_IE_SLAVE3_BUSER;
wire          AXI4L_IE_SLAVE3_BVALID;
wire   [31:0] AXI4L_IE_SLAVE3_RDATA;
wire   [8:0]  AXI4L_IE_SLAVE3_RID;
wire          AXI4L_IE_SLAVE3_RLAST;
wire          AXI4L_IE_RREADY;
wire   [1:0]  AXI4L_IE_SLAVE3_RRESP;
wire   [0:0]  AXI4L_IE_SLAVE3_RUSER;
wire          AXI4L_IE_SLAVE3_RVALID;
wire   [31:0] AXI4L_IE_WDATA;
wire          AXI4L_IE_WLAST;
wire          AXI4L_IE_SLAVE3_WREADY;
wire   [3:0]  AXI4L_IE_WSTRB;
wire   [0:0]  AXI4L_IE_WUSER;
wire          AXI4L_IE_WVALID;
wire   [37:0] AXI4L_MIPI_ARADDR;
wire   [1:0]  AXI4L_MIPI_ARBURST;
wire   [3:0]  AXI4L_MIPI_ARCACHE;
wire   [8:0]  AXI4L_MIPI_ARID;
wire   [7:0]  AXI4L_MIPI_ARLEN;
wire   [1:0]  AXI4L_MIPI_ARLOCK;
wire   [2:0]  AXI4L_MIPI_ARPROT;
wire   [3:0]  AXI4L_MIPI_ARQOS;
wire          AXI4L_MIPI_SLAVE1_ARREADY;
wire   [3:0]  AXI4L_MIPI_ARREGION;
wire   [2:0]  AXI4L_MIPI_ARSIZE;
wire   [0:0]  AXI4L_MIPI_ARUSER;
wire          AXI4L_MIPI_ARVALID;
wire   [37:0] AXI4L_MIPI_AWADDR;
wire   [1:0]  AXI4L_MIPI_AWBURST;
wire   [3:0]  AXI4L_MIPI_AWCACHE;
wire   [8:0]  AXI4L_MIPI_AWID;
wire   [7:0]  AXI4L_MIPI_AWLEN;
wire   [1:0]  AXI4L_MIPI_AWLOCK;
wire   [2:0]  AXI4L_MIPI_AWPROT;
wire   [3:0]  AXI4L_MIPI_AWQOS;
wire          AXI4L_MIPI_SLAVE1_AWREADY;
wire   [3:0]  AXI4L_MIPI_AWREGION;
wire   [2:0]  AXI4L_MIPI_AWSIZE;
wire   [0:0]  AXI4L_MIPI_AWUSER;
wire          AXI4L_MIPI_AWVALID;
wire   [8:0]  AXI4L_MIPI_SLAVE1_BID;
wire          AXI4L_MIPI_BREADY;
wire   [1:0]  AXI4L_MIPI_SLAVE1_BRESP;
wire   [0:0]  AXI4L_MIPI_SLAVE1_BUSER;
wire          AXI4L_MIPI_SLAVE1_BVALID;
wire   [31:0] AXI4L_MIPI_SLAVE1_RDATA;
wire   [8:0]  AXI4L_MIPI_SLAVE1_RID;
wire          AXI4L_MIPI_SLAVE1_RLAST;
wire          AXI4L_MIPI_RREADY;
wire   [1:0]  AXI4L_MIPI_SLAVE1_RRESP;
wire   [0:0]  AXI4L_MIPI_SLAVE1_RUSER;
wire          AXI4L_MIPI_SLAVE1_RVALID;
wire   [31:0] AXI4L_MIPI_WDATA;
wire          AXI4L_MIPI_WLAST;
wire          AXI4L_MIPI_SLAVE1_WREADY;
wire   [3:0]  AXI4L_MIPI_WSTRB;
wire   [0:0]  AXI4L_MIPI_WUSER;
wire          AXI4L_MIPI_WVALID;
wire   [37:0] AXI4L_OSD_ARADDR;
wire   [1:0]  AXI4L_OSD_ARBURST;
wire   [3:0]  AXI4L_OSD_ARCACHE;
wire   [8:0]  AXI4L_OSD_ARID;
wire   [7:0]  AXI4L_OSD_ARLEN;
wire   [1:0]  AXI4L_OSD_ARLOCK;
wire   [2:0]  AXI4L_OSD_ARPROT;
wire   [3:0]  AXI4L_OSD_ARQOS;
wire          AXI4L_OSD_SLAVE5_ARREADY;
wire   [3:0]  AXI4L_OSD_ARREGION;
wire   [2:0]  AXI4L_OSD_ARSIZE;
wire   [0:0]  AXI4L_OSD_ARUSER;
wire          AXI4L_OSD_ARVALID;
wire   [37:0] AXI4L_OSD_AWADDR;
wire   [1:0]  AXI4L_OSD_AWBURST;
wire   [3:0]  AXI4L_OSD_AWCACHE;
wire   [8:0]  AXI4L_OSD_AWID;
wire   [7:0]  AXI4L_OSD_AWLEN;
wire   [1:0]  AXI4L_OSD_AWLOCK;
wire   [2:0]  AXI4L_OSD_AWPROT;
wire   [3:0]  AXI4L_OSD_AWQOS;
wire          AXI4L_OSD_SLAVE5_AWREADY;
wire   [3:0]  AXI4L_OSD_AWREGION;
wire   [2:0]  AXI4L_OSD_AWSIZE;
wire   [0:0]  AXI4L_OSD_AWUSER;
wire          AXI4L_OSD_AWVALID;
wire   [8:0]  AXI4L_OSD_SLAVE5_BID;
wire          AXI4L_OSD_BREADY;
wire   [1:0]  AXI4L_OSD_SLAVE5_BRESP;
wire   [0:0]  AXI4L_OSD_SLAVE5_BUSER;
wire          AXI4L_OSD_SLAVE5_BVALID;
wire   [63:0] AXI4L_OSD_SLAVE5_RDATA;
wire   [8:0]  AXI4L_OSD_SLAVE5_RID;
wire          AXI4L_OSD_SLAVE5_RLAST;
wire          AXI4L_OSD_RREADY;
wire   [1:0]  AXI4L_OSD_SLAVE5_RRESP;
wire   [0:0]  AXI4L_OSD_SLAVE5_RUSER;
wire          AXI4L_OSD_SLAVE5_RVALID;
wire   [63:0] AXI4L_OSD_WDATA;
wire          AXI4L_OSD_WLAST;
wire          AXI4L_OSD_SLAVE5_WREADY;
wire   [7:0]  AXI4L_OSD_WSTRB;
wire   [0:0]  AXI4L_OSD_WUSER;
wire          AXI4L_OSD_WVALID;
wire   [37:0] AXI4L_SCALER_ARADDR;
wire   [1:0]  AXI4L_SCALER_ARBURST;
wire   [3:0]  AXI4L_SCALER_ARCACHE;
wire   [8:0]  AXI4L_SCALER_ARID;
wire   [7:0]  AXI4L_SCALER_ARLEN;
wire   [1:0]  AXI4L_SCALER_ARLOCK;
wire   [2:0]  AXI4L_SCALER_ARPROT;
wire   [3:0]  AXI4L_SCALER_ARQOS;
wire          AXI4L_SCALER_SLAVE4_ARREADY;
wire   [3:0]  AXI4L_SCALER_ARREGION;
wire   [2:0]  AXI4L_SCALER_ARSIZE;
wire   [0:0]  AXI4L_SCALER_ARUSER;
wire          AXI4L_SCALER_ARVALID;
wire   [37:0] AXI4L_SCALER_AWADDR;
wire   [1:0]  AXI4L_SCALER_AWBURST;
wire   [3:0]  AXI4L_SCALER_AWCACHE;
wire   [8:0]  AXI4L_SCALER_AWID;
wire   [7:0]  AXI4L_SCALER_AWLEN;
wire   [1:0]  AXI4L_SCALER_AWLOCK;
wire   [2:0]  AXI4L_SCALER_AWPROT;
wire   [3:0]  AXI4L_SCALER_AWQOS;
wire          AXI4L_SCALER_SLAVE4_AWREADY;
wire   [3:0]  AXI4L_SCALER_AWREGION;
wire   [2:0]  AXI4L_SCALER_AWSIZE;
wire   [0:0]  AXI4L_SCALER_AWUSER;
wire          AXI4L_SCALER_AWVALID;
wire   [8:0]  AXI4L_SCALER_SLAVE4_BID;
wire          AXI4L_SCALER_BREADY;
wire   [1:0]  AXI4L_SCALER_SLAVE4_BRESP;
wire   [0:0]  AXI4L_SCALER_SLAVE4_BUSER;
wire          AXI4L_SCALER_SLAVE4_BVALID;
wire   [63:0] AXI4L_SCALER_SLAVE4_RDATA;
wire   [8:0]  AXI4L_SCALER_SLAVE4_RID;
wire          AXI4L_SCALER_SLAVE4_RLAST;
wire          AXI4L_SCALER_RREADY;
wire   [1:0]  AXI4L_SCALER_SLAVE4_RRESP;
wire   [0:0]  AXI4L_SCALER_SLAVE4_RUSER;
wire          AXI4L_SCALER_SLAVE4_RVALID;
wire   [63:0] AXI4L_SCALER_WDATA;
wire          AXI4L_SCALER_WLAST;
wire          AXI4L_SCALER_SLAVE4_WREADY;
wire   [7:0]  AXI4L_SCALER_WSTRB;
wire   [0:0]  AXI4L_SCALER_WUSER;
wire          AXI4L_SCALER_WVALID;
wire   [37:0] AXI4L_VDMA_ARADDR;
wire   [1:0]  AXI4L_VDMA_ARBURST;
wire   [3:0]  AXI4L_VDMA_ARCACHE;
wire   [8:0]  AXI4L_VDMA_ARID;
wire   [7:0]  AXI4L_VDMA_ARLEN;
wire   [1:0]  AXI4L_VDMA_ARLOCK;
wire   [2:0]  AXI4L_VDMA_ARPROT;
wire   [3:0]  AXI4L_VDMA_ARQOS;
wire          AXI4L_VDMA_SLAVE0_ARREADY;
wire   [3:0]  AXI4L_VDMA_ARREGION;
wire   [2:0]  AXI4L_VDMA_ARSIZE;
wire   [0:0]  AXI4L_VDMA_ARUSER;
wire          AXI4L_VDMA_ARVALID;
wire   [37:0] AXI4L_VDMA_AWADDR;
wire   [1:0]  AXI4L_VDMA_AWBURST;
wire   [3:0]  AXI4L_VDMA_AWCACHE;
wire   [8:0]  AXI4L_VDMA_AWID;
wire   [7:0]  AXI4L_VDMA_AWLEN;
wire   [1:0]  AXI4L_VDMA_AWLOCK;
wire   [2:0]  AXI4L_VDMA_AWPROT;
wire   [3:0]  AXI4L_VDMA_AWQOS;
wire          AXI4L_VDMA_SLAVE0_AWREADY;
wire   [3:0]  AXI4L_VDMA_AWREGION;
wire   [2:0]  AXI4L_VDMA_AWSIZE;
wire   [0:0]  AXI4L_VDMA_AWUSER;
wire          AXI4L_VDMA_AWVALID;
wire   [8:0]  AXI4L_VDMA_SLAVE0_BID;
wire          AXI4L_VDMA_BREADY;
wire   [1:0]  AXI4L_VDMA_SLAVE0_BRESP;
wire   [0:0]  AXI4L_VDMA_SLAVE0_BUSER;
wire          AXI4L_VDMA_SLAVE0_BVALID;
wire   [31:0] AXI4L_VDMA_SLAVE0_RDATA;
wire   [8:0]  AXI4L_VDMA_SLAVE0_RID;
wire          AXI4L_VDMA_SLAVE0_RLAST;
wire          AXI4L_VDMA_RREADY;
wire   [1:0]  AXI4L_VDMA_SLAVE0_RRESP;
wire   [0:0]  AXI4L_VDMA_SLAVE0_RUSER;
wire          AXI4L_VDMA_SLAVE0_RVALID;
wire   [31:0] AXI4L_VDMA_WDATA;
wire          AXI4L_VDMA_WLAST;
wire          AXI4L_VDMA_SLAVE0_WREADY;
wire   [3:0]  AXI4L_VDMA_WSTRB;
wire   [0:0]  AXI4L_VDMA_WUSER;
wire          AXI4L_VDMA_WVALID;
wire          AXI4L_H264_ARVALID_net_0;
wire          AXI4L_H264_AWVALID_net_0;
wire          AXI4L_H264_BREADY_net_0;
wire          AXI4L_H264_RREADY_net_0;
wire          AXI4L_H264_WLAST_net_0;
wire          AXI4L_H264_WVALID_net_0;
wire          AXI4L_IE_ARVALID_net_0;
wire          AXI4L_IE_AWVALID_net_0;
wire          AXI4L_IE_BREADY_net_0;
wire          AXI4L_IE_RREADY_net_0;
wire          AXI4L_IE_WLAST_net_0;
wire          AXI4L_IE_WVALID_net_0;
wire          AXI4L_ARREADY_net_0;
wire          AXI4L_AWREADY_net_0;
wire          AXI4L_BVALID_net_0;
wire          AXI4L_RLAST_net_0;
wire          AXI4L_RVALID_net_0;
wire          AXI4L_WREADY_net_0;
wire          AXI4L_MIPI_ARVALID_net_0;
wire          AXI4L_MIPI_AWVALID_net_0;
wire          AXI4L_MIPI_BREADY_net_0;
wire          AXI4L_MIPI_RREADY_net_0;
wire          AXI4L_MIPI_WLAST_net_0;
wire          AXI4L_MIPI_WVALID_net_0;
wire          AXI4L_OSD_ARVALID_net_0;
wire          AXI4L_OSD_AWVALID_net_0;
wire          AXI4L_OSD_BREADY_net_0;
wire          AXI4L_OSD_RREADY_net_0;
wire          AXI4L_OSD_WLAST_net_0;
wire          AXI4L_OSD_WVALID_net_0;
wire          AXI4L_SCALER_ARVALID_net_0;
wire          AXI4L_SCALER_AWVALID_net_0;
wire          AXI4L_SCALER_BREADY_net_0;
wire          AXI4L_SCALER_RREADY_net_0;
wire          AXI4L_SCALER_WLAST_net_0;
wire          AXI4L_SCALER_WVALID_net_0;
wire          AXI4L_VDMA_ARVALID_net_0;
wire          AXI4L_VDMA_AWVALID_net_0;
wire          AXI4L_VDMA_BREADY_net_0;
wire          AXI4L_VDMA_RREADY_net_0;
wire          AXI4L_VDMA_WLAST_net_0;
wire          AXI4L_VDMA_WVALID_net_0;
wire   [37:0] AXI4L_H264_ARADDR_net_0;
wire   [1:0]  AXI4L_H264_ARBURST_net_0;
wire   [3:0]  AXI4L_H264_ARCACHE_net_0;
wire   [8:0]  AXI4L_H264_ARID_net_0;
wire   [7:0]  AXI4L_H264_ARLEN_net_0;
wire   [1:0]  AXI4L_H264_ARLOCK_net_0;
wire   [2:0]  AXI4L_H264_ARPROT_net_0;
wire   [3:0]  AXI4L_H264_ARQOS_net_0;
wire   [3:0]  AXI4L_H264_ARREGION_net_0;
wire   [2:0]  AXI4L_H264_ARSIZE_net_0;
wire   [0:0]  AXI4L_H264_ARUSER_net_0;
wire   [37:0] AXI4L_H264_AWADDR_net_0;
wire   [1:0]  AXI4L_H264_AWBURST_net_0;
wire   [3:0]  AXI4L_H264_AWCACHE_net_0;
wire   [8:0]  AXI4L_H264_AWID_net_0;
wire   [7:0]  AXI4L_H264_AWLEN_net_0;
wire   [1:0]  AXI4L_H264_AWLOCK_net_0;
wire   [2:0]  AXI4L_H264_AWPROT_net_0;
wire   [3:0]  AXI4L_H264_AWQOS_net_0;
wire   [3:0]  AXI4L_H264_AWREGION_net_0;
wire   [2:0]  AXI4L_H264_AWSIZE_net_0;
wire   [0:0]  AXI4L_H264_AWUSER_net_0;
wire   [31:0] AXI4L_H264_WDATA_net_0;
wire   [3:0]  AXI4L_H264_WSTRB_net_0;
wire   [0:0]  AXI4L_H264_WUSER_net_0;
wire   [37:0] AXI4L_IE_ARADDR_net_0;
wire   [1:0]  AXI4L_IE_ARBURST_net_0;
wire   [3:0]  AXI4L_IE_ARCACHE_net_0;
wire   [8:0]  AXI4L_IE_ARID_net_0;
wire   [7:0]  AXI4L_IE_ARLEN_net_0;
wire   [1:0]  AXI4L_IE_ARLOCK_net_0;
wire   [2:0]  AXI4L_IE_ARPROT_net_0;
wire   [3:0]  AXI4L_IE_ARQOS_net_0;
wire   [3:0]  AXI4L_IE_ARREGION_net_0;
wire   [2:0]  AXI4L_IE_ARSIZE_net_0;
wire   [0:0]  AXI4L_IE_ARUSER_net_0;
wire   [37:0] AXI4L_IE_AWADDR_net_0;
wire   [1:0]  AXI4L_IE_AWBURST_net_0;
wire   [3:0]  AXI4L_IE_AWCACHE_net_0;
wire   [8:0]  AXI4L_IE_AWID_net_0;
wire   [7:0]  AXI4L_IE_AWLEN_net_0;
wire   [1:0]  AXI4L_IE_AWLOCK_net_0;
wire   [2:0]  AXI4L_IE_AWPROT_net_0;
wire   [3:0]  AXI4L_IE_AWQOS_net_0;
wire   [3:0]  AXI4L_IE_AWREGION_net_0;
wire   [2:0]  AXI4L_IE_AWSIZE_net_0;
wire   [0:0]  AXI4L_IE_AWUSER_net_0;
wire   [31:0] AXI4L_IE_WDATA_net_0;
wire   [3:0]  AXI4L_IE_WSTRB_net_0;
wire   [0:0]  AXI4L_IE_WUSER_net_0;
wire   [7:0]  AXI4L_BID_net_0;
wire   [1:0]  AXI4L_BRESP_net_0;
wire   [0:0]  AXI4L_BUSER_net_0;
wire   [63:0] AXI4L_RDATA_net_0;
wire   [7:0]  AXI4L_RID_net_0;
wire   [1:0]  AXI4L_RRESP_net_0;
wire   [0:0]  AXI4L_RUSER_net_0;
wire   [37:0] AXI4L_MIPI_ARADDR_net_0;
wire   [1:0]  AXI4L_MIPI_ARBURST_net_0;
wire   [3:0]  AXI4L_MIPI_ARCACHE_net_0;
wire   [8:0]  AXI4L_MIPI_ARID_net_0;
wire   [7:0]  AXI4L_MIPI_ARLEN_net_0;
wire   [1:0]  AXI4L_MIPI_ARLOCK_net_0;
wire   [2:0]  AXI4L_MIPI_ARPROT_net_0;
wire   [3:0]  AXI4L_MIPI_ARQOS_net_0;
wire   [3:0]  AXI4L_MIPI_ARREGION_net_0;
wire   [2:0]  AXI4L_MIPI_ARSIZE_net_0;
wire   [0:0]  AXI4L_MIPI_ARUSER_net_0;
wire   [37:0] AXI4L_MIPI_AWADDR_net_0;
wire   [1:0]  AXI4L_MIPI_AWBURST_net_0;
wire   [3:0]  AXI4L_MIPI_AWCACHE_net_0;
wire   [8:0]  AXI4L_MIPI_AWID_net_0;
wire   [7:0]  AXI4L_MIPI_AWLEN_net_0;
wire   [1:0]  AXI4L_MIPI_AWLOCK_net_0;
wire   [2:0]  AXI4L_MIPI_AWPROT_net_0;
wire   [3:0]  AXI4L_MIPI_AWQOS_net_0;
wire   [3:0]  AXI4L_MIPI_AWREGION_net_0;
wire   [2:0]  AXI4L_MIPI_AWSIZE_net_0;
wire   [0:0]  AXI4L_MIPI_AWUSER_net_0;
wire   [31:0] AXI4L_MIPI_WDATA_net_0;
wire   [3:0]  AXI4L_MIPI_WSTRB_net_0;
wire   [0:0]  AXI4L_MIPI_WUSER_net_0;
wire   [37:0] AXI4L_OSD_ARADDR_net_0;
wire   [1:0]  AXI4L_OSD_ARBURST_net_0;
wire   [3:0]  AXI4L_OSD_ARCACHE_net_0;
wire   [8:0]  AXI4L_OSD_ARID_net_0;
wire   [7:0]  AXI4L_OSD_ARLEN_net_0;
wire   [1:0]  AXI4L_OSD_ARLOCK_net_0;
wire   [2:0]  AXI4L_OSD_ARPROT_net_0;
wire   [3:0]  AXI4L_OSD_ARQOS_net_0;
wire   [3:0]  AXI4L_OSD_ARREGION_net_0;
wire   [2:0]  AXI4L_OSD_ARSIZE_net_0;
wire   [0:0]  AXI4L_OSD_ARUSER_net_0;
wire   [37:0] AXI4L_OSD_AWADDR_net_0;
wire   [1:0]  AXI4L_OSD_AWBURST_net_0;
wire   [3:0]  AXI4L_OSD_AWCACHE_net_0;
wire   [8:0]  AXI4L_OSD_AWID_net_0;
wire   [7:0]  AXI4L_OSD_AWLEN_net_0;
wire   [1:0]  AXI4L_OSD_AWLOCK_net_0;
wire   [2:0]  AXI4L_OSD_AWPROT_net_0;
wire   [3:0]  AXI4L_OSD_AWQOS_net_0;
wire   [3:0]  AXI4L_OSD_AWREGION_net_0;
wire   [2:0]  AXI4L_OSD_AWSIZE_net_0;
wire   [0:0]  AXI4L_OSD_AWUSER_net_0;
wire   [63:0] AXI4L_OSD_WDATA_net_0;
wire   [7:0]  AXI4L_OSD_WSTRB_net_0;
wire   [0:0]  AXI4L_OSD_WUSER_net_0;
wire   [37:0] AXI4L_SCALER_ARADDR_net_0;
wire   [1:0]  AXI4L_SCALER_ARBURST_net_0;
wire   [3:0]  AXI4L_SCALER_ARCACHE_net_0;
wire   [8:0]  AXI4L_SCALER_ARID_net_0;
wire   [7:0]  AXI4L_SCALER_ARLEN_net_0;
wire   [1:0]  AXI4L_SCALER_ARLOCK_net_0;
wire   [2:0]  AXI4L_SCALER_ARPROT_net_0;
wire   [3:0]  AXI4L_SCALER_ARQOS_net_0;
wire   [3:0]  AXI4L_SCALER_ARREGION_net_0;
wire   [2:0]  AXI4L_SCALER_ARSIZE_net_0;
wire   [0:0]  AXI4L_SCALER_ARUSER_net_0;
wire   [37:0] AXI4L_SCALER_AWADDR_net_0;
wire   [1:0]  AXI4L_SCALER_AWBURST_net_0;
wire   [3:0]  AXI4L_SCALER_AWCACHE_net_0;
wire   [8:0]  AXI4L_SCALER_AWID_net_0;
wire   [7:0]  AXI4L_SCALER_AWLEN_net_0;
wire   [1:0]  AXI4L_SCALER_AWLOCK_net_0;
wire   [2:0]  AXI4L_SCALER_AWPROT_net_0;
wire   [3:0]  AXI4L_SCALER_AWQOS_net_0;
wire   [3:0]  AXI4L_SCALER_AWREGION_net_0;
wire   [2:0]  AXI4L_SCALER_AWSIZE_net_0;
wire   [0:0]  AXI4L_SCALER_AWUSER_net_0;
wire   [63:0] AXI4L_SCALER_WDATA_net_0;
wire   [7:0]  AXI4L_SCALER_WSTRB_net_0;
wire   [0:0]  AXI4L_SCALER_WUSER_net_0;
wire   [37:0] AXI4L_VDMA_ARADDR_net_0;
wire   [1:0]  AXI4L_VDMA_ARBURST_net_0;
wire   [3:0]  AXI4L_VDMA_ARCACHE_net_0;
wire   [8:0]  AXI4L_VDMA_ARID_net_0;
wire   [7:0]  AXI4L_VDMA_ARLEN_net_0;
wire   [1:0]  AXI4L_VDMA_ARLOCK_net_0;
wire   [2:0]  AXI4L_VDMA_ARPROT_net_0;
wire   [3:0]  AXI4L_VDMA_ARQOS_net_0;
wire   [3:0]  AXI4L_VDMA_ARREGION_net_0;
wire   [2:0]  AXI4L_VDMA_ARSIZE_net_0;
wire   [0:0]  AXI4L_VDMA_ARUSER_net_0;
wire   [37:0] AXI4L_VDMA_AWADDR_net_0;
wire   [1:0]  AXI4L_VDMA_AWBURST_net_0;
wire   [3:0]  AXI4L_VDMA_AWCACHE_net_0;
wire   [8:0]  AXI4L_VDMA_AWID_net_0;
wire   [7:0]  AXI4L_VDMA_AWLEN_net_0;
wire   [1:0]  AXI4L_VDMA_AWLOCK_net_0;
wire   [2:0]  AXI4L_VDMA_AWPROT_net_0;
wire   [3:0]  AXI4L_VDMA_AWQOS_net_0;
wire   [3:0]  AXI4L_VDMA_AWREGION_net_0;
wire   [2:0]  AXI4L_VDMA_AWSIZE_net_0;
wire   [0:0]  AXI4L_VDMA_AWUSER_net_0;
wire   [31:0] AXI4L_VDMA_WDATA_net_0;
wire   [3:0]  AXI4L_VDMA_WSTRB_net_0;
wire   [0:0]  AXI4L_VDMA_WUSER_net_0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign AXI4L_H264_ARVALID_net_0          = AXI4L_H264_ARVALID;
assign AXI4L_H264_SLAVE2_ARVALID         = AXI4L_H264_ARVALID_net_0;
assign AXI4L_H264_AWVALID_net_0          = AXI4L_H264_AWVALID;
assign AXI4L_H264_SLAVE2_AWVALID         = AXI4L_H264_AWVALID_net_0;
assign AXI4L_H264_BREADY_net_0           = AXI4L_H264_BREADY;
assign AXI4L_H264_SLAVE2_BREADY          = AXI4L_H264_BREADY_net_0;
assign AXI4L_H264_RREADY_net_0           = AXI4L_H264_RREADY;
assign AXI4L_H264_SLAVE2_RREADY          = AXI4L_H264_RREADY_net_0;
assign AXI4L_H264_WLAST_net_0            = AXI4L_H264_WLAST;
assign AXI4L_H264_SLAVE2_WLAST           = AXI4L_H264_WLAST_net_0;
assign AXI4L_H264_WVALID_net_0           = AXI4L_H264_WVALID;
assign AXI4L_H264_SLAVE2_WVALID          = AXI4L_H264_WVALID_net_0;
assign AXI4L_IE_ARVALID_net_0            = AXI4L_IE_ARVALID;
assign AXI4L_IE_SLAVE3_ARVALID           = AXI4L_IE_ARVALID_net_0;
assign AXI4L_IE_AWVALID_net_0            = AXI4L_IE_AWVALID;
assign AXI4L_IE_SLAVE3_AWVALID           = AXI4L_IE_AWVALID_net_0;
assign AXI4L_IE_BREADY_net_0             = AXI4L_IE_BREADY;
assign AXI4L_IE_SLAVE3_BREADY            = AXI4L_IE_BREADY_net_0;
assign AXI4L_IE_RREADY_net_0             = AXI4L_IE_RREADY;
assign AXI4L_IE_SLAVE3_RREADY            = AXI4L_IE_RREADY_net_0;
assign AXI4L_IE_WLAST_net_0              = AXI4L_IE_WLAST;
assign AXI4L_IE_SLAVE3_WLAST             = AXI4L_IE_WLAST_net_0;
assign AXI4L_IE_WVALID_net_0             = AXI4L_IE_WVALID;
assign AXI4L_IE_SLAVE3_WVALID            = AXI4L_IE_WVALID_net_0;
assign AXI4L_ARREADY_net_0               = AXI4L_ARREADY;
assign AXI4L_MASTER0_ARREADY             = AXI4L_ARREADY_net_0;
assign AXI4L_AWREADY_net_0               = AXI4L_AWREADY;
assign AXI4L_MASTER0_AWREADY             = AXI4L_AWREADY_net_0;
assign AXI4L_BVALID_net_0                = AXI4L_BVALID;
assign AXI4L_MASTER0_BVALID              = AXI4L_BVALID_net_0;
assign AXI4L_RLAST_net_0                 = AXI4L_RLAST;
assign AXI4L_MASTER0_RLAST               = AXI4L_RLAST_net_0;
assign AXI4L_RVALID_net_0                = AXI4L_RVALID;
assign AXI4L_MASTER0_RVALID              = AXI4L_RVALID_net_0;
assign AXI4L_WREADY_net_0                = AXI4L_WREADY;
assign AXI4L_MASTER0_WREADY              = AXI4L_WREADY_net_0;
assign AXI4L_MIPI_ARVALID_net_0          = AXI4L_MIPI_ARVALID;
assign AXI4L_MIPI_SLAVE1_ARVALID         = AXI4L_MIPI_ARVALID_net_0;
assign AXI4L_MIPI_AWVALID_net_0          = AXI4L_MIPI_AWVALID;
assign AXI4L_MIPI_SLAVE1_AWVALID         = AXI4L_MIPI_AWVALID_net_0;
assign AXI4L_MIPI_BREADY_net_0           = AXI4L_MIPI_BREADY;
assign AXI4L_MIPI_SLAVE1_BREADY          = AXI4L_MIPI_BREADY_net_0;
assign AXI4L_MIPI_RREADY_net_0           = AXI4L_MIPI_RREADY;
assign AXI4L_MIPI_SLAVE1_RREADY          = AXI4L_MIPI_RREADY_net_0;
assign AXI4L_MIPI_WLAST_net_0            = AXI4L_MIPI_WLAST;
assign AXI4L_MIPI_SLAVE1_WLAST           = AXI4L_MIPI_WLAST_net_0;
assign AXI4L_MIPI_WVALID_net_0           = AXI4L_MIPI_WVALID;
assign AXI4L_MIPI_SLAVE1_WVALID          = AXI4L_MIPI_WVALID_net_0;
assign AXI4L_OSD_ARVALID_net_0           = AXI4L_OSD_ARVALID;
assign AXI4L_OSD_SLAVE5_ARVALID          = AXI4L_OSD_ARVALID_net_0;
assign AXI4L_OSD_AWVALID_net_0           = AXI4L_OSD_AWVALID;
assign AXI4L_OSD_SLAVE5_AWVALID          = AXI4L_OSD_AWVALID_net_0;
assign AXI4L_OSD_BREADY_net_0            = AXI4L_OSD_BREADY;
assign AXI4L_OSD_SLAVE5_BREADY           = AXI4L_OSD_BREADY_net_0;
assign AXI4L_OSD_RREADY_net_0            = AXI4L_OSD_RREADY;
assign AXI4L_OSD_SLAVE5_RREADY           = AXI4L_OSD_RREADY_net_0;
assign AXI4L_OSD_WLAST_net_0             = AXI4L_OSD_WLAST;
assign AXI4L_OSD_SLAVE5_WLAST            = AXI4L_OSD_WLAST_net_0;
assign AXI4L_OSD_WVALID_net_0            = AXI4L_OSD_WVALID;
assign AXI4L_OSD_SLAVE5_WVALID           = AXI4L_OSD_WVALID_net_0;
assign AXI4L_SCALER_ARVALID_net_0        = AXI4L_SCALER_ARVALID;
assign AXI4L_SCALER_SLAVE4_ARVALID       = AXI4L_SCALER_ARVALID_net_0;
assign AXI4L_SCALER_AWVALID_net_0        = AXI4L_SCALER_AWVALID;
assign AXI4L_SCALER_SLAVE4_AWVALID       = AXI4L_SCALER_AWVALID_net_0;
assign AXI4L_SCALER_BREADY_net_0         = AXI4L_SCALER_BREADY;
assign AXI4L_SCALER_SLAVE4_BREADY        = AXI4L_SCALER_BREADY_net_0;
assign AXI4L_SCALER_RREADY_net_0         = AXI4L_SCALER_RREADY;
assign AXI4L_SCALER_SLAVE4_RREADY        = AXI4L_SCALER_RREADY_net_0;
assign AXI4L_SCALER_WLAST_net_0          = AXI4L_SCALER_WLAST;
assign AXI4L_SCALER_SLAVE4_WLAST         = AXI4L_SCALER_WLAST_net_0;
assign AXI4L_SCALER_WVALID_net_0         = AXI4L_SCALER_WVALID;
assign AXI4L_SCALER_SLAVE4_WVALID        = AXI4L_SCALER_WVALID_net_0;
assign AXI4L_VDMA_ARVALID_net_0          = AXI4L_VDMA_ARVALID;
assign AXI4L_VDMA_SLAVE0_ARVALID         = AXI4L_VDMA_ARVALID_net_0;
assign AXI4L_VDMA_AWVALID_net_0          = AXI4L_VDMA_AWVALID;
assign AXI4L_VDMA_SLAVE0_AWVALID         = AXI4L_VDMA_AWVALID_net_0;
assign AXI4L_VDMA_BREADY_net_0           = AXI4L_VDMA_BREADY;
assign AXI4L_VDMA_SLAVE0_BREADY          = AXI4L_VDMA_BREADY_net_0;
assign AXI4L_VDMA_RREADY_net_0           = AXI4L_VDMA_RREADY;
assign AXI4L_VDMA_SLAVE0_RREADY          = AXI4L_VDMA_RREADY_net_0;
assign AXI4L_VDMA_WLAST_net_0            = AXI4L_VDMA_WLAST;
assign AXI4L_VDMA_SLAVE0_WLAST           = AXI4L_VDMA_WLAST_net_0;
assign AXI4L_VDMA_WVALID_net_0           = AXI4L_VDMA_WVALID;
assign AXI4L_VDMA_SLAVE0_WVALID          = AXI4L_VDMA_WVALID_net_0;
assign AXI4L_H264_ARADDR_net_0           = AXI4L_H264_ARADDR;
assign AXI4L_H264_SLAVE2_ARADDR[37:0]    = AXI4L_H264_ARADDR_net_0;
assign AXI4L_H264_ARBURST_net_0          = AXI4L_H264_ARBURST;
assign AXI4L_H264_SLAVE2_ARBURST[1:0]    = AXI4L_H264_ARBURST_net_0;
assign AXI4L_H264_ARCACHE_net_0          = AXI4L_H264_ARCACHE;
assign AXI4L_H264_SLAVE2_ARCACHE[3:0]    = AXI4L_H264_ARCACHE_net_0;
assign AXI4L_H264_ARID_net_0             = AXI4L_H264_ARID;
assign AXI4L_H264_SLAVE2_ARID[8:0]       = AXI4L_H264_ARID_net_0;
assign AXI4L_H264_ARLEN_net_0            = AXI4L_H264_ARLEN;
assign AXI4L_H264_SLAVE2_ARLEN[7:0]      = AXI4L_H264_ARLEN_net_0;
assign AXI4L_H264_ARLOCK_net_0           = AXI4L_H264_ARLOCK;
assign AXI4L_H264_SLAVE2_ARLOCK[1:0]     = AXI4L_H264_ARLOCK_net_0;
assign AXI4L_H264_ARPROT_net_0           = AXI4L_H264_ARPROT;
assign AXI4L_H264_SLAVE2_ARPROT[2:0]     = AXI4L_H264_ARPROT_net_0;
assign AXI4L_H264_ARQOS_net_0            = AXI4L_H264_ARQOS;
assign AXI4L_H264_SLAVE2_ARQOS[3:0]      = AXI4L_H264_ARQOS_net_0;
assign AXI4L_H264_ARREGION_net_0         = AXI4L_H264_ARREGION;
assign AXI4L_H264_SLAVE2_ARREGION[3:0]   = AXI4L_H264_ARREGION_net_0;
assign AXI4L_H264_ARSIZE_net_0           = AXI4L_H264_ARSIZE;
assign AXI4L_H264_SLAVE2_ARSIZE[2:0]     = AXI4L_H264_ARSIZE_net_0;
assign AXI4L_H264_ARUSER_net_0[0]        = AXI4L_H264_ARUSER[0];
assign AXI4L_H264_SLAVE2_ARUSER[0:0]     = AXI4L_H264_ARUSER_net_0[0];
assign AXI4L_H264_AWADDR_net_0           = AXI4L_H264_AWADDR;
assign AXI4L_H264_SLAVE2_AWADDR[37:0]    = AXI4L_H264_AWADDR_net_0;
assign AXI4L_H264_AWBURST_net_0          = AXI4L_H264_AWBURST;
assign AXI4L_H264_SLAVE2_AWBURST[1:0]    = AXI4L_H264_AWBURST_net_0;
assign AXI4L_H264_AWCACHE_net_0          = AXI4L_H264_AWCACHE;
assign AXI4L_H264_SLAVE2_AWCACHE[3:0]    = AXI4L_H264_AWCACHE_net_0;
assign AXI4L_H264_AWID_net_0             = AXI4L_H264_AWID;
assign AXI4L_H264_SLAVE2_AWID[8:0]       = AXI4L_H264_AWID_net_0;
assign AXI4L_H264_AWLEN_net_0            = AXI4L_H264_AWLEN;
assign AXI4L_H264_SLAVE2_AWLEN[7:0]      = AXI4L_H264_AWLEN_net_0;
assign AXI4L_H264_AWLOCK_net_0           = AXI4L_H264_AWLOCK;
assign AXI4L_H264_SLAVE2_AWLOCK[1:0]     = AXI4L_H264_AWLOCK_net_0;
assign AXI4L_H264_AWPROT_net_0           = AXI4L_H264_AWPROT;
assign AXI4L_H264_SLAVE2_AWPROT[2:0]     = AXI4L_H264_AWPROT_net_0;
assign AXI4L_H264_AWQOS_net_0            = AXI4L_H264_AWQOS;
assign AXI4L_H264_SLAVE2_AWQOS[3:0]      = AXI4L_H264_AWQOS_net_0;
assign AXI4L_H264_AWREGION_net_0         = AXI4L_H264_AWREGION;
assign AXI4L_H264_SLAVE2_AWREGION[3:0]   = AXI4L_H264_AWREGION_net_0;
assign AXI4L_H264_AWSIZE_net_0           = AXI4L_H264_AWSIZE;
assign AXI4L_H264_SLAVE2_AWSIZE[2:0]     = AXI4L_H264_AWSIZE_net_0;
assign AXI4L_H264_AWUSER_net_0[0]        = AXI4L_H264_AWUSER[0];
assign AXI4L_H264_SLAVE2_AWUSER[0:0]     = AXI4L_H264_AWUSER_net_0[0];
assign AXI4L_H264_WDATA_net_0            = AXI4L_H264_WDATA;
assign AXI4L_H264_SLAVE2_WDATA[31:0]     = AXI4L_H264_WDATA_net_0;
assign AXI4L_H264_WSTRB_net_0            = AXI4L_H264_WSTRB;
assign AXI4L_H264_SLAVE2_WSTRB[3:0]      = AXI4L_H264_WSTRB_net_0;
assign AXI4L_H264_WUSER_net_0[0]         = AXI4L_H264_WUSER[0];
assign AXI4L_H264_SLAVE2_WUSER[0:0]      = AXI4L_H264_WUSER_net_0[0];
assign AXI4L_IE_ARADDR_net_0             = AXI4L_IE_ARADDR;
assign AXI4L_IE_SLAVE3_ARADDR[37:0]      = AXI4L_IE_ARADDR_net_0;
assign AXI4L_IE_ARBURST_net_0            = AXI4L_IE_ARBURST;
assign AXI4L_IE_SLAVE3_ARBURST[1:0]      = AXI4L_IE_ARBURST_net_0;
assign AXI4L_IE_ARCACHE_net_0            = AXI4L_IE_ARCACHE;
assign AXI4L_IE_SLAVE3_ARCACHE[3:0]      = AXI4L_IE_ARCACHE_net_0;
assign AXI4L_IE_ARID_net_0               = AXI4L_IE_ARID;
assign AXI4L_IE_SLAVE3_ARID[8:0]         = AXI4L_IE_ARID_net_0;
assign AXI4L_IE_ARLEN_net_0              = AXI4L_IE_ARLEN;
assign AXI4L_IE_SLAVE3_ARLEN[7:0]        = AXI4L_IE_ARLEN_net_0;
assign AXI4L_IE_ARLOCK_net_0             = AXI4L_IE_ARLOCK;
assign AXI4L_IE_SLAVE3_ARLOCK[1:0]       = AXI4L_IE_ARLOCK_net_0;
assign AXI4L_IE_ARPROT_net_0             = AXI4L_IE_ARPROT;
assign AXI4L_IE_SLAVE3_ARPROT[2:0]       = AXI4L_IE_ARPROT_net_0;
assign AXI4L_IE_ARQOS_net_0              = AXI4L_IE_ARQOS;
assign AXI4L_IE_SLAVE3_ARQOS[3:0]        = AXI4L_IE_ARQOS_net_0;
assign AXI4L_IE_ARREGION_net_0           = AXI4L_IE_ARREGION;
assign AXI4L_IE_SLAVE3_ARREGION[3:0]     = AXI4L_IE_ARREGION_net_0;
assign AXI4L_IE_ARSIZE_net_0             = AXI4L_IE_ARSIZE;
assign AXI4L_IE_SLAVE3_ARSIZE[2:0]       = AXI4L_IE_ARSIZE_net_0;
assign AXI4L_IE_ARUSER_net_0[0]          = AXI4L_IE_ARUSER[0];
assign AXI4L_IE_SLAVE3_ARUSER[0:0]       = AXI4L_IE_ARUSER_net_0[0];
assign AXI4L_IE_AWADDR_net_0             = AXI4L_IE_AWADDR;
assign AXI4L_IE_SLAVE3_AWADDR[37:0]      = AXI4L_IE_AWADDR_net_0;
assign AXI4L_IE_AWBURST_net_0            = AXI4L_IE_AWBURST;
assign AXI4L_IE_SLAVE3_AWBURST[1:0]      = AXI4L_IE_AWBURST_net_0;
assign AXI4L_IE_AWCACHE_net_0            = AXI4L_IE_AWCACHE;
assign AXI4L_IE_SLAVE3_AWCACHE[3:0]      = AXI4L_IE_AWCACHE_net_0;
assign AXI4L_IE_AWID_net_0               = AXI4L_IE_AWID;
assign AXI4L_IE_SLAVE3_AWID[8:0]         = AXI4L_IE_AWID_net_0;
assign AXI4L_IE_AWLEN_net_0              = AXI4L_IE_AWLEN;
assign AXI4L_IE_SLAVE3_AWLEN[7:0]        = AXI4L_IE_AWLEN_net_0;
assign AXI4L_IE_AWLOCK_net_0             = AXI4L_IE_AWLOCK;
assign AXI4L_IE_SLAVE3_AWLOCK[1:0]       = AXI4L_IE_AWLOCK_net_0;
assign AXI4L_IE_AWPROT_net_0             = AXI4L_IE_AWPROT;
assign AXI4L_IE_SLAVE3_AWPROT[2:0]       = AXI4L_IE_AWPROT_net_0;
assign AXI4L_IE_AWQOS_net_0              = AXI4L_IE_AWQOS;
assign AXI4L_IE_SLAVE3_AWQOS[3:0]        = AXI4L_IE_AWQOS_net_0;
assign AXI4L_IE_AWREGION_net_0           = AXI4L_IE_AWREGION;
assign AXI4L_IE_SLAVE3_AWREGION[3:0]     = AXI4L_IE_AWREGION_net_0;
assign AXI4L_IE_AWSIZE_net_0             = AXI4L_IE_AWSIZE;
assign AXI4L_IE_SLAVE3_AWSIZE[2:0]       = AXI4L_IE_AWSIZE_net_0;
assign AXI4L_IE_AWUSER_net_0[0]          = AXI4L_IE_AWUSER[0];
assign AXI4L_IE_SLAVE3_AWUSER[0:0]       = AXI4L_IE_AWUSER_net_0[0];
assign AXI4L_IE_WDATA_net_0              = AXI4L_IE_WDATA;
assign AXI4L_IE_SLAVE3_WDATA[31:0]       = AXI4L_IE_WDATA_net_0;
assign AXI4L_IE_WSTRB_net_0              = AXI4L_IE_WSTRB;
assign AXI4L_IE_SLAVE3_WSTRB[3:0]        = AXI4L_IE_WSTRB_net_0;
assign AXI4L_IE_WUSER_net_0[0]           = AXI4L_IE_WUSER[0];
assign AXI4L_IE_SLAVE3_WUSER[0:0]        = AXI4L_IE_WUSER_net_0[0];
assign AXI4L_BID_net_0                   = AXI4L_BID;
assign AXI4L_MASTER0_BID[7:0]            = AXI4L_BID_net_0;
assign AXI4L_BRESP_net_0                 = AXI4L_BRESP;
assign AXI4L_MASTER0_BRESP[1:0]          = AXI4L_BRESP_net_0;
assign AXI4L_BUSER_net_0[0]              = AXI4L_BUSER[0];
assign AXI4L_MASTER0_BUSER[0:0]          = AXI4L_BUSER_net_0[0];
assign AXI4L_RDATA_net_0                 = AXI4L_RDATA;
assign AXI4L_MASTER0_RDATA[63:0]         = AXI4L_RDATA_net_0;
assign AXI4L_RID_net_0                   = AXI4L_RID;
assign AXI4L_MASTER0_RID[7:0]            = AXI4L_RID_net_0;
assign AXI4L_RRESP_net_0                 = AXI4L_RRESP;
assign AXI4L_MASTER0_RRESP[1:0]          = AXI4L_RRESP_net_0;
assign AXI4L_RUSER_net_0[0]              = AXI4L_RUSER[0];
assign AXI4L_MASTER0_RUSER[0:0]          = AXI4L_RUSER_net_0[0];
assign AXI4L_MIPI_ARADDR_net_0           = AXI4L_MIPI_ARADDR;
assign AXI4L_MIPI_SLAVE1_ARADDR[37:0]    = AXI4L_MIPI_ARADDR_net_0;
assign AXI4L_MIPI_ARBURST_net_0          = AXI4L_MIPI_ARBURST;
assign AXI4L_MIPI_SLAVE1_ARBURST[1:0]    = AXI4L_MIPI_ARBURST_net_0;
assign AXI4L_MIPI_ARCACHE_net_0          = AXI4L_MIPI_ARCACHE;
assign AXI4L_MIPI_SLAVE1_ARCACHE[3:0]    = AXI4L_MIPI_ARCACHE_net_0;
assign AXI4L_MIPI_ARID_net_0             = AXI4L_MIPI_ARID;
assign AXI4L_MIPI_SLAVE1_ARID[8:0]       = AXI4L_MIPI_ARID_net_0;
assign AXI4L_MIPI_ARLEN_net_0            = AXI4L_MIPI_ARLEN;
assign AXI4L_MIPI_SLAVE1_ARLEN[7:0]      = AXI4L_MIPI_ARLEN_net_0;
assign AXI4L_MIPI_ARLOCK_net_0           = AXI4L_MIPI_ARLOCK;
assign AXI4L_MIPI_SLAVE1_ARLOCK[1:0]     = AXI4L_MIPI_ARLOCK_net_0;
assign AXI4L_MIPI_ARPROT_net_0           = AXI4L_MIPI_ARPROT;
assign AXI4L_MIPI_SLAVE1_ARPROT[2:0]     = AXI4L_MIPI_ARPROT_net_0;
assign AXI4L_MIPI_ARQOS_net_0            = AXI4L_MIPI_ARQOS;
assign AXI4L_MIPI_SLAVE1_ARQOS[3:0]      = AXI4L_MIPI_ARQOS_net_0;
assign AXI4L_MIPI_ARREGION_net_0         = AXI4L_MIPI_ARREGION;
assign AXI4L_MIPI_SLAVE1_ARREGION[3:0]   = AXI4L_MIPI_ARREGION_net_0;
assign AXI4L_MIPI_ARSIZE_net_0           = AXI4L_MIPI_ARSIZE;
assign AXI4L_MIPI_SLAVE1_ARSIZE[2:0]     = AXI4L_MIPI_ARSIZE_net_0;
assign AXI4L_MIPI_ARUSER_net_0[0]        = AXI4L_MIPI_ARUSER[0];
assign AXI4L_MIPI_SLAVE1_ARUSER[0:0]     = AXI4L_MIPI_ARUSER_net_0[0];
assign AXI4L_MIPI_AWADDR_net_0           = AXI4L_MIPI_AWADDR;
assign AXI4L_MIPI_SLAVE1_AWADDR[37:0]    = AXI4L_MIPI_AWADDR_net_0;
assign AXI4L_MIPI_AWBURST_net_0          = AXI4L_MIPI_AWBURST;
assign AXI4L_MIPI_SLAVE1_AWBURST[1:0]    = AXI4L_MIPI_AWBURST_net_0;
assign AXI4L_MIPI_AWCACHE_net_0          = AXI4L_MIPI_AWCACHE;
assign AXI4L_MIPI_SLAVE1_AWCACHE[3:0]    = AXI4L_MIPI_AWCACHE_net_0;
assign AXI4L_MIPI_AWID_net_0             = AXI4L_MIPI_AWID;
assign AXI4L_MIPI_SLAVE1_AWID[8:0]       = AXI4L_MIPI_AWID_net_0;
assign AXI4L_MIPI_AWLEN_net_0            = AXI4L_MIPI_AWLEN;
assign AXI4L_MIPI_SLAVE1_AWLEN[7:0]      = AXI4L_MIPI_AWLEN_net_0;
assign AXI4L_MIPI_AWLOCK_net_0           = AXI4L_MIPI_AWLOCK;
assign AXI4L_MIPI_SLAVE1_AWLOCK[1:0]     = AXI4L_MIPI_AWLOCK_net_0;
assign AXI4L_MIPI_AWPROT_net_0           = AXI4L_MIPI_AWPROT;
assign AXI4L_MIPI_SLAVE1_AWPROT[2:0]     = AXI4L_MIPI_AWPROT_net_0;
assign AXI4L_MIPI_AWQOS_net_0            = AXI4L_MIPI_AWQOS;
assign AXI4L_MIPI_SLAVE1_AWQOS[3:0]      = AXI4L_MIPI_AWQOS_net_0;
assign AXI4L_MIPI_AWREGION_net_0         = AXI4L_MIPI_AWREGION;
assign AXI4L_MIPI_SLAVE1_AWREGION[3:0]   = AXI4L_MIPI_AWREGION_net_0;
assign AXI4L_MIPI_AWSIZE_net_0           = AXI4L_MIPI_AWSIZE;
assign AXI4L_MIPI_SLAVE1_AWSIZE[2:0]     = AXI4L_MIPI_AWSIZE_net_0;
assign AXI4L_MIPI_AWUSER_net_0[0]        = AXI4L_MIPI_AWUSER[0];
assign AXI4L_MIPI_SLAVE1_AWUSER[0:0]     = AXI4L_MIPI_AWUSER_net_0[0];
assign AXI4L_MIPI_WDATA_net_0            = AXI4L_MIPI_WDATA;
assign AXI4L_MIPI_SLAVE1_WDATA[31:0]     = AXI4L_MIPI_WDATA_net_0;
assign AXI4L_MIPI_WSTRB_net_0            = AXI4L_MIPI_WSTRB;
assign AXI4L_MIPI_SLAVE1_WSTRB[3:0]      = AXI4L_MIPI_WSTRB_net_0;
assign AXI4L_MIPI_WUSER_net_0[0]         = AXI4L_MIPI_WUSER[0];
assign AXI4L_MIPI_SLAVE1_WUSER[0:0]      = AXI4L_MIPI_WUSER_net_0[0];
assign AXI4L_OSD_ARADDR_net_0            = AXI4L_OSD_ARADDR;
assign AXI4L_OSD_SLAVE5_ARADDR[37:0]     = AXI4L_OSD_ARADDR_net_0;
assign AXI4L_OSD_ARBURST_net_0           = AXI4L_OSD_ARBURST;
assign AXI4L_OSD_SLAVE5_ARBURST[1:0]     = AXI4L_OSD_ARBURST_net_0;
assign AXI4L_OSD_ARCACHE_net_0           = AXI4L_OSD_ARCACHE;
assign AXI4L_OSD_SLAVE5_ARCACHE[3:0]     = AXI4L_OSD_ARCACHE_net_0;
assign AXI4L_OSD_ARID_net_0              = AXI4L_OSD_ARID;
assign AXI4L_OSD_SLAVE5_ARID[8:0]        = AXI4L_OSD_ARID_net_0;
assign AXI4L_OSD_ARLEN_net_0             = AXI4L_OSD_ARLEN;
assign AXI4L_OSD_SLAVE5_ARLEN[7:0]       = AXI4L_OSD_ARLEN_net_0;
assign AXI4L_OSD_ARLOCK_net_0            = AXI4L_OSD_ARLOCK;
assign AXI4L_OSD_SLAVE5_ARLOCK[1:0]      = AXI4L_OSD_ARLOCK_net_0;
assign AXI4L_OSD_ARPROT_net_0            = AXI4L_OSD_ARPROT;
assign AXI4L_OSD_SLAVE5_ARPROT[2:0]      = AXI4L_OSD_ARPROT_net_0;
assign AXI4L_OSD_ARQOS_net_0             = AXI4L_OSD_ARQOS;
assign AXI4L_OSD_SLAVE5_ARQOS[3:0]       = AXI4L_OSD_ARQOS_net_0;
assign AXI4L_OSD_ARREGION_net_0          = AXI4L_OSD_ARREGION;
assign AXI4L_OSD_SLAVE5_ARREGION[3:0]    = AXI4L_OSD_ARREGION_net_0;
assign AXI4L_OSD_ARSIZE_net_0            = AXI4L_OSD_ARSIZE;
assign AXI4L_OSD_SLAVE5_ARSIZE[2:0]      = AXI4L_OSD_ARSIZE_net_0;
assign AXI4L_OSD_ARUSER_net_0[0]         = AXI4L_OSD_ARUSER[0];
assign AXI4L_OSD_SLAVE5_ARUSER[0:0]      = AXI4L_OSD_ARUSER_net_0[0];
assign AXI4L_OSD_AWADDR_net_0            = AXI4L_OSD_AWADDR;
assign AXI4L_OSD_SLAVE5_AWADDR[37:0]     = AXI4L_OSD_AWADDR_net_0;
assign AXI4L_OSD_AWBURST_net_0           = AXI4L_OSD_AWBURST;
assign AXI4L_OSD_SLAVE5_AWBURST[1:0]     = AXI4L_OSD_AWBURST_net_0;
assign AXI4L_OSD_AWCACHE_net_0           = AXI4L_OSD_AWCACHE;
assign AXI4L_OSD_SLAVE5_AWCACHE[3:0]     = AXI4L_OSD_AWCACHE_net_0;
assign AXI4L_OSD_AWID_net_0              = AXI4L_OSD_AWID;
assign AXI4L_OSD_SLAVE5_AWID[8:0]        = AXI4L_OSD_AWID_net_0;
assign AXI4L_OSD_AWLEN_net_0             = AXI4L_OSD_AWLEN;
assign AXI4L_OSD_SLAVE5_AWLEN[7:0]       = AXI4L_OSD_AWLEN_net_0;
assign AXI4L_OSD_AWLOCK_net_0            = AXI4L_OSD_AWLOCK;
assign AXI4L_OSD_SLAVE5_AWLOCK[1:0]      = AXI4L_OSD_AWLOCK_net_0;
assign AXI4L_OSD_AWPROT_net_0            = AXI4L_OSD_AWPROT;
assign AXI4L_OSD_SLAVE5_AWPROT[2:0]      = AXI4L_OSD_AWPROT_net_0;
assign AXI4L_OSD_AWQOS_net_0             = AXI4L_OSD_AWQOS;
assign AXI4L_OSD_SLAVE5_AWQOS[3:0]       = AXI4L_OSD_AWQOS_net_0;
assign AXI4L_OSD_AWREGION_net_0          = AXI4L_OSD_AWREGION;
assign AXI4L_OSD_SLAVE5_AWREGION[3:0]    = AXI4L_OSD_AWREGION_net_0;
assign AXI4L_OSD_AWSIZE_net_0            = AXI4L_OSD_AWSIZE;
assign AXI4L_OSD_SLAVE5_AWSIZE[2:0]      = AXI4L_OSD_AWSIZE_net_0;
assign AXI4L_OSD_AWUSER_net_0[0]         = AXI4L_OSD_AWUSER[0];
assign AXI4L_OSD_SLAVE5_AWUSER[0:0]      = AXI4L_OSD_AWUSER_net_0[0];
assign AXI4L_OSD_WDATA_net_0             = AXI4L_OSD_WDATA;
assign AXI4L_OSD_SLAVE5_WDATA[63:0]      = AXI4L_OSD_WDATA_net_0;
assign AXI4L_OSD_WSTRB_net_0             = AXI4L_OSD_WSTRB;
assign AXI4L_OSD_SLAVE5_WSTRB[7:0]       = AXI4L_OSD_WSTRB_net_0;
assign AXI4L_OSD_WUSER_net_0[0]          = AXI4L_OSD_WUSER[0];
assign AXI4L_OSD_SLAVE5_WUSER[0:0]       = AXI4L_OSD_WUSER_net_0[0];
assign AXI4L_SCALER_ARADDR_net_0         = AXI4L_SCALER_ARADDR;
assign AXI4L_SCALER_SLAVE4_ARADDR[37:0]  = AXI4L_SCALER_ARADDR_net_0;
assign AXI4L_SCALER_ARBURST_net_0        = AXI4L_SCALER_ARBURST;
assign AXI4L_SCALER_SLAVE4_ARBURST[1:0]  = AXI4L_SCALER_ARBURST_net_0;
assign AXI4L_SCALER_ARCACHE_net_0        = AXI4L_SCALER_ARCACHE;
assign AXI4L_SCALER_SLAVE4_ARCACHE[3:0]  = AXI4L_SCALER_ARCACHE_net_0;
assign AXI4L_SCALER_ARID_net_0           = AXI4L_SCALER_ARID;
assign AXI4L_SCALER_SLAVE4_ARID[8:0]     = AXI4L_SCALER_ARID_net_0;
assign AXI4L_SCALER_ARLEN_net_0          = AXI4L_SCALER_ARLEN;
assign AXI4L_SCALER_SLAVE4_ARLEN[7:0]    = AXI4L_SCALER_ARLEN_net_0;
assign AXI4L_SCALER_ARLOCK_net_0         = AXI4L_SCALER_ARLOCK;
assign AXI4L_SCALER_SLAVE4_ARLOCK[1:0]   = AXI4L_SCALER_ARLOCK_net_0;
assign AXI4L_SCALER_ARPROT_net_0         = AXI4L_SCALER_ARPROT;
assign AXI4L_SCALER_SLAVE4_ARPROT[2:0]   = AXI4L_SCALER_ARPROT_net_0;
assign AXI4L_SCALER_ARQOS_net_0          = AXI4L_SCALER_ARQOS;
assign AXI4L_SCALER_SLAVE4_ARQOS[3:0]    = AXI4L_SCALER_ARQOS_net_0;
assign AXI4L_SCALER_ARREGION_net_0       = AXI4L_SCALER_ARREGION;
assign AXI4L_SCALER_SLAVE4_ARREGION[3:0] = AXI4L_SCALER_ARREGION_net_0;
assign AXI4L_SCALER_ARSIZE_net_0         = AXI4L_SCALER_ARSIZE;
assign AXI4L_SCALER_SLAVE4_ARSIZE[2:0]   = AXI4L_SCALER_ARSIZE_net_0;
assign AXI4L_SCALER_ARUSER_net_0[0]      = AXI4L_SCALER_ARUSER[0];
assign AXI4L_SCALER_SLAVE4_ARUSER[0:0]   = AXI4L_SCALER_ARUSER_net_0[0];
assign AXI4L_SCALER_AWADDR_net_0         = AXI4L_SCALER_AWADDR;
assign AXI4L_SCALER_SLAVE4_AWADDR[37:0]  = AXI4L_SCALER_AWADDR_net_0;
assign AXI4L_SCALER_AWBURST_net_0        = AXI4L_SCALER_AWBURST;
assign AXI4L_SCALER_SLAVE4_AWBURST[1:0]  = AXI4L_SCALER_AWBURST_net_0;
assign AXI4L_SCALER_AWCACHE_net_0        = AXI4L_SCALER_AWCACHE;
assign AXI4L_SCALER_SLAVE4_AWCACHE[3:0]  = AXI4L_SCALER_AWCACHE_net_0;
assign AXI4L_SCALER_AWID_net_0           = AXI4L_SCALER_AWID;
assign AXI4L_SCALER_SLAVE4_AWID[8:0]     = AXI4L_SCALER_AWID_net_0;
assign AXI4L_SCALER_AWLEN_net_0          = AXI4L_SCALER_AWLEN;
assign AXI4L_SCALER_SLAVE4_AWLEN[7:0]    = AXI4L_SCALER_AWLEN_net_0;
assign AXI4L_SCALER_AWLOCK_net_0         = AXI4L_SCALER_AWLOCK;
assign AXI4L_SCALER_SLAVE4_AWLOCK[1:0]   = AXI4L_SCALER_AWLOCK_net_0;
assign AXI4L_SCALER_AWPROT_net_0         = AXI4L_SCALER_AWPROT;
assign AXI4L_SCALER_SLAVE4_AWPROT[2:0]   = AXI4L_SCALER_AWPROT_net_0;
assign AXI4L_SCALER_AWQOS_net_0          = AXI4L_SCALER_AWQOS;
assign AXI4L_SCALER_SLAVE4_AWQOS[3:0]    = AXI4L_SCALER_AWQOS_net_0;
assign AXI4L_SCALER_AWREGION_net_0       = AXI4L_SCALER_AWREGION;
assign AXI4L_SCALER_SLAVE4_AWREGION[3:0] = AXI4L_SCALER_AWREGION_net_0;
assign AXI4L_SCALER_AWSIZE_net_0         = AXI4L_SCALER_AWSIZE;
assign AXI4L_SCALER_SLAVE4_AWSIZE[2:0]   = AXI4L_SCALER_AWSIZE_net_0;
assign AXI4L_SCALER_AWUSER_net_0[0]      = AXI4L_SCALER_AWUSER[0];
assign AXI4L_SCALER_SLAVE4_AWUSER[0:0]   = AXI4L_SCALER_AWUSER_net_0[0];
assign AXI4L_SCALER_WDATA_net_0          = AXI4L_SCALER_WDATA;
assign AXI4L_SCALER_SLAVE4_WDATA[63:0]   = AXI4L_SCALER_WDATA_net_0;
assign AXI4L_SCALER_WSTRB_net_0          = AXI4L_SCALER_WSTRB;
assign AXI4L_SCALER_SLAVE4_WSTRB[7:0]    = AXI4L_SCALER_WSTRB_net_0;
assign AXI4L_SCALER_WUSER_net_0[0]       = AXI4L_SCALER_WUSER[0];
assign AXI4L_SCALER_SLAVE4_WUSER[0:0]    = AXI4L_SCALER_WUSER_net_0[0];
assign AXI4L_VDMA_ARADDR_net_0           = AXI4L_VDMA_ARADDR;
assign AXI4L_VDMA_SLAVE0_ARADDR[37:0]    = AXI4L_VDMA_ARADDR_net_0;
assign AXI4L_VDMA_ARBURST_net_0          = AXI4L_VDMA_ARBURST;
assign AXI4L_VDMA_SLAVE0_ARBURST[1:0]    = AXI4L_VDMA_ARBURST_net_0;
assign AXI4L_VDMA_ARCACHE_net_0          = AXI4L_VDMA_ARCACHE;
assign AXI4L_VDMA_SLAVE0_ARCACHE[3:0]    = AXI4L_VDMA_ARCACHE_net_0;
assign AXI4L_VDMA_ARID_net_0             = AXI4L_VDMA_ARID;
assign AXI4L_VDMA_SLAVE0_ARID[8:0]       = AXI4L_VDMA_ARID_net_0;
assign AXI4L_VDMA_ARLEN_net_0            = AXI4L_VDMA_ARLEN;
assign AXI4L_VDMA_SLAVE0_ARLEN[7:0]      = AXI4L_VDMA_ARLEN_net_0;
assign AXI4L_VDMA_ARLOCK_net_0           = AXI4L_VDMA_ARLOCK;
assign AXI4L_VDMA_SLAVE0_ARLOCK[1:0]     = AXI4L_VDMA_ARLOCK_net_0;
assign AXI4L_VDMA_ARPROT_net_0           = AXI4L_VDMA_ARPROT;
assign AXI4L_VDMA_SLAVE0_ARPROT[2:0]     = AXI4L_VDMA_ARPROT_net_0;
assign AXI4L_VDMA_ARQOS_net_0            = AXI4L_VDMA_ARQOS;
assign AXI4L_VDMA_SLAVE0_ARQOS[3:0]      = AXI4L_VDMA_ARQOS_net_0;
assign AXI4L_VDMA_ARREGION_net_0         = AXI4L_VDMA_ARREGION;
assign AXI4L_VDMA_SLAVE0_ARREGION[3:0]   = AXI4L_VDMA_ARREGION_net_0;
assign AXI4L_VDMA_ARSIZE_net_0           = AXI4L_VDMA_ARSIZE;
assign AXI4L_VDMA_SLAVE0_ARSIZE[2:0]     = AXI4L_VDMA_ARSIZE_net_0;
assign AXI4L_VDMA_ARUSER_net_0[0]        = AXI4L_VDMA_ARUSER[0];
assign AXI4L_VDMA_SLAVE0_ARUSER[0:0]     = AXI4L_VDMA_ARUSER_net_0[0];
assign AXI4L_VDMA_AWADDR_net_0           = AXI4L_VDMA_AWADDR;
assign AXI4L_VDMA_SLAVE0_AWADDR[37:0]    = AXI4L_VDMA_AWADDR_net_0;
assign AXI4L_VDMA_AWBURST_net_0          = AXI4L_VDMA_AWBURST;
assign AXI4L_VDMA_SLAVE0_AWBURST[1:0]    = AXI4L_VDMA_AWBURST_net_0;
assign AXI4L_VDMA_AWCACHE_net_0          = AXI4L_VDMA_AWCACHE;
assign AXI4L_VDMA_SLAVE0_AWCACHE[3:0]    = AXI4L_VDMA_AWCACHE_net_0;
assign AXI4L_VDMA_AWID_net_0             = AXI4L_VDMA_AWID;
assign AXI4L_VDMA_SLAVE0_AWID[8:0]       = AXI4L_VDMA_AWID_net_0;
assign AXI4L_VDMA_AWLEN_net_0            = AXI4L_VDMA_AWLEN;
assign AXI4L_VDMA_SLAVE0_AWLEN[7:0]      = AXI4L_VDMA_AWLEN_net_0;
assign AXI4L_VDMA_AWLOCK_net_0           = AXI4L_VDMA_AWLOCK;
assign AXI4L_VDMA_SLAVE0_AWLOCK[1:0]     = AXI4L_VDMA_AWLOCK_net_0;
assign AXI4L_VDMA_AWPROT_net_0           = AXI4L_VDMA_AWPROT;
assign AXI4L_VDMA_SLAVE0_AWPROT[2:0]     = AXI4L_VDMA_AWPROT_net_0;
assign AXI4L_VDMA_AWQOS_net_0            = AXI4L_VDMA_AWQOS;
assign AXI4L_VDMA_SLAVE0_AWQOS[3:0]      = AXI4L_VDMA_AWQOS_net_0;
assign AXI4L_VDMA_AWREGION_net_0         = AXI4L_VDMA_AWREGION;
assign AXI4L_VDMA_SLAVE0_AWREGION[3:0]   = AXI4L_VDMA_AWREGION_net_0;
assign AXI4L_VDMA_AWSIZE_net_0           = AXI4L_VDMA_AWSIZE;
assign AXI4L_VDMA_SLAVE0_AWSIZE[2:0]     = AXI4L_VDMA_AWSIZE_net_0;
assign AXI4L_VDMA_AWUSER_net_0[0]        = AXI4L_VDMA_AWUSER[0];
assign AXI4L_VDMA_SLAVE0_AWUSER[0:0]     = AXI4L_VDMA_AWUSER_net_0[0];
assign AXI4L_VDMA_WDATA_net_0            = AXI4L_VDMA_WDATA;
assign AXI4L_VDMA_SLAVE0_WDATA[31:0]     = AXI4L_VDMA_WDATA_net_0;
assign AXI4L_VDMA_WSTRB_net_0            = AXI4L_VDMA_WSTRB;
assign AXI4L_VDMA_SLAVE0_WSTRB[3:0]      = AXI4L_VDMA_WSTRB_net_0;
assign AXI4L_VDMA_WUSER_net_0[0]         = AXI4L_VDMA_WUSER[0];
assign AXI4L_VDMA_SLAVE0_WUSER[0:0]      = AXI4L_VDMA_WUSER_net_0[0];
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------COREAXI4INTERCONNECT_C0
COREAXI4INTERCONNECT_C0 COREAXI4INTERCONNECT_C0_0(
        // Inputs
        .ACLK             ( ACLK ),
        .ARESETN          ( ARESETN ),
        .SLAVE0_AWREADY   ( AXI4L_VDMA_SLAVE0_AWREADY ),
        .SLAVE0_WREADY    ( AXI4L_VDMA_SLAVE0_WREADY ),
        .SLAVE0_BID       ( AXI4L_VDMA_SLAVE0_BID ),
        .SLAVE0_BRESP     ( AXI4L_VDMA_SLAVE0_BRESP ),
        .SLAVE0_BVALID    ( AXI4L_VDMA_SLAVE0_BVALID ),
        .SLAVE0_ARREADY   ( AXI4L_VDMA_SLAVE0_ARREADY ),
        .SLAVE0_RID       ( AXI4L_VDMA_SLAVE0_RID ),
        .SLAVE0_RDATA     ( AXI4L_VDMA_SLAVE0_RDATA ),
        .SLAVE0_RRESP     ( AXI4L_VDMA_SLAVE0_RRESP ),
        .SLAVE0_RLAST     ( AXI4L_VDMA_SLAVE0_RLAST ),
        .SLAVE0_RVALID    ( AXI4L_VDMA_SLAVE0_RVALID ),
        .SLAVE0_BUSER     ( AXI4L_VDMA_SLAVE0_BUSER ),
        .SLAVE0_RUSER     ( AXI4L_VDMA_SLAVE0_RUSER ),
        .SLAVE1_AWREADY   ( AXI4L_MIPI_SLAVE1_AWREADY ),
        .SLAVE1_WREADY    ( AXI4L_MIPI_SLAVE1_WREADY ),
        .SLAVE1_BID       ( AXI4L_MIPI_SLAVE1_BID ),
        .SLAVE1_BRESP     ( AXI4L_MIPI_SLAVE1_BRESP ),
        .SLAVE1_BVALID    ( AXI4L_MIPI_SLAVE1_BVALID ),
        .SLAVE1_ARREADY   ( AXI4L_MIPI_SLAVE1_ARREADY ),
        .SLAVE1_RID       ( AXI4L_MIPI_SLAVE1_RID ),
        .SLAVE1_RDATA     ( AXI4L_MIPI_SLAVE1_RDATA ),
        .SLAVE1_RRESP     ( AXI4L_MIPI_SLAVE1_RRESP ),
        .SLAVE1_RLAST     ( AXI4L_MIPI_SLAVE1_RLAST ),
        .SLAVE1_RVALID    ( AXI4L_MIPI_SLAVE1_RVALID ),
        .SLAVE1_BUSER     ( AXI4L_MIPI_SLAVE1_BUSER ),
        .SLAVE1_RUSER     ( AXI4L_MIPI_SLAVE1_RUSER ),
        .SLAVE2_AWREADY   ( AXI4L_H264_SLAVE2_AWREADY ),
        .SLAVE2_WREADY    ( AXI4L_H264_SLAVE2_WREADY ),
        .SLAVE2_BID       ( AXI4L_H264_SLAVE2_BID ),
        .SLAVE2_BRESP     ( AXI4L_H264_SLAVE2_BRESP ),
        .SLAVE2_BVALID    ( AXI4L_H264_SLAVE2_BVALID ),
        .SLAVE2_ARREADY   ( AXI4L_H264_SLAVE2_ARREADY ),
        .SLAVE2_RID       ( AXI4L_H264_SLAVE2_RID ),
        .SLAVE2_RDATA     ( AXI4L_H264_SLAVE2_RDATA ),
        .SLAVE2_RRESP     ( AXI4L_H264_SLAVE2_RRESP ),
        .SLAVE2_RLAST     ( AXI4L_H264_SLAVE2_RLAST ),
        .SLAVE2_RVALID    ( AXI4L_H264_SLAVE2_RVALID ),
        .SLAVE2_BUSER     ( AXI4L_H264_SLAVE2_BUSER ),
        .SLAVE2_RUSER     ( AXI4L_H264_SLAVE2_RUSER ),
        .SLAVE3_AWREADY   ( AXI4L_IE_SLAVE3_AWREADY ),
        .SLAVE3_WREADY    ( AXI4L_IE_SLAVE3_WREADY ),
        .SLAVE3_BID       ( AXI4L_IE_SLAVE3_BID ),
        .SLAVE3_BRESP     ( AXI4L_IE_SLAVE3_BRESP ),
        .SLAVE3_BVALID    ( AXI4L_IE_SLAVE3_BVALID ),
        .SLAVE3_ARREADY   ( AXI4L_IE_SLAVE3_ARREADY ),
        .SLAVE3_RID       ( AXI4L_IE_SLAVE3_RID ),
        .SLAVE3_RDATA     ( AXI4L_IE_SLAVE3_RDATA ),
        .SLAVE3_RRESP     ( AXI4L_IE_SLAVE3_RRESP ),
        .SLAVE3_RLAST     ( AXI4L_IE_SLAVE3_RLAST ),
        .SLAVE3_RVALID    ( AXI4L_IE_SLAVE3_RVALID ),
        .SLAVE3_BUSER     ( AXI4L_IE_SLAVE3_BUSER ),
        .SLAVE3_RUSER     ( AXI4L_IE_SLAVE3_RUSER ),
        .SLAVE4_AWREADY   ( AXI4L_SCALER_SLAVE4_AWREADY ),
        .SLAVE4_WREADY    ( AXI4L_SCALER_SLAVE4_WREADY ),
        .SLAVE4_BID       ( AXI4L_SCALER_SLAVE4_BID ),
        .SLAVE4_BRESP     ( AXI4L_SCALER_SLAVE4_BRESP ),
        .SLAVE4_BVALID    ( AXI4L_SCALER_SLAVE4_BVALID ),
        .SLAVE4_ARREADY   ( AXI4L_SCALER_SLAVE4_ARREADY ),
        .SLAVE4_RID       ( AXI4L_SCALER_SLAVE4_RID ),
        .SLAVE4_RDATA     ( AXI4L_SCALER_SLAVE4_RDATA ),
        .SLAVE4_RRESP     ( AXI4L_SCALER_SLAVE4_RRESP ),
        .SLAVE4_RLAST     ( AXI4L_SCALER_SLAVE4_RLAST ),
        .SLAVE4_RVALID    ( AXI4L_SCALER_SLAVE4_RVALID ),
        .SLAVE4_BUSER     ( AXI4L_SCALER_SLAVE4_BUSER ),
        .SLAVE4_RUSER     ( AXI4L_SCALER_SLAVE4_RUSER ),
        .SLAVE5_AWREADY   ( AXI4L_OSD_SLAVE5_AWREADY ),
        .SLAVE5_WREADY    ( AXI4L_OSD_SLAVE5_WREADY ),
        .SLAVE5_BID       ( AXI4L_OSD_SLAVE5_BID ),
        .SLAVE5_BRESP     ( AXI4L_OSD_SLAVE5_BRESP ),
        .SLAVE5_BVALID    ( AXI4L_OSD_SLAVE5_BVALID ),
        .SLAVE5_ARREADY   ( AXI4L_OSD_SLAVE5_ARREADY ),
        .SLAVE5_RID       ( AXI4L_OSD_SLAVE5_RID ),
        .SLAVE5_RDATA     ( AXI4L_OSD_SLAVE5_RDATA ),
        .SLAVE5_RRESP     ( AXI4L_OSD_SLAVE5_RRESP ),
        .SLAVE5_RLAST     ( AXI4L_OSD_SLAVE5_RLAST ),
        .SLAVE5_RVALID    ( AXI4L_OSD_SLAVE5_RVALID ),
        .SLAVE5_BUSER     ( AXI4L_OSD_SLAVE5_BUSER ),
        .SLAVE5_RUSER     ( AXI4L_OSD_SLAVE5_RUSER ),
        .MASTER0_AWID     ( AXI4L_MASTER0_AWID ),
        .MASTER0_AWADDR   ( AXI4L_MASTER0_AWADDR ),
        .MASTER0_AWLEN    ( AXI4L_MASTER0_AWLEN ),
        .MASTER0_AWSIZE   ( AXI4L_MASTER0_AWSIZE ),
        .MASTER0_AWBURST  ( AXI4L_MASTER0_AWBURST ),
        .MASTER0_AWLOCK   ( AXI4L_MASTER0_AWLOCK ),
        .MASTER0_AWCACHE  ( AXI4L_MASTER0_AWCACHE ),
        .MASTER0_AWPROT   ( AXI4L_MASTER0_AWPROT ),
        .MASTER0_AWQOS    ( AXI4L_MASTER0_AWQOS ),
        .MASTER0_AWREGION ( AXI4L_MASTER0_AWREGION ),
        .MASTER0_AWVALID  ( AXI4L_MASTER0_AWVALID ),
        .MASTER0_WDATA    ( AXI4L_MASTER0_WDATA ),
        .MASTER0_WSTRB    ( AXI4L_MASTER0_WSTRB ),
        .MASTER0_WLAST    ( AXI4L_MASTER0_WLAST ),
        .MASTER0_WVALID   ( AXI4L_MASTER0_WVALID ),
        .MASTER0_BREADY   ( AXI4L_MASTER0_BREADY ),
        .MASTER0_ARID     ( AXI4L_MASTER0_ARID ),
        .MASTER0_ARADDR   ( AXI4L_MASTER0_ARADDR ),
        .MASTER0_ARLEN    ( AXI4L_MASTER0_ARLEN ),
        .MASTER0_ARSIZE   ( AXI4L_MASTER0_ARSIZE ),
        .MASTER0_ARBURST  ( AXI4L_MASTER0_ARBURST ),
        .MASTER0_ARLOCK   ( AXI4L_MASTER0_ARLOCK ),
        .MASTER0_ARCACHE  ( AXI4L_MASTER0_ARCACHE ),
        .MASTER0_ARPROT   ( AXI4L_MASTER0_ARPROT ),
        .MASTER0_ARQOS    ( AXI4L_MASTER0_ARQOS ),
        .MASTER0_ARREGION ( AXI4L_MASTER0_ARREGION ),
        .MASTER0_ARVALID  ( AXI4L_MASTER0_ARVALID ),
        .MASTER0_RREADY   ( AXI4L_MASTER0_RREADY ),
        .MASTER0_AWUSER   ( AXI4L_MASTER0_AWUSER ),
        .MASTER0_WUSER    ( AXI4L_MASTER0_WUSER ),
        .MASTER0_ARUSER   ( AXI4L_MASTER0_ARUSER ),
        // Outputs
        .SLAVE0_AWID      ( AXI4L_VDMA_AWID ),
        .SLAVE0_AWADDR    ( AXI4L_VDMA_AWADDR ),
        .SLAVE0_AWLEN     ( AXI4L_VDMA_AWLEN ),
        .SLAVE0_AWSIZE    ( AXI4L_VDMA_AWSIZE ),
        .SLAVE0_AWBURST   ( AXI4L_VDMA_AWBURST ),
        .SLAVE0_AWLOCK    ( AXI4L_VDMA_AWLOCK ),
        .SLAVE0_AWCACHE   ( AXI4L_VDMA_AWCACHE ),
        .SLAVE0_AWPROT    ( AXI4L_VDMA_AWPROT ),
        .SLAVE0_AWQOS     ( AXI4L_VDMA_AWQOS ),
        .SLAVE0_AWREGION  ( AXI4L_VDMA_AWREGION ),
        .SLAVE0_AWVALID   ( AXI4L_VDMA_AWVALID ),
        .SLAVE0_WDATA     ( AXI4L_VDMA_WDATA ),
        .SLAVE0_WSTRB     ( AXI4L_VDMA_WSTRB ),
        .SLAVE0_WLAST     ( AXI4L_VDMA_WLAST ),
        .SLAVE0_WVALID    ( AXI4L_VDMA_WVALID ),
        .SLAVE0_BREADY    ( AXI4L_VDMA_BREADY ),
        .SLAVE0_ARID      ( AXI4L_VDMA_ARID ),
        .SLAVE0_ARADDR    ( AXI4L_VDMA_ARADDR ),
        .SLAVE0_ARLEN     ( AXI4L_VDMA_ARLEN ),
        .SLAVE0_ARSIZE    ( AXI4L_VDMA_ARSIZE ),
        .SLAVE0_ARBURST   ( AXI4L_VDMA_ARBURST ),
        .SLAVE0_ARLOCK    ( AXI4L_VDMA_ARLOCK ),
        .SLAVE0_ARCACHE   ( AXI4L_VDMA_ARCACHE ),
        .SLAVE0_ARPROT    ( AXI4L_VDMA_ARPROT ),
        .SLAVE0_ARQOS     ( AXI4L_VDMA_ARQOS ),
        .SLAVE0_ARREGION  ( AXI4L_VDMA_ARREGION ),
        .SLAVE0_ARVALID   ( AXI4L_VDMA_ARVALID ),
        .SLAVE0_RREADY    ( AXI4L_VDMA_RREADY ),
        .SLAVE0_AWUSER    ( AXI4L_VDMA_AWUSER ),
        .SLAVE0_WUSER     ( AXI4L_VDMA_WUSER ),
        .SLAVE0_ARUSER    ( AXI4L_VDMA_ARUSER ),
        .SLAVE1_AWID      ( AXI4L_MIPI_AWID ),
        .SLAVE1_AWADDR    ( AXI4L_MIPI_AWADDR ),
        .SLAVE1_AWLEN     ( AXI4L_MIPI_AWLEN ),
        .SLAVE1_AWSIZE    ( AXI4L_MIPI_AWSIZE ),
        .SLAVE1_AWBURST   ( AXI4L_MIPI_AWBURST ),
        .SLAVE1_AWLOCK    ( AXI4L_MIPI_AWLOCK ),
        .SLAVE1_AWCACHE   ( AXI4L_MIPI_AWCACHE ),
        .SLAVE1_AWPROT    ( AXI4L_MIPI_AWPROT ),
        .SLAVE1_AWQOS     ( AXI4L_MIPI_AWQOS ),
        .SLAVE1_AWREGION  ( AXI4L_MIPI_AWREGION ),
        .SLAVE1_AWVALID   ( AXI4L_MIPI_AWVALID ),
        .SLAVE1_WDATA     ( AXI4L_MIPI_WDATA ),
        .SLAVE1_WSTRB     ( AXI4L_MIPI_WSTRB ),
        .SLAVE1_WLAST     ( AXI4L_MIPI_WLAST ),
        .SLAVE1_WVALID    ( AXI4L_MIPI_WVALID ),
        .SLAVE1_BREADY    ( AXI4L_MIPI_BREADY ),
        .SLAVE1_ARID      ( AXI4L_MIPI_ARID ),
        .SLAVE1_ARADDR    ( AXI4L_MIPI_ARADDR ),
        .SLAVE1_ARLEN     ( AXI4L_MIPI_ARLEN ),
        .SLAVE1_ARSIZE    ( AXI4L_MIPI_ARSIZE ),
        .SLAVE1_ARBURST   ( AXI4L_MIPI_ARBURST ),
        .SLAVE1_ARLOCK    ( AXI4L_MIPI_ARLOCK ),
        .SLAVE1_ARCACHE   ( AXI4L_MIPI_ARCACHE ),
        .SLAVE1_ARPROT    ( AXI4L_MIPI_ARPROT ),
        .SLAVE1_ARQOS     ( AXI4L_MIPI_ARQOS ),
        .SLAVE1_ARREGION  ( AXI4L_MIPI_ARREGION ),
        .SLAVE1_ARVALID   ( AXI4L_MIPI_ARVALID ),
        .SLAVE1_RREADY    ( AXI4L_MIPI_RREADY ),
        .SLAVE1_AWUSER    ( AXI4L_MIPI_AWUSER ),
        .SLAVE1_WUSER     ( AXI4L_MIPI_WUSER ),
        .SLAVE1_ARUSER    ( AXI4L_MIPI_ARUSER ),
        .SLAVE2_AWID      ( AXI4L_H264_AWID ),
        .SLAVE2_AWADDR    ( AXI4L_H264_AWADDR ),
        .SLAVE2_AWLEN     ( AXI4L_H264_AWLEN ),
        .SLAVE2_AWSIZE    ( AXI4L_H264_AWSIZE ),
        .SLAVE2_AWBURST   ( AXI4L_H264_AWBURST ),
        .SLAVE2_AWLOCK    ( AXI4L_H264_AWLOCK ),
        .SLAVE2_AWCACHE   ( AXI4L_H264_AWCACHE ),
        .SLAVE2_AWPROT    ( AXI4L_H264_AWPROT ),
        .SLAVE2_AWQOS     ( AXI4L_H264_AWQOS ),
        .SLAVE2_AWREGION  ( AXI4L_H264_AWREGION ),
        .SLAVE2_AWVALID   ( AXI4L_H264_AWVALID ),
        .SLAVE2_WDATA     ( AXI4L_H264_WDATA ),
        .SLAVE2_WSTRB     ( AXI4L_H264_WSTRB ),
        .SLAVE2_WLAST     ( AXI4L_H264_WLAST ),
        .SLAVE2_WVALID    ( AXI4L_H264_WVALID ),
        .SLAVE2_BREADY    ( AXI4L_H264_BREADY ),
        .SLAVE2_ARID      ( AXI4L_H264_ARID ),
        .SLAVE2_ARADDR    ( AXI4L_H264_ARADDR ),
        .SLAVE2_ARLEN     ( AXI4L_H264_ARLEN ),
        .SLAVE2_ARSIZE    ( AXI4L_H264_ARSIZE ),
        .SLAVE2_ARBURST   ( AXI4L_H264_ARBURST ),
        .SLAVE2_ARLOCK    ( AXI4L_H264_ARLOCK ),
        .SLAVE2_ARCACHE   ( AXI4L_H264_ARCACHE ),
        .SLAVE2_ARPROT    ( AXI4L_H264_ARPROT ),
        .SLAVE2_ARQOS     ( AXI4L_H264_ARQOS ),
        .SLAVE2_ARREGION  ( AXI4L_H264_ARREGION ),
        .SLAVE2_ARVALID   ( AXI4L_H264_ARVALID ),
        .SLAVE2_RREADY    ( AXI4L_H264_RREADY ),
        .SLAVE2_AWUSER    ( AXI4L_H264_AWUSER ),
        .SLAVE2_WUSER     ( AXI4L_H264_WUSER ),
        .SLAVE2_ARUSER    ( AXI4L_H264_ARUSER ),
        .SLAVE3_AWID      ( AXI4L_IE_AWID ),
        .SLAVE3_AWADDR    ( AXI4L_IE_AWADDR ),
        .SLAVE3_AWLEN     ( AXI4L_IE_AWLEN ),
        .SLAVE3_AWSIZE    ( AXI4L_IE_AWSIZE ),
        .SLAVE3_AWBURST   ( AXI4L_IE_AWBURST ),
        .SLAVE3_AWLOCK    ( AXI4L_IE_AWLOCK ),
        .SLAVE3_AWCACHE   ( AXI4L_IE_AWCACHE ),
        .SLAVE3_AWPROT    ( AXI4L_IE_AWPROT ),
        .SLAVE3_AWQOS     ( AXI4L_IE_AWQOS ),
        .SLAVE3_AWREGION  ( AXI4L_IE_AWREGION ),
        .SLAVE3_AWVALID   ( AXI4L_IE_AWVALID ),
        .SLAVE3_WDATA     ( AXI4L_IE_WDATA ),
        .SLAVE3_WSTRB     ( AXI4L_IE_WSTRB ),
        .SLAVE3_WLAST     ( AXI4L_IE_WLAST ),
        .SLAVE3_WVALID    ( AXI4L_IE_WVALID ),
        .SLAVE3_BREADY    ( AXI4L_IE_BREADY ),
        .SLAVE3_ARID      ( AXI4L_IE_ARID ),
        .SLAVE3_ARADDR    ( AXI4L_IE_ARADDR ),
        .SLAVE3_ARLEN     ( AXI4L_IE_ARLEN ),
        .SLAVE3_ARSIZE    ( AXI4L_IE_ARSIZE ),
        .SLAVE3_ARBURST   ( AXI4L_IE_ARBURST ),
        .SLAVE3_ARLOCK    ( AXI4L_IE_ARLOCK ),
        .SLAVE3_ARCACHE   ( AXI4L_IE_ARCACHE ),
        .SLAVE3_ARPROT    ( AXI4L_IE_ARPROT ),
        .SLAVE3_ARQOS     ( AXI4L_IE_ARQOS ),
        .SLAVE3_ARREGION  ( AXI4L_IE_ARREGION ),
        .SLAVE3_ARVALID   ( AXI4L_IE_ARVALID ),
        .SLAVE3_RREADY    ( AXI4L_IE_RREADY ),
        .SLAVE3_AWUSER    ( AXI4L_IE_AWUSER ),
        .SLAVE3_WUSER     ( AXI4L_IE_WUSER ),
        .SLAVE3_ARUSER    ( AXI4L_IE_ARUSER ),
        .SLAVE4_AWID      ( AXI4L_SCALER_AWID ),
        .SLAVE4_AWADDR    ( AXI4L_SCALER_AWADDR ),
        .SLAVE4_AWLEN     ( AXI4L_SCALER_AWLEN ),
        .SLAVE4_AWSIZE    ( AXI4L_SCALER_AWSIZE ),
        .SLAVE4_AWBURST   ( AXI4L_SCALER_AWBURST ),
        .SLAVE4_AWLOCK    ( AXI4L_SCALER_AWLOCK ),
        .SLAVE4_AWCACHE   ( AXI4L_SCALER_AWCACHE ),
        .SLAVE4_AWPROT    ( AXI4L_SCALER_AWPROT ),
        .SLAVE4_AWQOS     ( AXI4L_SCALER_AWQOS ),
        .SLAVE4_AWREGION  ( AXI4L_SCALER_AWREGION ),
        .SLAVE4_AWVALID   ( AXI4L_SCALER_AWVALID ),
        .SLAVE4_WDATA     ( AXI4L_SCALER_WDATA ),
        .SLAVE4_WSTRB     ( AXI4L_SCALER_WSTRB ),
        .SLAVE4_WLAST     ( AXI4L_SCALER_WLAST ),
        .SLAVE4_WVALID    ( AXI4L_SCALER_WVALID ),
        .SLAVE4_BREADY    ( AXI4L_SCALER_BREADY ),
        .SLAVE4_ARID      ( AXI4L_SCALER_ARID ),
        .SLAVE4_ARADDR    ( AXI4L_SCALER_ARADDR ),
        .SLAVE4_ARLEN     ( AXI4L_SCALER_ARLEN ),
        .SLAVE4_ARSIZE    ( AXI4L_SCALER_ARSIZE ),
        .SLAVE4_ARBURST   ( AXI4L_SCALER_ARBURST ),
        .SLAVE4_ARLOCK    ( AXI4L_SCALER_ARLOCK ),
        .SLAVE4_ARCACHE   ( AXI4L_SCALER_ARCACHE ),
        .SLAVE4_ARPROT    ( AXI4L_SCALER_ARPROT ),
        .SLAVE4_ARQOS     ( AXI4L_SCALER_ARQOS ),
        .SLAVE4_ARREGION  ( AXI4L_SCALER_ARREGION ),
        .SLAVE4_ARVALID   ( AXI4L_SCALER_ARVALID ),
        .SLAVE4_RREADY    ( AXI4L_SCALER_RREADY ),
        .SLAVE4_AWUSER    ( AXI4L_SCALER_AWUSER ),
        .SLAVE4_WUSER     ( AXI4L_SCALER_WUSER ),
        .SLAVE4_ARUSER    ( AXI4L_SCALER_ARUSER ),
        .SLAVE5_AWID      ( AXI4L_OSD_AWID ),
        .SLAVE5_AWADDR    ( AXI4L_OSD_AWADDR ),
        .SLAVE5_AWLEN     ( AXI4L_OSD_AWLEN ),
        .SLAVE5_AWSIZE    ( AXI4L_OSD_AWSIZE ),
        .SLAVE5_AWBURST   ( AXI4L_OSD_AWBURST ),
        .SLAVE5_AWLOCK    ( AXI4L_OSD_AWLOCK ),
        .SLAVE5_AWCACHE   ( AXI4L_OSD_AWCACHE ),
        .SLAVE5_AWPROT    ( AXI4L_OSD_AWPROT ),
        .SLAVE5_AWQOS     ( AXI4L_OSD_AWQOS ),
        .SLAVE5_AWREGION  ( AXI4L_OSD_AWREGION ),
        .SLAVE5_AWVALID   ( AXI4L_OSD_AWVALID ),
        .SLAVE5_WDATA     ( AXI4L_OSD_WDATA ),
        .SLAVE5_WSTRB     ( AXI4L_OSD_WSTRB ),
        .SLAVE5_WLAST     ( AXI4L_OSD_WLAST ),
        .SLAVE5_WVALID    ( AXI4L_OSD_WVALID ),
        .SLAVE5_BREADY    ( AXI4L_OSD_BREADY ),
        .SLAVE5_ARID      ( AXI4L_OSD_ARID ),
        .SLAVE5_ARADDR    ( AXI4L_OSD_ARADDR ),
        .SLAVE5_ARLEN     ( AXI4L_OSD_ARLEN ),
        .SLAVE5_ARSIZE    ( AXI4L_OSD_ARSIZE ),
        .SLAVE5_ARBURST   ( AXI4L_OSD_ARBURST ),
        .SLAVE5_ARLOCK    ( AXI4L_OSD_ARLOCK ),
        .SLAVE5_ARCACHE   ( AXI4L_OSD_ARCACHE ),
        .SLAVE5_ARPROT    ( AXI4L_OSD_ARPROT ),
        .SLAVE5_ARQOS     ( AXI4L_OSD_ARQOS ),
        .SLAVE5_ARREGION  ( AXI4L_OSD_ARREGION ),
        .SLAVE5_ARVALID   ( AXI4L_OSD_ARVALID ),
        .SLAVE5_RREADY    ( AXI4L_OSD_RREADY ),
        .SLAVE5_AWUSER    ( AXI4L_OSD_AWUSER ),
        .SLAVE5_WUSER     ( AXI4L_OSD_WUSER ),
        .SLAVE5_ARUSER    ( AXI4L_OSD_ARUSER ),
        .MASTER0_AWREADY  ( AXI4L_AWREADY ),
        .MASTER0_WREADY   ( AXI4L_WREADY ),
        .MASTER0_BID      ( AXI4L_BID ),
        .MASTER0_BRESP    ( AXI4L_BRESP ),
        .MASTER0_BVALID   ( AXI4L_BVALID ),
        .MASTER0_ARREADY  ( AXI4L_ARREADY ),
        .MASTER0_RID      ( AXI4L_RID ),
        .MASTER0_RDATA    ( AXI4L_RDATA ),
        .MASTER0_RRESP    ( AXI4L_RRESP ),
        .MASTER0_RLAST    ( AXI4L_RLAST ),
        .MASTER0_RVALID   ( AXI4L_RVALID ),
        .MASTER0_BUSER    ( AXI4L_BUSER ),
        .MASTER0_RUSER    ( AXI4L_RUSER ) 
        );


endmodule
