// --************************************************************************************************
// -- File Name                           : H264_Iframe_Encoder_Eval.v
// -- Targeted device                     : Microsemi-SoC
// -- Author                              : India Solutions Team
// --
// -- COPYRIGHT 2021 BY MICROSEMI
// -- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS FROM MICROSEMI
// -- CORP. IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM MICROSEMI FOR USE OF THIS
// -- FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND NO BACK-UP OF THE FILE SHOULD BE MADE.
// --
// --*************************************************************************************************

module H264_Iframe_Encoder #(
			     parameter G_DW 	  = 8,
			     parameter G_C_TYPE = 1,  // 0 - 400, 1 - 420
			     parameter G_16x16_INTRA_PRED = 1,
			     parameter G_HRES = 16'h780,
			     parameter G_VRES = 16'h430,
			     parameter G_QFACTOR = 6'h1E				     
			     )
   (
    // Clock and Reset interface----------------------------------------------------
    input wire 	      ACLK_I, // clock
    input wire 	      ARESETN_I, // This active-low reset
    //write address channel
    input wire 	      awvalid, // AXI4-Lite write address valid. This signal indicates that valid write address and control information are available.
    output reg 	      awready, // AXI4-Lite write address ready. This signal indicates that the target is ready to accept an address and associated control signals.
    input wire [31:0] awaddr, // AXI4-Lite write address.
    //write data channel
    input wire [31:0] wdata, // AXI4-Lite write data.
    input wire 	      wvalid, // AXI4-Lite write valid.
    output reg 	      wready, // AXI4-Lite Write ready.
    //write response channel
    output [1:0]      bresp, // AXI4-Lite write response.
    output reg 	      bvalid, // AXI4-Lite write response valid.
    input wire 	      bready, // AXI4-Lite response ready.
    //read address channel
    input wire [31:0] araddr, // AXI4-Lite read address. The read address gives the address of the first transfer in a read burst transaction.  
    input wire 	      arvalid, // AXI4-Lite read address valid. This signal indicates that the channel is signaling valid read address and control information. 
    output reg 	      arready, // AXI4-Lite response ready. This signal indicates that the slave is ready to accept an address and associated control signals.
    //read data and response channel
    input wire 	      rready, 
    output [31:0]     rdata, // AXI4-Lite read data.
    output [1:0]      rresp, // AXI4-Lite read response.
    output reg 	      rvalid, // AXI4-Lite read valid. This signal indicates that the channel is signaling the required read data.
    
    input 	      RESETN_I, 
    input 	      PIX_CLK_I,
    input 	      FRAME_START_I, // must be before frame start
    input 	      DATA_VALID_I,
    input [G_DW-1:0]  DATA_Y_I,
    input [G_DW-1:0]  DATA_C_I,
    output 	      FRAME_START_O,
    output 	      DATA_VALID_O,
    output [15:0]     DATA_O
    );   

   wire 	      resetn;
   wire 	      w_h264_ip_en;   
   wire 	      h264_ip_rstn;
   wire [5:0] 	      w_q_factor;
   wire [5:0] 	      w_ip_frame_gap;
   wire [15:0] 	      w_hres;
   wire [15:0] 	      w_vres;
   
   assign resetn = !h264_ip_rstn & RESETN_I;
   
   generate 
      H264_Iframe_Encoder_top #(
				 .G_DW(G_DW),
				 .G_C_TYPE(G_C_TYPE),
				 .G_16x16_INTRA_PRED(G_16x16_INTRA_PRED)
				 ) 
      H264_Iframe_Encoder_inst (
				.PIX_CLK(PIX_CLK_I),
				.RESET_N(resetn),
				.EN_I(w_h264_ip_en),
				.VRES_I(w_vres),
				.HRES_I(w_hres),
				.QP_I(w_q_factor),
				.FRAME_START_I(FRAME_START_I),
				.DATA_VALID_I(DATA_VALID_I),
				.DATA_Y_I(DATA_Y_I),
				.DATA_C_I(DATA_C_I),
				.FRAME_START_O(FRAME_START_O),
				.DATA_VALID_O(DATA_VALID_O),
				.DATA_O(DATA_O)
				);

      axi4lite_if_h264 #(.G_HRES(G_HRES), 
			 .G_VRES(G_VRES), 
			 .G_QFACTOR(G_QFACTOR)
			 )
      axi4lite_if_h264_inst
	(.*,
	 .h264_ip_en(w_h264_ip_en),
	 .h264_ip_rstn(h264_ip_rstn),
	 .q_factor(w_q_factor),
	 .i_p_frame_gap(w_ip_frame_gap),
	 .h_res(w_hres),
	 .v_res(w_vres)
	 );

   endgenerate
   
   
endmodule // H264_Iframe_Encoder






// --*************************************************************************************************
// -- File Name                           : axi4lite_if_h264.v
// -- Targeted device                     : Microsemi-SoC
// -- Author                              : India Solutions Team
// --
// -- COPYRIGHT 2021 BY MICROSEMI
// -- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS FROM MICROSEMI
// -- CORP. IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM MICROSEMI FOR USE OF THIS
// -- FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND NO BACK-UP OF THE FILE SHOULD BE MADE.
// --
// --*************************************************************************************************



localparam ADDR_DECODER_WIDTH = 8; //Address values of the registers
localparam IP_VER = 32'h0; //Read Only
localparam CTRL_REG = 32'h4; //Read Write
localparam IP_TYPE = 32'h8; //Read Only
localparam Q_FACTOR = 32'hC; //Write Only
localparam IN_FORMAT = 32'h10; //Read Only
localparam I_P_FRAME_GAP = 32'h14; //Write Only
localparam H_RES = 32'h18; //Write Only
localparam V_RES = 32'h1C; //Write Only


module axi4lite_if_h264 #(
			parameter G_HRES,
			parameter G_VRES,
			parameter G_QFACTOR
			)
  (
   // Clock and Reset interface----------------------------------------------------
   input wire 	     ACLK_I, // clock
   input wire 	     ARESETN_I, // This active-low reset
   //write address channel
   input wire 	     awvalid, // AXI4-Lite write address valid. This signal indicates that valid write address and control information are available.
   output reg 	     awready, // AXI4-Lite write address ready. This signal indicates that the target is ready to accept an address and associated control signals.
   input wire [31:0] awaddr, // AXI4-Lite write address.
   //write data channel
   input wire [31:0] wdata, // AXI4-Lite write data.
   input wire 	     wvalid, // AXI4-Lite write valid.
   output reg 	     wready, // AXI4-Lite Write ready.
   //write response channel
   output [1:0]      bresp, // AXI4-Lite write response.
   output reg 	     bvalid, // AXI4-Lite write response valid.
   input wire 	     bready, // AXI4-Lite response ready.
   //read address channel
   input wire [31:0] araddr, // AXI4-Lite read address. The read address gives the address of the first transfer in a read burst transaction.  
   input wire 	     arvalid, // AXI4-Lite read address valid. This signal indicates that the channel is signaling valid read address and control information. 
   output reg 	     arready, // AXI4-Lite response ready. This signal indicates that the slave is ready to accept an address and associated control signals.
   //read data and response channel
   input wire 	     rready, 
   output  [31:0] rdata, // AXI4-Lite read data.
   output  [1:0] rresp, // AXI4-Lite read response.
   output reg 	     rvalid, // AXI4-Lite read valid. This signal indicates that the channel is signaling the required read data.

   input 	     FRAME_START_I,
   output reg 	     h264_ip_en,
   output reg 	     h264_ip_rstn,
   output reg [5:0]  q_factor,
   output reg [5:0]  i_p_frame_gap,
   output [15:0]     h_res,
   output [15:0]     v_res
   );      

   wire 	     mem_wr_valid;
   wire [31:0] 	     mem_wr_addr;
   wire [31:0] 	     mem_wr_data;
   wire [31:0] 	     mem_rd_data;
   wire [31:0] 	     mem_rd_addr;   
   wire [1:0] 	     ctrl_reg;
   wire [1:0] 	     ip_type;
   wire [3:0] 	     in_format;
   
   assign ip_type = 2'h0;

   
   axi4lite_adapter_h264 axi4lite_adapter_h264_inst (.*);
   read_reg_h264 read_reg_h264_inst (.*);
   write_reg_h264 #(.G_HRES(G_HRES), 
		    .G_VRES(G_VRES), 
		    .G_QFACTOR(G_QFACTOR)) write_reg_h264_inst (.*);
   
endmodule // axi4lite_if_h264


// --*************************************************************************************************
// -- File Name                           : axi4lite_adapter_h264.v
// -- Targeted device                     : Microsemi-SoC
// -- Author                              : India Solutions Team
// --
// -- COPYRIGHT 2021 BY MICROSEMI
// -- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS FROM MICROSEMI
// -- CORP. IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM MICROSEMI FOR USE OF THIS
// -- FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND NO BACK-UP OF THE FILE SHOULD BE MADE.
// --
// --*************************************************************************************************

module axi4lite_adapter_h264  
  (
   // Clock and Reset interface----------------------------------------------------
   input wire 	     ACLK_I, // clock
   input wire 	     ARESETN_I, // This active-low reset
   //write address channel
   input wire 	     awvalid, // AXI4-Lite write address valid. This signal indicates that valid write address and control information are available.
   output reg 	     awready, // AXI4-Lite write address ready. This signal indicates that the target is ready to accept an address and associated control signals.
   input wire [31:0] awaddr, // AXI4-Lite write address.
   //write data channel
   input wire [31:0] wdata, // AXI4-Lite write data.
   input wire 	     wvalid, // AXI4-Lite write valid.
   output reg 	     wready, // AXI4-Lite Write ready.
   //write response channel
   output [1:0]      bresp, // AXI4-Lite write response.
   output reg 	     bvalid, // AXI4-Lite write response valid.
   input wire 	     bready, // AXI4-Lite response ready.
   //read address channel
   input wire [31:0] araddr, // AXI4-Lite read address. The read address gives the address of the first transfer in a read burst transaction.  
   input wire 	     arvalid, // AXI4-Lite read address valid. This signal indicates that the channel is signaling valid read address and control information. 
   output reg 	     arready, // AXI4-Lite response ready. This signal indicates that the slave is ready to accept an address and associated control signals.
   //read data and response channel
   input wire 	     rready, 
   output [31:0]     rdata, // AXI4-Lite read data.
   output [1:0]      rresp, // AXI4-Lite read response.
   output reg 	     rvalid, // AXI4-Lite read valid. This signal indicates that the channel is signaling the required read data.
   //Memory interface
   output reg 	     mem_wr_valid,
   output reg [31:0] mem_wr_addr,
   output reg [31:0] mem_wr_data,
   output [31:0]     mem_rd_addr,
   input [31:0]      mem_rd_data
   );      

   reg [31:0] 	     awaddr_reg;
   reg [31:0] 	     araddr_reg;            
   wire 	     raddr_phs_cmp;   

   //------------------------------------------------------------------------------------
   // AXI4 Lite Write Address channel
   //------------------------------------------------------------------------------------   

   ////////////////////////////////////////////////
   // AWREADY generation
   ////////////////////////////////////////////////
   always@(posedge ACLK_I  or negedge ARESETN_I)
     begin
	if(!ARESETN_I)
     	  awready  <= 1'b1;
	else if (bvalid && bready)
          awready  <= 1'b1;
	else if(awvalid && awready)
          awready  <= 1'b0;
     end
   

   ////////////////////////////////////////////////
   // Storing the valid AWADDR 
   ////////////////////////////////////////////////
   always@(posedge ACLK_I or negedge ARESETN_I)
     begin
	if(!ARESETN_I)
          awaddr_reg  <= 'd0;
	else if(awvalid && awready)
          awaddr_reg  <= awaddr;
     end


   //------------------------------------------------------------------------------------
   // AXI4 Lite Write Data channel
   //------------------------------------------------------------------------------------   

   ////////////////////////////////////////////////
   // Generating WREADY
   ////////////////////////////////////////////////
   always@(posedge ACLK_I or negedge ARESETN_I)
     begin
	if(!ARESETN_I)
          wready  <= 1'd0;
	else if (wvalid && wready)
          wready  <= 1'd0;
	else if(awvalid && awready)
          wready  <= 1'd1;
     end


   ////////////////////////////////////////////////
   // Writing the memory with valid data 
   ////////////////////////////////////////////////   
   assign mem_wr_addr = awaddr_reg;
   assign mem_wr_data = wdata;
   assign mem_wr_valid = (wvalid == 1'b1 && wready == 1'b1);


   //------------------------------------------------------------------------------------
   // AXI4 Lite Write Response channel
   //------------------------------------------------------------------------------------   

   ////////////////////////////////////////////////
   // Generating BVALID
   ////////////////////////////////////////////////   
   always@(posedge ACLK_I or negedge ARESETN_I)
     begin
	if(!ARESETN_I)
          bvalid  <= 1'd0;
	else if(bvalid == 1'b1 && bready == 1'b1)
          bvalid  <= 1'd0;
	else if(wvalid == 1'b1 && wready == 1'b1 )
          bvalid  <= 1'b1;
     end

   assign bresp = 'd0; //Giving OK response for all strobe and protection conditions
   
   //------------------------------------------------------------------------------------
   // AXI4 Lite Read Address channel
   //------------------------------------------------------------------------------------   

   ////////////////////////////////////////////////
   // Generating ARREADY
   ////////////////////////////////////////////////      
   always@(posedge ACLK_I or negedge ARESETN_I)
     begin
	if(!ARESETN_I)
          arready  <= 1'd1;
	else if(rvalid && rready)
          arready  <= 1'd1;
	else if(raddr_phs_cmp)
          arready  <= 1'b0;
     end

   assign raddr_phs_cmp = (arvalid && arready); 

   ////////////////////////////////////////////////
   // Registering valid read address
   ////////////////////////////////////////////////         
   always@(posedge ACLK_I or negedge ARESETN_I)
     if(!ARESETN_I)
       araddr_reg <= 'd0;
     else if(arvalid && arready)
       araddr_reg <= araddr; 

   assign mem_rd_addr = araddr_reg; 
   
   //------------------------------------------------------------------------------------
   // AXI4 Lite Read Data channel
   //------------------------------------------------------------------------------------   

   ////////////////////////////////////////////////
   // RVALID generation
   ////////////////////////////////////////////////         
   always@(posedge ACLK_I or negedge ARESETN_I)
     if(!ARESETN_I)
       rvalid <= 'b0;   
     else if(arvalid && arready) 
       rvalid <= 'b1;
     else if(rvalid && rready) //hold rvalid high till rready is asserted
       rvalid <= 'b0;   

   assign rdata = mem_rd_data; //connect the the mem data directly to axi4 lite bus
   assign rresp = 2'h0; //return read OK response
   
endmodule // axi4lite_adapter_h264


// --*************************************************************************************************
// -- File Name                           : write_reg_h264.v
// -- Targeted device                     : Microsemi-SoC
// -- Author                              : India Solutions Team
// --
// -- COPYRIGHT 2021 BY MICROSEMI
// -- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS FROM MICROSEMI
// -- CORP. IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM MICROSEMI FOR USE OF THIS
// -- FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND NO BACK-UP OF THE FILE SHOULD BE MADE.
// --
// --*************************************************************************************************



module write_reg_h264 #(
			parameter G_HRES = 16'h780,
			parameter G_VRES = 16'h430,
			parameter G_QFACTOR = 6'h1E	
			)
   (
    ACLK_I,
    ARESETN_I,

    mem_wr_valid,
    mem_wr_addr,
    mem_wr_data,

    FRAME_START_I,
    h264_ip_en,
    h264_ip_rstn,
    q_factor,
    i_p_frame_gap,
    h_res,
    v_res
    );
   

   // Clock and Reset interface----------------------------------------------------
   input 	     ACLK_I; // clock
   input 	     ARESETN_I; // This active-low reset

   //Memory interface
   input 	     mem_wr_valid;
   input [31:0]      mem_wr_addr;
   input [31:0]      mem_wr_data;
   input 	     FRAME_START_I;
   
   output reg 	     h264_ip_en;
   output 	     h264_ip_rstn;
   output reg [5:0]  q_factor;
   output reg [5:0]  i_p_frame_gap;
   output reg [15:0] h_res;
   output reg [15:0] v_res;   

   reg [1:0] 	     ctrl_reg;
   reg [15:0] 	     h_res_tmp;
   reg [15:0] 	     v_res_tmp;   
   
   assign h264_ip_en = ctrl_reg[0];
   assign h264_ip_rstn = ctrl_reg[1];

   ////////////////////////////////////////////////
   // Update registers at the end of frame
   ////////////////////////////////////////////////
   always@(posedge ACLK_I  or negedge ARESETN_I)
     if(!ARESETN_I) begin
	h_res <= G_HRES;
	v_res <= G_VRES;
     end
     else if (FRAME_START_I)
       begin
	  h_res <= h_res_tmp;
	  v_res <= v_res_tmp;	  
       end

   
   ////////////////////////////////////////////////
   // Write registers
   ////////////////////////////////////////////////
   always@(posedge ACLK_I  or negedge ARESETN_I)
     if(!ARESETN_I) begin
	ctrl_reg <= 'h1;
	q_factor <= G_QFACTOR;
	i_p_frame_gap <= 'h0;
	h_res_tmp <= G_HRES;
	v_res_tmp <= G_VRES;
     end
     else if (mem_wr_valid) 
       case (mem_wr_addr[ADDR_DECODER_WIDTH-1:0])
	 
	 CTRL_REG:
	   ctrl_reg <= mem_wr_data[1:0];

	 Q_FACTOR:
	   q_factor <= mem_wr_data[5:0];

	 I_P_FRAME_GAP:
	   i_p_frame_gap <= mem_wr_data[5:0];
	 
	 H_RES:
	   h_res_tmp <= mem_wr_data[15:0];
	 
	 V_RES:
	   v_res_tmp <= mem_wr_data[15:0];

	 default:
	   ctrl_reg[1:1] <= 'h0;	    
	 
       endcase // case (mem_wr_addr)
     else
       ctrl_reg[1:1] <= 'h0;

endmodule


// --*************************************************************************************************
// -- File Name                           : read_reg_h264.v
// -- Targeted device                     : Microsemi-SoC
// -- Author                              : India Solutions Team
// --
// -- COPYRIGHT 2021 BY MICROSEMI
// -- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS FROM MICROSEMI
// -- CORP. IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM MICROSEMI FOR USE OF THIS
// -- FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND NO BACK-UP OF THE FILE SHOULD BE MADE.
// --
// --*************************************************************************************************

module read_reg_h264 (
		      mem_rd_addr,
		      mem_rd_data,

		      ctrl_reg,
		      ip_type,
		      in_format
		      );
   
   
   //Memory interface
   input [31:0] 	  mem_rd_addr;
   output reg [31:0] 	  mem_rd_data;

   input [1:0] 		  ctrl_reg;   
   input [1:0] 		  ip_type;
   input [3:0] 		  in_format;


   ////////////////////////////////////////////////
   // Read registers based on input address
   ////////////////////////////////////////////////
   always@(mem_rd_addr[ADDR_DECODER_WIDTH-1:0])
     case (mem_rd_addr[ADDR_DECODER_WIDTH-1:0])
       
       IP_VER: begin
	  mem_rd_data[31:24] = 0;	    
	  mem_rd_data[23:16] <= 'h1;
	  mem_rd_data[15:8] <= 'h5;
	  mem_rd_data[7:0] <= 'h0;	    
       end

       CTRL_REG:
	 mem_rd_data <= ctrl_reg;

       IP_TYPE:
	 mem_rd_data <= ip_type;

       IN_FORMAT:
	 mem_rd_data <= in_format;

       default:
	 mem_rd_data <= 32'h0;

     endcase // case (mem_rd_addr)

endmodule


/*************************************************************************************************************************************
 --
 -- File Name    : h264_I_Encoder.v 
 -- Description  : The IP compresses the video as per H.264 standard by using only I frames. 
 The IP expects the input in YUV422 format and implements compression in YUV420 format.

 -- COPYRIGHT 2021 BY MICROSEMI 
 -- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS 
 -- FROM MICROSEMI CORP.  IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM 
 -- MICROSEMI FOR USE OF THIS FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND 
 -- NO BACK-UP OF THE FILE SHOULD BE MADE. 
 --
 --*************************************************************************************************************************************/
`timescale 1ns/1ps
module H264_Iframe_Encoder_top #(
				 parameter G_DW 	  = 8,
				 parameter G_C_TYPE = 1,  // 0 - 400, 1 - 420
				 parameter G_16x16_INTRA_PRED = 1
				 )
   (
    input 	     PIX_CLK,
    input 	     RESET_N,
    input 	     EN_I,
    input [15:0]     VRES_I,
    input [15:0]     HRES_I,
    input [5:0]      QP_I,
    input 	     FRAME_START_I, // must be before frame start
    input 	     DATA_VALID_I,
    input [G_DW-1:0] DATA_Y_I,
    input [G_DW-1:0] DATA_C_I,
    output reg 	     FRAME_START_O,
    output 	     DATA_VALID_O,
    output [15:0]    DATA_O
    );

`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="author-a", author_info="author-a-details"
`pragma protect encrypt_agent="encryptP1735.pl", encrypt_agent_info="Synplify encryption scripts"

`pragma protect key_keyowner="Synplicity", key_keyname="SYNP05_001", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_block
PYoGJ7hZnclIgpohET95yULywieqeyip6U+2CSYpgL5ll7/4CJ0Q6MqgEHW2mu2zjMxzG9G5JEoN
4HwnQIS3EwzNkXq2qvC8mYNNlttKD6Z/UIUXdIkkfQPnWb+W4UrTCnevOHEXVJLyaqp4OBK1ZAdJ
QpldE3dA6gyMIqV8g3ozH/VnZmGp9GEnOFT3qF8+Qp2A4af2eQ0UHo6SLuvHmORsf0Zc52p8MIdx
HWIJN9tt9SUAZ7fTyu1PzOnDdg5qPY8rehU3h1Ejagbv4kLgHcUNUeLPTFy/RSNk0S9abr4NREKS
8eGD1QV+C6BUEJNjtxgN4YnqyPWp7gNCryJ7JA==

`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_block
Xe7/fd7gns/MtXIg1BUoxQi/8zHnQ7gPrvkmmRNFv76gYVVrPhNtZJk0yGarFuSZjNlT91IfcPoO
LfPoNstQd+GdwAnw2C4ujr1bzViuvLxsjMOURczu6/VrV5h24TlKaWN2NNv/VZ3lSYseMURAktSP
g4K2rimmupY+GCN7Dg0=

`pragma protect key_keyowner="Microsemi Corporation", key_keyname="MSC-IP-KEY-RSA", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=960)
`pragma protect key_block
GAJNiAqFgfUNuh2EmxhMrcl9jAZmP5iw7D7cT9b+V3Nt+JyxS4t7OFE8gG5owAEk8SPWzHksL2T/
Nvzuk4xvNcSMqPRXgKOx7XB4ZUDFZ1M7oearK6W1kdLCs7f93WZM9zumZ70DAOw0r9OEUH80na0m
yJg+7SuzO9/SgdXMipsYSsgUMLW7YObeR9MZhoS1uIWb1Cvfm3z4bxLGM0sc1BTeSp3ZB5koN/TP
k00aJt99iQV8JAi6okjPmD1U9xirLi/I46sacPbTrT1u29ZgbXxNSwvXysMG63moADGWynUZaC9t
I5L8MnuRivB7ZRn9N+6QbH6keVbH3wHm8Y+3jdVmv0KwSeq2e1P08DGU4eNbRsW9hUOc985NGodz
tYbvCFF9pyQvzgWMr0JXD8zcOHHOh2yPyH9pxkqaJzhadW+Szaqpb9QxPHArmFQw7ZUcBD1Klesy
7CvRozb2DjpDyx79dTeaEPWE21FRtMfKS1lS3TaEK0YoljZSpK5j5Snlh9rYvL96SBwjVg+PT8t5
vwtl1OJTJ2s/WHZHMaxDPeo5QaAmYvRF6sSkj94ayaRm3Pp7DzAG9Sq+eMLBWeHYkxX01snnHTZz
ywpzK/vxPfzOEXyNIcK2/n4kjDHJGBbD0C7DWzDcDqvK+wt7xwf1pF9DUHBL0NUo3bVvHZdHvm7h
j4wT+8VIYG5EFL2xHcC2l8K01l5QvrBzDAOLKj9JbOpXaCrHHv9KP7f26YRKeZDSMmvj2O/ykGL2
YfCl4OEyTu0vgK+eZ580K8wMEs/S83siQ13ldvbVG9PEleXkzy+WGWVwjzwSVxY65lfXxWJGbbuG
xs43TNe1hhunzlb+HTMk04mfEYibj00UH0XktZzlsrK7RiZUXx5jdQXx3YM8mtEE36NGgEO+dw5u
7EtLF6DNVDhbg1gVZX7kD5EMXa4xUzfBTTDK0CJGEpmdsq4OUYOUR/3lFAU0ogrDqqkZ1kXZTjyJ
+p45NYpqy+Oba1gBRCnKgDG54OeIzLe/bzYXsbdeHcLxN+dHJ64OKm+zn/s6jI5Vhzvp+d92E3FE
IcUk6j7WXbhlyabPLZ0C9tj0QLNlJ/Puy8Y9K9JTlDdXZ7oJT1XEgfLB0FaWgBhQCiAESL/AV9PY
fWieS9NM4c8f61aQs86ch9Dp+gm6ltHVEsNlyQDUqw78pYSTNyIdxaIJcxPmyA+Hdbo5NQGOmvNR
VC38tczndGMd3NLUKitY8BhyuSSK5271L0vhyyDNhN46R9ntdJhv0VSvqhs/km5w

`pragma protect data_keyowner="ip-vendor-a", data_keyname="fpga-ip", data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=583600)
`pragma protect data_block
J03eHscCMGBmJofC52PVsJEWmm84m6dOGNP6TphVadwGOBGAcXpmNXslqxQ4asKK5S9wXmaZNb1f
VW9N+VVBvjoNXbFCV3EdEfj9j9xbaVUOcr8U1ZJqvKg2Ly0skXaDIHzGbueoUSSPwPBcNWfnqw5G
1W7G/SWBaALgygSPeSSmnvgE9Py3xqG5h5xznvUh2vTcDeAmY+C3A9DyWuv6ftG4mWFnk82+sYyy
t1sRN0zksgBLPBoQXjFl7eOBvFNGB5VJYxEtEwKpYBzj6dBhrDkX5rEHa6mMSawICM8bs8Mckgwl
4HLbIy7i0UNoJgVc1GuDJxKty56k4E3FnbRQnG7QrOBP1S/OZ13xmZ4m2zAgKNpRQPPx71Se/Q7t
UTiv0scVrr9JbBxcQZ+n0EdlYYXL9QQijFzgUNOyNjbHOxjKbdtNGkgAlqKnxiFeoQdV/ezkHA9C
7/EQM3Zgl8ZWvq1L0LogMxKP6Hj4LrpcnQI5ZqwlnaCWTNMjW0y1HacwF8TsT7U1xoUfRrb9au3j
ZYVGN23E6YmzY4EE09soGC5ww49w4SdEsRgrkEWiJaWitGekR6FzJxRwtMfwDuALrgME/c4yis1l
q7ywclnxsepRzfeGNdkS8IOxC8HNE5h0l+6d6cxMONqEnhrQuN0ikXiL8vmvtVh7bVIvQRSz/hq6
n+fDtIQC7zQxOFSDyC8DyQjQZt49x0z6OWAIR9/x82qPutGwP4opca3QMS/UvFkKqvUFsHjAXI5B
suLUsu6ewLw7mJA+bX0pfyEJz3Nc4IWBgfm3oZBlVBDv+5dqpBfENVhy1/QTUByljO8cspgbyvbH
KK5TIhW40TWCVnl1iJqji/DUX67y8SzFNMPqB1pPRyV8bJtzvVP8b1DCZtHTK5AFI19eMRCtFu8z
nNnCkkZPAZzP2aiEYimk4XKLrVfQp3/UgvDwGGtkaPbQueROOG8RzS+AbxBT5uq15pQsEkXlWC51
o3jzHldaFhSh9zadbLqecURWMmcEts2TaKAcfMIg35J4s8AL32UjTg/YS4wJb8CAq+0DMzCTGBC5
hYKzgO1sirQp3Im4tclMOqQje5D07FKbcSAMVgzXD2B7l1xTXBiEO62NhpngYGoK4EJCoDw1U2ei
VIwktM0hpTh2E0HxZt6+Z1oV1VUHyLoMba4+gysj8pwPjZqVeXQuEdDbNmx8awkkjbKWbZxfG/wV
Bd+kXK8aDh55EySwA+AFjQwN/6fDBVhnfs6v/2Zxd+/HXCrDHoD7NZaTkNUAMAJBOJwaQj1Fg7fT
ethxn+yvUcYUKdxCkQKtuW6WtfFZaBGJ2DhV+Kh11CEEx1ZyRPWB88cIyKiIwQdC6ldp///Vi2B8
LYV2cZNDIDe/r2NOdk7wLmJwakdMxjMB0zy02jQsZNNq4FB9+TGRhrYumMFmLNpUonyokxlUYfjH
IEWTkhVsH5ND339jNMUdqQs7Fwf7sEVWloo1O0ZdpVouH7JLVOom44XGsGYHThez3VN5awOniEUE
PLG0eyG/BAc8BMxVhnFDsAnaI5pzmlKL9xCVC1P+OWie2x5gzTM8SwsAVE356xwI8DXvZTVXav/J
07i2Jg7Z0+BET2x+tdxHIFrfKQoVV6Y2BkDUrEF2l94oWzwU6g+ONZvUrBz1aiInuLEmRyhVTd9q
5LfU8GS5zFXYAOJVZUWjTe9rXLXzafsn9W5W2NuGFaEzHOZ+vOSQMXjYBf5F0pywzLE6ZX6t0+Rm
BzuoYASQ2uN1D4kI0z+8S4OZ5ACgc8LxjKizhHwLxnzbGV5kM+FfHnxKmF+0jf6cPbuGTJNEjVId
ty/sLCaEWAQ6lMuH9rb3naoS0PiJwfcWOZ2/op3W/QVDWsUkWxBAKG2ECg/3ni75NrR8nixf6GqA
646O71SX6pfOp2xVWV3Uxh4m5V5kQ4BGZc66TQ/DB6wTpc/Z8e8uucPKmRoEJxHrwI/bm9VwelyX
9DD4aheIocYnlkcapx+A5WTkvmfJmZc1/d2oSP8sz9CCupZXkd+g0wSy9rYUVL0VnQ6KyQPPjX9V
9qMW94UyIx9fxs7/RjKzraHjSVPY+GXf0scogi08/aEsba0IczUlcPOEwN8Q4zzEd/9OUl2Sn+nr
yup11Pmo2UmnOjrbx+28RgdGpyzSOUPA1Lo8apoN1P1Qq79r+OwIaMRkOpSnaLsHIZV1bN9glkWS
qtBAKQq8Prz4gqoAAHkjUnFe9f+LDXLlbmHEZUNkF6kargSNFcKxpnoKlR5ckHSJYp//8LSUeI5h
HhXYPti9ChyhCT9fUmPcpMYh44ozb3QDEHLFrCf1cFo03RgCRMsxvHd6oAghdbG96JMSIMYbcMag
8Z6gu9jBrzTJWbRvU2FI7pmin1HsHr/AI8y0DJ52d0e9S/6kZ7QDkvU0Nd/+6Ieq8uwNumep+XCr
Sg7950r3q+eC1dBnvSHQZB7l/kGhkq3CgY76ZUkFqTu6UooRznnKAgjLV5ZZJ5tv+JuWlrPpqZf2
bd8HDVQpm2TPzE28M9FMfGQUamaKuucz0C9pd/X1gaITAfjzNLPvZaDQOSe7U3oM/k8C+j9WHZhE
6idpgz4u+yiWzrhYsznqlhu25KHtFWVnDP84TTJeP2RarVj2arJnQZUeLK9oxJB++S+CsEGEzw/g
k+61qH13xGYR7y11gdzpkmPq/QojLJTK70w+zm93jjtsMmsmA9v9JYNYt1qbMp6R4E19QjWcS/pP
1pCvzun0hfk/W87Vlnj19+RW2dFZKQyKa2WzzwAEAog92KtN9pRA+XN9u5ads5K/lNGV23ySwvSJ
g/Rt5+mDwLSeFcD6e581SOlL9GB2VwSAlTs4G5Eyarropn1eF1idY9yjoeVymd+CM1aYPY22FwCh
FPzlzQDn5Y4BGuzVsm3XYLiIW6cRJYGfb3Jc5bbcT4LdvikGQKAPsmQayCOVYs8NLzSmdEfgA52I
Upk9oceSs85SbF3IxFQGnO/0kWLDefWquFSAU106cOonUzvuJMrSHGWtxJNMg3+4i4jyWOavvArO
cuU6KBmPjFM6XqTvRMfD4i5Vs1ef5lRIhYNrC+ZSM2Tm6uPY5cvKl9Jblunl1OISvjxA/RFU4rp9
4KzcAQv4CpVii4JWDms8MdsoJspbVGlis29vf4eofxy9XscaR0s4Kx+bj+NBRvMUd+YBA4pUrARj
7SEyoQh21k8tOG+WwxF38/GbBvL3SELMI/Xi5Z4xDUVrpU3/7H0n4cwTtiFxmF0nVZ9LSxN0cMYJ
MC14di7cJsYLYCHpKQhU8y130IdDiPHyhjWe1UDi3NREwVryTNPe8OhS8gQkpSzEdY5eetDFFpIP
aczLPvVJk433NibvnTSl3YAKAjb6q/AeOlnmebnbg/r6dZ7A8yxYEM117ZGEj+BSk+9J0ZaNx723
3EN4KaOpc43iY9shLbPMA+i967IHBz+lIlOSaxAJaZoIg4wiT20m+egRZpLEMr4NjIMOaV0ettbh
XFuE6i7tYy9CUsASJ7IdK+O1Qa6npQU3KTplutQ3MtyZJ4g++P329JEEJW+mm9eE9wNcrZZGDYk0
4t4UwPtskf3AQ9eRF+YPxQi+5iq3Ef5XRxI2PkVpx5qpBAEfukBdkPtOt6/v2yssWzBouUd6YZ9A
o4vbbFKqoKRaxkKdPzFliCFfR7dP8IpeZG2iD8bFFYQyNwhAP/s22l36WOvVCCKLJckK3CarWoLw
EJI6tOMCxYAW6SdrAYGnrWhzWn7J21GpRxFeKcyr5i3mh3MKWrGjhhVRt+LrPcbwFZrCyo4+ipaE
x5lclyqvZzkBpWPBM9yJGpSbS/PEwqbRhfVp45DmDsX0z451DnlXpqJwKuhH+s0v38Ih5NzZgZU9
/KBi/a+NhU7Q39KlUbP0YHC/WY4crCWj0xQPmiEIN9uDDzXMey1IatC9FrMylpXMmjrK1vsFzTTQ
4fFLAfsBkyNGulczhjTUZQ/QJMfiqp9t9vTus3iERngRzCR/e8264gK3be7EN43g4ceDoZgacl5Q
lK208sf48Q2y4GwokIwh88C+dIShyDCmGW2Zq7YoS/v313/eh907VchHdDoeJ/OXn6PqBaaO+eS4
+OXnIGN9ixQzTZOH0FnDbWYq0CKCQFP/VG9iuaE+MId10kQ+KFD41RIqBt+75pFchG9rpuhHr/3b
cIe/7iMM7+UuSNckGMQNjDiNu0xQsDPfr+ooLbU/9eWPZr55kOgLxcs0I/J+Ax9uCtVGGhwop+L5
3BrB061+gT47aNsYIXoREeAGouGKOBJl2QtmXyyfXoHgvjekdsroBDb/hRrHi0R+eSPzOVsnnv5I
jQb0SEHsxjUN1PNWpZru7/RQU2I55kO0VDCBoVHs24u/f055Vg7qtFfY1RJvbAUWe07kD0EndVqw
5QVSzYoQaFL251jvW8mrLTvHxDIGx4zaOuD7ZLnyutwOpIA5JmSy4dM3fbS5/Ufz+YVSGajAa85B
AtBF81BwuNLMuTFuY0ozgt1RuCS3gHtSsYF05yeQP4L0Nr3mIMGqJ6yyMHUGR0Nqtc31mvPgYPPb
15a0cDeupB2MvVlbbJ+1nGBREkmdahf2GhpfROwc191dabNs0+kWOHdmobj+0//TT6LjegjRRCfn
N3wwmUMtUORBII86uooGmbHetAaz335/52Gl3yHzadvMtuOC7E2XqZWxzfS2XmhMnzdyiOBSGfAG
8r6UyQ0BkCYrbnv1A2ZyEOyg93I7lJ1I4rVNTQhut/Mpeq8XaxTEHCVaMul0PTwP9CUU94+V7p3P
CzBZpjL4bQqko+3g2cqEPiLJnDz87LfQg7GILBKI7NWcU6/fwi5TcQZezoewVfIN/sBzpy5ZIWzA
+jaRv7tuHRpx+2ecwRaQrhMVweDltkSUlRHJRXyik9HvnY2Xdg1JqANUESclQMvshjHsj7aeZRdN
Qyblk6QK4NIHDA/XR2YhXl2EyFTwGYcKa2DfFl6OYtIbeVPUE/G7VYcz4tpyVx5nF2eHppqTGVYj
r3wkCrOYzD0dYL6jC4cIg1MZ+HvHA6itrRSTyztBWrmPBxV1Q5nZJvEoEVPLoSGi7W34q4wtfnJX
b3d/gwpXkQ+ly3uSjfJZ53PuIEzzfD526Hfex73fZ/8DSiTyW51Pm6zVhCCCPnyjne/b8/uMj/YI
6Db5cbRyDDc/dXzIyZ0aqTdofPZgkED4hkobCeiAV465zoLgzxDli82PRMHV/UHxgEfnnJN/d2CM
rV9fqiDBG5NPto8+7MG3yXDFs7s426XX15Iso0Uz+FDCfd7WTJiFDhrh3az3vaQbyLuts+Ou7UHD
glpFzMjUGEWYy7AJh470d4K4j5kd2bASKa2uC9arV/yoaBNl56t0szb+2hElXmJ8LBjGYBoUEVe6
wb0XEuySUxJdckMMuUxDo0P1fPB67e/Z+oylSMAj1hOfwiCinDZaZGbAbe16/vaLKLknWcVrEN3S
xFwqZpq87rRoLnjLQ2+kYcdBEL8ISjC8PdIEV610KiZ9Uf+8JIqcG8hUU7l8D/T/DkoVyoFLwKyV
nd1tguJXej6qkT/dYkeXCj51WQhM83CKInjOwqo3YqI2m3cvjKJJ5aV88UUZ3K3zfXPPTyfKtbOT
Xp5aEL8+RXwYIfTSixeEjyuNJ4lPF8R/YbFq+JPvRqnZPmVtelNs52G7tMsZmpp+CSBwvUDVbMi7
kxwSo6vN1UsJZBVzYmmmRGyklX12CANXyLm+r2DOsdSzrz/YA8jmL/7fCxrzD6pa3RXDhXt9NWe6
Y73RnigCndoBo7ukSeS7p01wwGJngSMNhVRIcOhW8VvtCYMhvXvJeEVgW4/uv+DQLwpfDrbb/zjX
vaiSf/i/aXoGqKZWA8CnWYK/9ugjZp3zRK4JVCh8JDqc5UwngcjGhHCNoZlNN03HM3L5D8lK/9o/
D8rntTHpsx4RPsphThAFziX/GxX+usNO5l4f+qCoU1MG98AC5q4r37EbPA8BxgZIQzuAateD61wL
DUbT2z4FhOPwIt2Hznwt8/077D+ebueJD8QFRUHzbmoC6Nk/oDlHJ1T23JMSWKXg4Jq8EaLACesR
Lr7hEObPi2JUeaoIpYP/1ggSoMD8qq+vygyb/EZpfmTnD53SWeqKJIDmfTSDyKySJyxv/poJyOkY
iG2HIpR0PJg5QrEOdLLtHkSoawNZ/cBnn8Mse7oCZabJ2fXNYKrGqorhbbbyNRPnEQZjwJWoA41/
0zzc7wjdSdTtBECESVcQVhAh4XGmmejGhzuqRZ9jaUfvAQcvr5R1vauHpV2wD+I+knbvPwJvT+2V
FnTv+Bh3W7QZvukNuIkC8Ugr+A7x6orVbXbJ9Fe6rRsdpNJ2EDbcXt0+WPtPfaYJnUXbmtjJ9eG1
858yoogmbOuScdn+TVexs3fumbaPIBw9rgm33k5iAcPgrilmUuRR1PyvAOtfZjDAv7dd+ESqzFKo
r2jnXlGZOjX59bVw473p33bYk6ye0feTG7zVDuC0xju/faAyUPNM288awLFTqEyqhPBNkWVpG9eh
foJnIlVHAe3ntGG06iMcZmXSEjRRBQ888cs8ldLFmaUJPu0qJo5jJ49KCGpcjmOP9CkM+eYmb0mH
OoeaXT0fpUy/YmFwo1Fol04lyVnBPlq3KbYM7634Tk1AYsXUKIJ3hXmdVipgnqmDL7TjTcDN/Lk2
KBlRM2WvMJ7N8TgSR/804h91kppTEIHCDp9J7z+6eD7KZruUBNhkexCyH4/9RVxtjkfBmZJSq+B4
WcQMTnGfauf5ZjIP7XyUyw0eVAK7mQs1k7HsvfZEJFBoXkTSdnePqepVF5bXLNKo1YtU18ex0U0n
uXePy1OVExmiN4f7+CSDloc8nmIuCNnI++CGWZ5Y/VUXJodEAB2xMSTe6oUIKEsvk7Yp4wKzf4bu
mbHjZmzn5MPTo+Djq7qbc8xQGDylmQg5HjObtyel91BNLrQlW3+75u4MWUK/3KFgJluD1fvM9gYA
WX9lqytw6v0/EZoUUFOTgTcVYzKSdDN15NtVCz7QubMgASmsUFj6PRwwrHJdsCnQs1Auqy5yv/CR
oww48PLqq5UpiD2pgz/O8LP1FG2OWzVBLqztkHoFWnyiNG0JhnLBnJ4d91098EL0pWfN2CgniDoj
91C4b1743HOhiqGVInuDdJe4ykuQHGzt27DuYCwK1EhImemk+nZokqTEAvCJ0zJSLtpqISRMkLuP
uhiVULfbhlxo5ftqb0cyRtNW3oaYcq7mMrtyS2cBc31ViXT+2O7Z5dWnCckO6ImUxeTi318uHNHu
DIVTwjYw5vq+11Nv+2LY2JlyeiC+2XU1EGMOZqwzCZMjKjiYpZG4wxN7XfVoAnzn4JzU/Q6Ux3mW
LJYGvYhYA4yfGqIzDIl5vyohRncgabLKOWjWvOjiDiSbOu85kxoWlqF9bXbdg7aigTeWItPhVKz/
wJtQwopVTD+y5Y1CRKOeJRKOW7c4lUayeOSDLt95aA//By6Tk1+udOm4yKq/yzKq62dnVVLTynX2
LaDId7oOpR5zFwgokBNPpxSvN96KXEvELL/B7OqbQh4EdD8X2m/VoL+Mevzl9IYWaH2wlV95zFqd
ZKh5stYGT4pqqFPO4JrNIGjP+s23elfwnjLot1GOw9DlC7P+yNdnDx46qLxCSyRxoTLMM1bxcUka
Y4zpqmLsWU4Msk5IaBqKFQ2eTAZD/dco89hvdPgBIP319SrQhSoyCXOIFl8by6V7ZLK81L9vtL/B
zDoibLH+aytz63u4dIG5o3AtppoRNHkwrCbsmo3CXxrAdozUqRRZKNGbbVaO1FOS4ffUHTu671+F
+Mbo3IgmBnEbWJF08uaqrdEhQwTMXho7ON5uYrX/otTV8hyGFVwNBijB4w1Ghb3Q5iA4SXTmt6x2
2ccCZ7e9PiQiH36+QE+275WiZ+WMfn3xobK5r5RZQUJZhDycBR5LKT1xCR/DfsVlNQRg1dU4NAv1
L31wn+Z/GNnu2sEDv3jlf5swgIRLQMfdVW58SmVkP/24mQCyHKS0WgTASxjTyLZ9aBliB0B7Vnjs
O7YgLjyU4uHe+ZPbSfWWUvbHmn+5ZloByINX4D020p8R1ux17+VH+1FShcayDkWdmVwOtv2N+lfL
Bmi6miVBW05ACfRjSAkKcVeazoXYwljldSUfZ6wJDt8P0JPVj6GqbOKNfRJjXsFQDvQHEt2D7THU
kJi6iK5N/YovlgnNr91V7bzSqqFSF3jV8fqbjMDmcXKlDXFY3mQx2aVlJMip9qO2ywkDAUV/Efer
nnniU2+kvnO4r6TYXUK5UzcjbIMH5NrHvw5mrS4hKRJrP2A9yLnP/1GA22R07PWdzdMa9b9RwkKk
WheUs3duM5oim4tMc/2F8jl2Pbv0EQQ+ufror73LSagb0WJujzCSf7Foqc7JVoZyFBUC4C0mofp1
LZ7huRvPD3+NzunSedkeH0vDfkcWKtCaYxUn64zGMyMzOzY60DskzbUmBPRooQRNCpiKqQ3UQel6
aPi2VE1fubqN4dPITLg5i/wzPyKITxBmImu28Q291hS3M5M9TjXAXrpKBut3oNkTcITt26DSvx7O
JNMqPebhBrbuNFlJ2y1x/kzdgWXoNsKT9Xf/USYQISHBhQIwpbLeZh2GVNpDShvyB+HDMtyj/msM
FACDxHeMGHuCGA/XPBtnoErQjy82CZ3jg7RjrAsZ2EQhbU3odMcN618h+pTT8VRXiID1G6EncJXn
R57Ufw02G5lut+hy1Du8r7xZP/cdOLQAspWv9dBvKthCBJKY+oNr+JXfpIhdzv0HKXyrqMtlsk+p
7lxvT2G2NpdXu5+OI7RxWcyJ09TeH8STdByTRljlkCeIYqWh5fR7jlnovUIZ4S0IhqnFoejV4u5z
EIeKpStiLQx1JaOPyL0hR1BzDpK2d6Q0+WpRI+gxJ8SbOSuDbgmkUSfINlvvQyKjSkl0SjGHvsoE
5iXOQHSOONoh2VWZ1/Wya2/NDTmbSMONfsih8B3ZvpdCUZyd5xMFys97fNaOuERKlHSuEf5xLCWJ
Pov+EbujWIfefctf9zBrUm52OkkxXros+eIvCFWiiFtts0GtuCOhSnX8GA+H19Y4quGhP1GzNF+Y
MNvGAEtBTBSVOyAPADub21oswy41+vPvzgm5iAT7KOtlIaaTH+BvVlv9ktztWb9lw30yokUF9PN7
5Bb8GM+mgtnNQpBDBh4WWNnpNWtzffGdxvsFFxEcJT357I/Gt0yGnSAOr5sWmqE4RAzwJ4U7cvmk
Cgl6l6ltNo3X7sQMi2EKLvlR3/Z1qj5mVTadP08PgnTT02d9cdUT5PiZWSIMWi2s6gcpvP0xcpPq
5XbikhFPFk4MSs6liJE8qssW4tnLWlxWHnoBjSd2PFR9G9GVUlmIlAnTSRCHIlYJsnVI07IuZC5n
69AYQujfzVWeNdrQuPqbJw1DDl2xwJYtdH71ZAWLth4646wLQk0ZzUWvuuybp/oChisKRrJRa6/4
RTY7E1Nk/uE8eSpvQc1r4ebzdchkmzqYkqKHCKZDyM+JNfDDDXpPAQEiaiImObAauU8TVD/vXyLZ
cgpRCz192L2kswel6rehDhyeAgG4xwq1b/HbnXIsA/5GdRWUDUeOYQ7xRhiy/OC7d8is/NLQqJA2
Xv6Svd6yCLbYyGYy1rxC7DHoIen8OiCL75FzOgUrYRLSYe6jB95MQ5hNTZ4UM6xTEqr+V+YuSG3H
ThYEGp1mfqb7x7p2lfWTZR3GuIwV8jkpYCwyrjHLMVNr584ktohm/zdVUc+orGe/mbVFowkjpGbn
jxeeXS+XHOHem0iM2k0p2qmr9JjDg2uIw7Qm4Gz4ik2xsb9xRrNuvqoEANRrw6jU4WiOR/cWsT8v
/Ib7ZTx/M8Gw70Eea/IQaVUud/dW1cwm6DMMHHxTm3FNABko95yg2znAMve3s6JXaxcERnOaIBkG
LNXsdzWX4tnf1Pp+cRhEuenPHOC/rC4iusS725TjsDoDcR0NFlOPBo3erDQhGPKkz7JGpp/kFjE9
znIO1gGeDY8Ih97zzZDQjAqxKjbW32u0yOPHAwwoGSPk8I83tdcIF6KsKmcv481IeSIbV1qO5MAl
cwLVC7TD3O5Kzkjz7HUk2Ar0qnBMl4RbPG0BusykJMSWTOKEjxRwe/kX60+NQaY3e1CI3T4HlkKi
hD9ICkXylvAGhNIRJCDxUMOe0ztOPV0KIbeS+AlB9gp2Er+OViiMEdcmLUCxPnDOA8m2rBIAHvBM
bwpex28HOO9ueyW5gIN6XKDhA2bnFRGpqxQpPLcx9kVOw+oujiienrX6yxpmcjBjcC7gsh7WS0x5
x5hSw8yamDRwEMoL1p/MrEK6Ezc55mO5hjSbDbzESXlbc1S4wgZ1hF31l55Jq+52s0HUzsMiixCw
wm8RRa2eZNhh6GNlV1Fc/Vs1F4BGaQfW1JZxJR5JP1RPlaIO/fY6RqVcaAHEf1spGPght0XBMCmm
/2BWZ/w2mZhzOkVytzr/2rKYiOEfg8BIHRfOFr9voGs9tKBXmyT4YaT3YluLX4tz8CyPB+LEYJul
IXFLUKeEC+fFqxgfL6BBlt3TVW9P+AKsSecGpECn8feDPEUfN6KOHzrfyFM/+HOB9ok6QX34uX+C
rlcPY4/S/dvrXojZT2VOpXjl9HnIEQkkMGp5hDtjxvE4p6Vp8/rM7LoeF0e8iZsLhvaXwT2d0doa
QhoLjiarl7DotP9gEfwj4Aqva94iAiv/l5hIFmTVG8w9Xt/uTB0XEAPLzskXepg5xKk8ARnw5oJN
bKtejuynspToT0OASXZFOdli+IEze26TvLqz1FPwTfQkAxJbW6w/U5sW5bGoizT7b9NvBRVI8uu/
fbBEnD8Punx1kBnKvsYC4jeHxAiPiWi5GIpaXplE2JbyNopZMd3ctbUGnQXoteYeghB0EyxfPuVJ
tt2GBXFsRMYW8ocwZNNHjds1upgKQt7pb9W8IJssOuPA3cc8tyaEbMsqbSukYT2SR3YLPYEjAQ2N
NUd3WNRk9DA2s1n5XgItKEf6LLAq5N2HiSxDJtugBP10x2gxgAYwF0khqzCFe8q/L7YUX0P+hY62
o3GA8dpgG1dwfmAZH/ewLxC/9NDlSlg3iUZInDhirtNWBfSm6fix2VRHTAYIt7Wcan1Tc5aMSdmS
p5lGNQgR17f0X9y+L5CcZ71W2pDpkqatQ+5ef96uU49oJtqZQHNsD4pJgUP9GrOnEyjZDYutdWZ5
gWuyK5tWdImF+WMCP2qO2BXCM96QZomBooIUtVpiCJf/S9Tdz/qOi2KvPDxNk5lOL+DyadADlwR/
p1DFd+KdKctJGvJfEbDPDYQYmgUAMslsBLXHWSQKa0twzj2aBSMjjfe8nYRVCdSOPOF+0HsgwW5w
FAM+rUwFgFtxxqzhSkTIsG1gd1QyhvZdBbkCB/U337esFYTExndL4nFp3OZuiNNyg9/33NXfRwvq
tBQbIkJoG46Rh8ThVDOskYGgkkikngfjPednM5MqG6reNd3dWZi2LuvQ1HPY4NBWRV3FroiNJrt+
RJDWmn8KkhY8LGYswENKRIt9Rdv9KMNydo4V26kzi1tuSkQGQCq8OdiN9ULepVZEOTu7QMglF5dJ
tst/vDHr56xRIH2Syvth+lGg9UIZyh8+Iv6ogsbv01FCoutpjaXOVYaQmtfMupBCBH69y8nMK4aQ
5PTAnVASEw3fJy+JOGn+LU4BUgMms+OKZHsPT7Fo6+ZhkLkppSWXTddS/H9EuNEshPn9VD3b4iwx
b3hx64yn+HYvtPlotLTdUumXZzUrJN3eK9j5sljyWDxPW5ODTR0e59BX3ZFFwpHIWduX7J+zB5ND
mPVpy5FFowzZ0e7/xpE1YxrbKR/0/J/n/GKp+b4vGNsn+qgbCFC6yZnH6whReqMmBCjKyb5ZYwV6
okeERZVgU4pDW2q2aT/T2MoYdYWaEcqlg+mSyp4i92sYANWr26O/B/2RX20wIchAUsvap3ws0dGz
MwFO1zxff9LpD3pkX+DLzzQqoY9s8P4oDYCQsuesme79TBPTZNsoMZxJSfW7abFyJgwJZiWKu+Zq
WxxEsuA+SUmxze4RkdUzi7mpzwlgLJJvhMHKIyt02S6QhpMT3jo90BJyi8VsXUfwE8RPztD9Z8Nz
Qtzo3Zua4bs57ubtgruQbH1BB/kVUamV/lMYXZXABrUjOKYnHHRXdOBtPLDaVw+1H6TP0ypN7yrD
eyFWDfEna8B+dj7x9KyJel9hTJ+wq1LbMy36rGTGCahGuM+LMLymSmAwuZvyd8jLfmOuNW1Ow7PI
uk/2cAcslHlkG4IjbYpkkemddkANLoOSzw/LxLJWEXTTNuMTkmrp4X9yxecDQVMGE0/hozOPqv2K
OITc6i2YnJX+ZJk5/nnLNYDXcNbkrfoJp6nS7VbNv5fL2U9VGWI99c4ac2JkPOGyI1sQ6iZY9lPv
nFG5Y/akXz5O9s9eETkpwnk95MhbTXuAJ4YgKyeEqsX6gz8C4zg7Al8Y4SC7As/6aXXnvqDDDikO
2s7yQA+lTb0Ht72n8cQ91wpR1E2/cMlq9MpH/78Pf+noB9JsQrtYB2Qne+3pkeAC5Fqj4TFGJ8Hs
N14HFDhqXymQTPrvs3O+9c896QN4ERF96WPFwxp0u9HHSW9hx+ip8Or3DU/jTVZqJug19dl9f/Ld
mnEe4hScoG5jCKLjYKPMaXkhr3LI7guCg5mYoE36IrN51kF8uYPtpelsgaL3ryezZWh4bt76h+Cn
4E26pwYVAoePOqneVdt9fP29yxqv5++A/zgAaWFUogIqyXylMZcwZ2Uu1tLOmV/bZgbMbKHXYz2B
+GPu2ej/8tzEKKP7yeZGIL6GjkRRtAUBgmvGnqE2+aQqEsldCwuw8OtBs6klbiR8Hsl1OVmpZMvQ
TZN0PTDj5EQSitSXdr8imMm2Tc7EVX1AYrNlUIfWSNtKOYyoKtnYOQaWzCrqmAwS9NzQZN2aWJSu
LwH89jo2QaYAJX5SQAZLlBfSBAKcvS+IQmDW+g41EmvFhNHSOpOzeX0E/zwTMjTwrHUJ4Mp0ruQl
jOXMNnrUMNLXKe9iqM0/lDfE+7cFFmtG+BbTkS/yVV5TLVDBZFgR/7pQ0sP5jFcWc0NY6o2kL85N
3qvrJ1F3NBvbDASGabw/wtCejd4qfFvSueq8LYkqa8l9nmmWgdGXTlJsn+MrV4moYUbUvV6WJfiM
LlV89Qfh2hPb2fIz7ZFEngHWD2WlzPSBtOITKHZ/oSJT+Echu2Terzfeu7na6/3d6XLzxrKGblUT
aaHrvJgtfOPe6FIEt98CkBUV/irNiA1UnABw7m0COQRHwVi78MAkKoME7FdUTciSBcMdBEr7Gi7f
Mpul7NG7TTBM+geTva/fmzC/ecVyI7+ncPppwWLowdOc+uWUjXOVpDPs6/U0JdcCsfIamKREKX5B
wMX8sQAbOu3cHTxxwxjIgznYWgOLwjFC79LJqnqHc2839kY1fToAwgqNw6bZFZP5ajmQroEuj6Lb
ifVsfZIk2bFwo81OSUPqJHQBhI1k0+phHIXCa2GkWVP0CFc8sCZ5NK7L/nYZO0OzXMtml1yR4Y5P
XWkyk/zSHwUNbPyr/ya7DhBMbcw3BbeW7okEAkqA50kgPvCKVUYDdm8mYTzWbV79R3YVpstF/KwD
pHMC5Gy3WfSifx+DVcQ9Fi2762j0tdd9vZV/9gr/2kfnNeZbns3cjvr6i2G5kfP2w3UmMB8NIQI8
Kl0uFPmRZxsWnrmUue4R3kDb/aSm6otlrZcvyNBbsaJpMEu9RJvInPOAnsFXxKfiS02uB8xtO/5b
sKfAWhhZhYdqKCK/wUSR/qzr8Eic7tSQEZz3XNyCICGzQ3/1yLWPXCRjsOPxavzOIIcsjqjy7wlO
EkMAhEUHe/itF00M6o8bNGk25qvdyJT0Bv84EcqqBQ3p8zkAkF+DpJEE+BfO8KhSjXxy9bL+U3IX
GpZ73fOevnooRQqJm8zdNmUAAyQgVX6UYP8xhnNXHmqRME03MQhpTU6XEh/eZh89QX/BJxASitir
L/2U2jSL80Q5Vu0wFhBp5oB3lCFErPEGuV5AC1SIIWe+EeZQUq79HbLt+vEVsbPjCpCVBZObvbfT
PKGtSP76GhK17N1Ui3qZSYTIggx+Booyb6UXS7bR38BgP2JOqpgftvdFZJ7jPa7PCRQg1Iwy6d97
5rq3aH7n9n2/EaQQtCKX0nx9WgTuMl6DSn20KGJrx4a6PYi3L90dqEru/wCo1Ez+0XbeR9038Ps6
CuzOgaSIrWuW83FkiR7MEcaV2ych2jPV11lBE6SCdh1muCIFpWu1cGpFDp0JGpurr0bB5v3Wf2cD
uG5Pij+IVgkt7xO0/XVHv9hMqA9sekad4C6aaxY8yrK4vWrKvFT/qtCZPYrer5IcMOvQ2FAcOOZV
9Ka5GyQ6SXz8GTUnJycVO6sljtzEw4O2QzvN2hPTdtHuNI2SG1Ze7kxoTkE55mQTGMpdNvEdJV85
hndpjW+3WiYBrS67LtK7olSJApBwZib0AeVHO4ZDLO+0e8Kg8MXKR5iN8m5t3c+XDVoLFtbwgj+e
tq1hrT0KxxYc8kzlP1CoKE/bQjxWylB5j2+QVB+St2dgk7ghQZLlp2ODhyuhiceKTea7E8j9WM/Q
QE/HkfFrgSNCfytd5V6TogUe7p+VPY13yFl6CWAWKHJOWtmzeBRZy2usBhbuCnTeVbB5Q1Mgd2my
FFC3gG3YCywm+6hAyTiHLN9t7d60oedjoLUFUfXRnrDZ5+0iqPdPFCngqokxmk/3kdvkyVjJlgPG
0zPwC8plrfRBZLoyYE1t7UvKKoQg72jkJivyZq2rHL2Tl1/Dv/WIlUJpubJCBZ1Y1H0cZAlZOwMB
NqljfHfWQBYkuV1iAl780mewtCPjuHGzA8jv5tsoUMbfuT1bo8ZHEm6Aag1niylt/FoOEe7B7m5M
F/2xnJRetTxAVGB7Im/OyXWeiUz5j1r9otUX4Z3AxI/xykJDvXlYV6hi7vOevFWe2BFS3Z240zap
6hX2aA5Bsf9+nACkryA8p14nhm1OILiQav5DiLNHgEOUqmEOeqFKwy9wYh3qBt1jLGY+NjMtv0Sc
vgU5ZPaD39NBHMACdMriwOvfoHg4uSEwzjc/t6xXt55IHEePxaUvszdJlMfxUzEubNFt5jtFFZja
JoIxls17fsuhYi1xlyUnfx14iyid6U+5r/PNi05iVjuXLA5Mzf0Jxf4a9NRd6W34oudcBLd5x9AJ
fR+Vb2j0sXbUBMovAOIlh9sTGjur9mlsA0fqNrkR+cHBwdrT0QXs2En1QmWFIY4BiC2s2RVC4qTD
9dEgTbSb2jQA1q8MCXeKHA7qInRVKy4I1Zm4Mf9Aa8aCpsd8ny5rcoKuFROE+4nbl7jk7TXspkAB
hbcYvL34mmQ2JAPeW+46U4/iR5D0NXCcuR/TzpQj2L523sEHYqgPawcUIxCTjO9SYfnRize0VVDG
1nyWv+hnJJcKXEU5mF1gTBmsIz4qGi1vjtChppWqD/3257G11xAXJO8Fq2TzQL6SpqrjINoU2yEf
5sSgFKnf9/7oH9FQkrlcsKVzlqELx9Fb6M5BETjRCJuq6EuKT5oB4QFi+DoElKEroxLhYXbaFPTl
INNdpO8AOVcX1tsavMZA9CjDvJeaMXiOVHfXyiCTjq9+7U0R6SM5HAy/FDyupF+8F2geuWDDUgCR
/StozbUbOVLlxHFblic85qznrNexu8RCurYj8mBnKSNOT0fVozZXKw27j6vbObXYwlqtvPJeNeJ/
XntZ/nJhiEgPMGAk6V5auL3J6cMLP/HcQh1wKsVX3EJjSmV9xjrBJSbcAGSKMLIWsoMacWxHyufK
XWrAwVcgE+PWXru8NFjavkNmzHPQPU50g8V0nSMWQ4pdMZSQsZc8GHnISck6vImtNOWzNaKoI2A4
mNFa32w80qv1nYHk+yHvjcHMmVEASQzEZYDi8FbLRgO2SkXct2LVOXpSlFfMUQkoL/4F/VBG2S8K
9sN+gwaQhtyyTyDvXV+LftRXns0ZQlaifx02N/1SCgPkJZnejBQvWSUQIldlO63p8IPzimkfEA02
aoB4gJgbxpAGrYnr3OFdQBHw+mB/O++e744LyEsmfdluRjfMQ5eKWFRLM7sotezfzKLNSWwZ5xmy
kCReQgPhjiLhNClKhO9LRXJSMJFBdGbovCvGmqvgbQ8Sjqux0YPs7pkO5RSJ2H8BpDMsN2HTf1u9
ThiEwC9hl33i36tgu6DCgGfyLb9agXCKv9R7oqbSWl1G4MiaDwZ/jhM0wL647GUwngpPr6FumHCH
8WP4WzIe6ViYPji5GAFAjO8D2VuMe7MLLvxfHZBESKiE3MR61r7Wz6rthmof/3InQIy2oyrBaToZ
ggcdtFWEP0Qaq5idDqKsgLRt//jjP6ndPNnmYxpuJev4jYijitfbaHrkEhHb5DuEtLtMv/vVO+kp
q44Ss5cj6A70boKuu+7oB1Y1cR7eDr92TY0Rl5CZc9kQR4xmqeUayMiVPz2af/sGb1OCyvVjpgLt
43MH0W3lMm7oDH6hfzJKntXN7whoF8VW6XXENHlB4dsYrAD6qIor8TtWTYKByDN62ApltoRkDfc3
Th2rYMXN6b8DT36mFsXXKQh6EKKoTZOfJ5y3zPdo/yvzBpZUxB7Cm755fF3x59uS4qoEXs9Y5Or+
0ThowJa8no5Rotb+W+Y8mhw96Y1CWsr2xUPt5x0YQVMn9nzE2BB7IzKJ9WNCFy0BxnkGbQPIseUD
dDZ7FfJAj6dKrW3YrushdctNJLTfvE6xwxN6FdQf76wYj4WiC5EJvh12h6QpnWzHCQ7YM5IuWsyQ
Dpjt+GY5KQ+wVjmYLQbv8BTZ/MkH9s2y2Kz9nhNdWmVy6pv9QeodjPbLDvSFp1hXI3k2O6KjR7yB
niqzOdddL8ZJR18MdqicMSu//W4Cdav+zDpYYQe1YClZWGrGwkIofZJnkKYSVEoAGIrSqj+iLSF5
xLwDuDgCJALaMr6oYvW+TgXtSrJvSwZJREs8G5fqWE9AWIWufGhg/ZGKZqE3Ys+6vyXKztAZrzoe
Eluf9++/JppFw4T8QLriZxYt1rHnYtAJK3ZyG7JxAZbnld4MTYcg3n7D+ZOrG6T7wyrlsZAb18XC
Rb24R3+zyLZcUS/n5aKRBHnFiAH4wzcY/DhF3bQtoaR9TiqvJI8AlEtV1FZ7fj3HhZLn2WNehTfG
Mr+r7TDB6IHtnIVfHsUUOk2WTar9iUpHJfSa428qXgXjr9NHR5IIyYp3WeT7/n7vqfq0xSZWoh2O
WxoqGdYe7I1MMq2VKu9pTBMt/ZAHAPe4XOTr6pj1UahUnXDHioNAne7KY+gJ5dhQKkSy9stHUmYw
sTKMfwZrlgjl+P+cKbZLd+plZM9en/kBXCwY0F5zhAk7MX1K64fpcY0CJLED7oLuBACV/iTAplQ/
0H0pK6ky7sHaKmxJHe7xs1hyq+vbO1EhtSEPau6NRj7yUZlVVwTv3wWKdq6m6mfg4mNvIy1B7xPD
STImVNZqq0jfj2CEcJfQmuiWUVdCGro1yNmLrvZFlaTdHopX8YufS8Bx1p0AKtbf5WUopMlBA0Bi
xnkWzZGORNLn6gRoyRaKHE9LOUfjAqfAGcpzTRiHPJOxeRKXxDWVG5OUMR4ejU3wKAuizIZxu1Wz
PSb1RQ2bXkKwvTpxGyTUcwG3sWz4AeQwRT8asku7zzW0dLrM6txVaA5TaJo+HgBYhOsMpLQYN81N
b9dD+P+Xl3/nC9r8a6uRQQDarVKdGOJdxdoUCG2AdWt+PxqTGGhgzmShzNlKBPAQoVD7t73VsTPM
EYQUGVydOBv4re+fnzTJ0JRWGYXiueZ9x3/siAWrjLRjrfCTDeg8GzXCCx5PP4U2/BoxD37cqxTE
pJS1AjENRYVUMf93driBsp47qq/aGQviZ6YZs2bj6yxt3wXrFL9mcwApPaqs7qo2PzWUR4Sfgbpi
1XUpkJF3QWd8sMiPEZfBlaaeUwWeMI3EPT8kbE5RW2xJqchmCBwDxmvrqfgGDpZiEYhm3iqd/xIk
FhsEk2YjgzEozwQzkEJFijXheLRKl/weybERw94KRpTYUYKVbRT9wDYUSZ9+f0MKv+q2Jc24F0YR
TOXhwbbnXXUgGhIFZoHJ/cwPNfWKb6oVHCfUVPKGKfE/iwbg5LyICz/ZZOgGo0L6pbdsKAHlduWo
9+EtlkSPSovWS6VPSyvCVg5R6IhAGLD0GkLBp2dOyR0CCj2k1WSny2X8yzC0vSsrZKuoU60e0lIG
8Ep3sUWnFOFCUlPO9KBY5HhxyIxpjNrJX7T2P8D4R15Ioxlto7ts3mSpWfmOSTRt0tx4xFb/yIz5
BXM0YDK0LLszmh9irg3rkj/tcqBdWJNceIbJZoRvf8e21WCE1pSO7WaTmWLfTRGX+54ZcKLVAln+
yuN2gdLztD9AeFtOOT+64BRqRRC1BI5UdbSFSHLnaT2zRX6RENRE+t66kYhMzT6SD0XWhcs4B1sw
N1vP6mSs1ehcv5s9atAKyqVKLzlbwB5WEU66MdKryCkfEli3FyX+h/p6CV0klnS1yI4tAda+UEQF
RG6Cb2eWtM13eeWMWo7LxOPpl2nAqNm4BYWC5lnWcXTuUK1VeZ6iRwG/QN+l7Vv//PvhfrIJJ6r2
d0YZUBoOFXTkjubgjWOAA6d1uLVPX4stijITyfytKlmWiIPOsUPeWCgvZ1F9prLYUeSCoEVt1MSL
2clAS6EWqsmO63te4rz+FLtghxcFL6eAd44ScQ30hW1xdgOtJQAgERCQjpQQlnOnMLhD0wbGzCVR
/Ib22e2gT44fZmS8o9goyCp821LRNmqqYVs/fy6n5YD0l+xVxqFFfs9tcW7rjUJNzSCkwgCLBp7P
fg+8DYkbB1LbhOn+nW/fB9xvAeT8wSdVka/1VMXRdCh05COmWFO62xXbag4DsXhjj0Czq6Bnd2as
RBpvxv75o0oerMe64wevcl+nhO6HfPmofilmVqharEZAuX0MMQe/isokwgdgvrU9tpaWL7k2QqMf
ZDK7FjNBwe/XQRtOZzVHNmoHMUHms4HDRtOu19zkOyJxjIaCStI8REhixPmehWUXvNYZ8WTQogcT
TeQQJVjkP/MzYbD3sD/TvCw4eXLpfzazFrhB8hd2/dtKeYZXGf62jUSAoETiflySZ3GlBzbp/dJP
H0m5w+ihGMPICs5zL9bcKkincw5g3iuKGIVawv6g+UMVeSbXvD/H+heqVUeQXBt4hccxnqaZ9Uaa
Xh8Ql93LfdOKcXBc+7dE8E20Fis1mUN5xGtmChloTL3TY1yFdfRMddycuV6Axqkt3LdEfFJVr2Pv
snQU1xwKirvMDPZ3SJiH7mUVSjG67nCvwFC4q1JZV5iQ4ZijnUkvfFiX/URlx12jp9h7LNqhFXOT
1pLmRIo+T2Uo4bHah44w/rtEPJhAGEp+H7+36ki1yc6u8TVdwhSPdjsbdRE69H6PlR1+lcXyQJzF
CcaLjYXIY0zhhdgMn9Dbx8OKpKwsTR1kwPu9fmJLfxBu34nWfr/TuyYQfVoOJSU+j2ugjHk81Ks6
SNqFKmpCAEK0DZXG+q+kERRREGtLtkgCF0hF2uZd/evkAdRicq7DPFXQIndrokdWQlfH8/KWBPhd
Q8UXPjN7ciukQjybTNFJDHW3ZY7YNlpx0UF310K/P9V3siX2ny9wZp6twYIdUuB1ptTA/7XPNgMz
5KPs9RC2XuKhMs4HmY8BFWu3F2NTKqq+F56M4oMe0RU2cvZsotX+BAEt5snqs3bywN12sQDHEFN5
nRakqtANYpUnqnzHcj3DuRK4/2tBbOyUGaKNiUKYGMMoINR1wU1OryjCitkqtQU/aCsYMri/1nXn
qASnMNkAYz9WzUB+upqwcOcMLlZY310hqUFDo1ZObmRv1w66G5BYwS1sYyok59Iaix7a0XrcOYf3
Q5UmEQomwTFhHvJ0CALvYU3NKWFLvqLrgkvc4e77EeLIY7exOCp8o1KOu/lMRT2CFyvwFGSYdmZC
i4j+UQ0afES3WKUwgCIts8odkL7Up0/pdxDnhixI51GbqFPLvp2bgY020MQQkBxfhJXFm51j17mo
wlacA0SYoBiX8szlTWBTUMznNDV+gXUm7ZCQU4tQLXZjZkJAPHlEfzl4rcdpPRHGvdorAKzXNNSK
nUO+mkpJuF2z0t6hYmylJyHikMWOQOTFnmV0fYYS/O41T0NxhIqil93sN3yAr1taZY/Us3VlvyBC
YxK2LPaQZlf6YiPC0B/sRXooIijZ0ZQlTghl7LUYGzW8quoq2ggDL7gs6bwfacA4JEeh9tV8GnFY
VjYZ5Id4iP9G+4eh9dPbnsfh54GLzf5Q+nJj07k3dO2WsLOSzt0MbxCa6LeMRNz8jk+dWof7VFuI
7Q853QntFhZHqkoMbORjv973aK+FMNvVXm01BcVlhrLOpkirhvqIQXRbeS1dOF/44fDiyDIn2cPr
4UIR7Vnc8VFq+k6RRQthqK8iwuYEPPnnJt9x01nsJQeReCdKDjSVkKktGLQ9GvUePZJx25OvQIzI
hYIgQ8NUhnWuTUtcNHcS6v8QecjNyvzHxrD9e2LzYnxmCdLBYDiI/32Jt3Jf9Quh0vHieblfyABB
UcOSO/XNeJfsaM79e81QWfwX3ZvKEPEPEO6owkAyUs9C/R0lY0jzjmoNT5VIexJtP/bKfNeZnUaF
YYnlWO6bbT4QTrzWqlTWGEGJQNML7BneTlnmXimkQnUd0A2FJUb09FpPTrQ6uih26XuUP5cDfi1/
AVQCvPZAKqd9nolfExcMT6idw273j9jFidExBJEJpEPoxUUVanPH72UyyyKLfjGBvIQSQuuxGiZs
8JoOAAlLurkP9GeHkhuzvgfh1CDRNUmEd8ZE4b/YDr45KFCTbVWykSnC3n4HH+gU/QGvHrTPKtl1
6xOSU30rjBU/qV1lYctEPqcT2nWEj8Mc1hJ3n+5Jp++N8FhrUacOTADkMJlTUHihVoBLAa/PWZFy
xVq/qZvLcdLe4HgNJkW+FMQ6fca1LFgzEGsIXqvvip9P0GUAU1A6G1/AvYgWiHJB7AoV9SVH1YiM
y8Qf7puRHQjW8UIN4zzVoA32bLCMEd9cuQyc41mvR9UEUUIQ56rBmKmb4LSviOtLy9QRmhgDTYdl
aGJhoY5Kl8yQAeIrltKlBzvahExCWEg3Tu3nWzrwfaNkeUKoxfL0M/Qiz1aTmSIttSYMpY/snGYe
Tc4G8Sn0jNksUvzFEtO8rBrECKoLL/jhrqbPd0tTegdtdVgehPUO5g0ycweao6WLjhVllc1gsPwv
xUjnq8WTnezqZRsLXZypmTVl+Gbg7HX/6ot9FyVqhfCudwej74gATNqNv979pjwiykQNWkxp1nqk
2efCgkaRvSkdbXD0hKAs3aJ4KvVYndmMRfbFyCCW267atJCYrnLXf2yHXjQazTGhxw9zKjZaWUM1
13EPorSVVoGQQfyB3M23VSdIU7BGxGOHCg8cI6gEqVEY97Evmmh09Pv8ysXmIp+nGa6lPEqPqk0/
IwPhsyfYYj3u1QlUwa1pGLC0My9lvF/UR70sPqLHP9FRdXv0seqhoeCPZMLT8gitwGFR1DVWl0tq
AxoCJuYGDrhjzfDSI58ssse2ryt4xz7JlMKE3SDR765jFxclEwDoaPzMBrJFe78OQ4IwS7qQlvZ4
KHcxmovLumDcY2hSAl3qfPtL+CZzcvTcDYJNVpMDzZcGHGixRDaH8lY2r/i6S8X2Gt+nT1otNAu2
ViuPyzoW9xP5a47lyf4sdlBLFwtob8znbslb+yofYHW1QFXX8DU6KcWdjqUL9myGsKnPkYAVsslW
Mi+nuMtp5wPm8MruRbQdLXa1zqfoHH0l7+GRVvnm7gSj5eFrEH7X3i/0cRftUwiSaXYiqjVCfcQR
G+WAPGCPrif5z+dTZlxovMTQkwXsSFknyA/Cl65mY+GXil1XaBHbIgRdx+J37CuaxV3jO/VQI5a7
q/5qXx6V2dBRdt6bfyDJYUbGZs9lGe4vcd5mpmAuUXO8PwbJDi0kV2hMR/wazpBxIKncOuKc/Cpy
vq3gjcOWa2+zWm0UWJELizgBg9B2mHKBWgShZWmyYSY2vTCsfiHCBkbGhndoJXWorizlEo4+x+bo
uAW0ditnKeVTxW+6jSx1FD8bF2mLc1cX14EcI/dlT1oQ01Ucpt1pNSdz+Vv6Jie9XoZhU1q6MGGv
mJsvx7sjb+nHGuwLQUmwiH9VA6MTI+Y1YBsNiO/xfqPcGLpV3AmMoBrdpYOxlPjWoGgBjBofhXiV
YoGz/zla0kV0AMNUiWH9n70dgKROBRmxXHocNAWlnY4nho769bxbyw2acoVVAZThrjhJzemhbyyN
X317DqiSbPWOwiEM1YwmuAmrwdfwBMXRkiKiTMfbTsq21CsMvNZhWo18L6bRo0/Dp2H2qkTDQ3gA
VAvEbEIUpxYQFSKHWwd3PZ+5aZa7ogI+2e+FUGzIkH+nYoFG4KaISLi/3sY0JzCvyvM7Of78xUlw
WTznsLuif7YRKs3G+Ahg+PRAfu2wGQjetz88mGYMWld7FwJ4EO4ywEwg/AZk2TzLG391RlfopX/x
XKjsZrqUbonATX9dih539kOh9hkmakmP9Oew3Q2kMmaRzPCQNocPSEH5VroGqkSd1yWdfXJTf0M2
JOYLtiso8TNCYZesUnOE7qlv8FN0VKjzap0BzX2VssQzA38lRPKLpBoMB39wk8PnWfB6ihH5+e3A
mnPUjTcTv/9bn20vIs1s+HyRrynRl288pu5jJP5emoX1/wEPgiRaDj0gCn9L4fxrPAaGybXtQtID
G7uf/9gYpcrPcYki7p3N4/iJlU1/dUT2j9wbq1/7j44/HIXf5CE0n+Bd2srWGiz+nLJxExentJwT
0fSUuMi1AjvhrcYoFdod9yFyPOniRawOE617n0Yk8AH9aWAhvXjvUTmQlPBhSqamy/05/depyQ5X
xJKZJy7GDr4/n6XX2Rfy7aUIMKQz0kj21CFRtTqkTfJDFEy2YGNpFt/bYQANQjdrMsJyHvU2e0fp
EnLcOH/Hmc89rSrxv0kx2vkTehK5nGAp5SS64Vocy5tBAdjd6BqgMh2IJFI1kDeEFhgIx8wNmbNZ
KfWP8cOBkU6r8mK/v9UyBGB/k4iMZGNDcNNKXy8F7IsTMMTNS6dNHZnvUdq4kZmNu8rqPgI1lwVV
AswPtM/IxaMG68A9soYsYndP2pT4P4sb/KLA09+Grz4BMy3z5jzdPB/HSPnnvpVakh6C/aM270x7
2M5QZSErecTPOqO/hlA7iRWf5Ju8OKJMSAuVlPPgJOL4ZxGSqR6wqVzalIpxYFz+q/oGD7g+tXd2
lKf7sLU+pgczbH6nCjvpWxMbp/tLPmLWEQYIKz42c2hChsKEeU0TkwCLXxWOFJFUTN2lXCIbd3yM
cH1IHbPmhKWa5q2F1UFzZAWL7y0539kBQTveALp0RxMRveUDagAV1kkljj/4/ufs1wGEustm+pRa
nT8yc8kSPpBmvHKyDkTN0AIEBi+tGcamcI+pBj/v4UER9V/7YEzLo2bVANzxI9lZ+iDKSnvhSexY
XGCy7WU4w/dwTgvAwWco5hhLZHWP6wIGw5QLcVJt7CuybjxTpIgr4GaIC6SgutakGzEp9ZuYOYTC
bj5ZaXHWqakFlHzc/2NIxWNgZMvve3MlF80QnxipSPwCUiheCHTOwYUxCDXaJ0fNTX8KWLZemHok
5olDJE5ysXNOuCF+jvXgolNrR6g+6dt34CYHcoWGbyqRThG7o5LNBClRS4W4kJVMtZF4MnC8oS45
AREDHd119U5PfMsLBjfQtzSfVQKjHXUZ9CMEHd9//8SZi6xD61qJkT/D0OW0eBuMqxh0TdjDk3pF
YXtdioItOhQ1rJJhTLnoQdeRcIzOl7sirrwgr3Re9mgmeDK2I1HJkTBf81lKnGZIgsevBgVna+x+
8JONoBMORoay6RsWV8C7K181TKncNTFQRj8XRtDzVzXGP26wIG8qsngRTmtqDD9D+l1edjPt9PTq
7Z4B6iVYtiF+G/icBiCa76LM5s78Q5jHIhzT6zUTzl+Ul9Ztt8Aw0AKvAwUN+2rA871cotYLoZWv
4E8aeQed8U622QQgKRMkaTCbYrwIqRucqOcfnRFMLPJ2nwTrgGEm19xos/40+p28Anzvc6vg/z3F
ftmOsZBvjSKSktmsD11cre/Bwc9GF3/TFHJhitDWOWy4zoJQyXqayiRmC4nLHtQCOlprN1fAg3F/
6Jk02CTOwvzPm4yVrv1I4Wq4nOf4EziEe4Z2fgZoP7zf74Yy4cOlsPPmerIrhizEtfukxB2FiJWe
4kb9AN5dfUWinH4XryKpxbHNQE2nKF0TCTuM/k4tBPVpPFF//DaVCzHS8IXGwwOrR/uQzBdxYtsn
JnqOY2WHe4my6dsKVOY9iiFz119Q43vpoLRi6qZEfv1E16iomV30VShAN+IhASSEaHdurKLrhcS5
vnfGGwYSaexph5MCGkpcaD28wq8b4tngREz9S0NXinOn8DuAdJccnuLS63HA1cXMoAi/Y/ZQMmqU
vAipGtqbpWEqKxkxFo67VMFBle/++hkiWBBtw0w7RbQOU/OAMXWFM42ZXQ77Jl0WmRfoJpHriFCY
J9GIttRVFwzbHpnv3wFp9mmPRMOnolZtxKOnqNqhNBVxJVut8Cu2iKvRAR4o1h0iSM5TCnIwOcQ4
qTHkty16BMDpjS2iuNzmlYkcQbdi+ucOxRmkxwuLe2P/ywWKgF0oSuNjma1qdsH1rYJSuyvyFKFy
fSRj97xKArF3/CnzKsi/LEUoI76QsiUGWg2Iw6oNHNOIArDxVZqVvP6u3OJJ9YbPHYsim8jIGk90
UoybzlKfjkBVPJFnNdgHdY88y3d8+qu2fXcTnY6YTgRtpn/De1q4oDDHIHNizw5KhNZXmcmn11j3
NaHU0dIvqB5cgZZ7VsvF8nUAFYskZNIP1ehtrWVgwrwMAzp2SELtKS33TqFx02Gr4z5b2gj3pfHF
OXnKJQQFE7o4L4nZ8Y5e2rxHdW9GW1nagowhM1G89VdBy2WeHtv5+nNolzRWMJbLQHxNv6i64uGG
zayDBE1zX9jtIwNciTZVGv0qozCb07adpd4yTu6b/Xmk7XEOsRKthy/W+bUPjVeHdXE9ot3LYAfs
fU9wrDiZpANIavG9ryxzQs3mfntaubOmnwIeo82uMNld3cS+yAjyy3CvPA2HVePTIzagotLm5EGv
NTri5mfE17Xq4NZjgd0VEMCHXU+bLdQXviv+mrKFP4yIWdiQ42TVsxNVV5U8f+xjZih3rDxYCAFF
PiZd/Kb/U7rSTvcOdwBk7G3RH9k7cH6CFjT508h6VrD1VXud22mpQGAe476n6NviTkywuqm0+PNg
5OSWIfGsSyqgX9dlCt6TPMxrXg2Odwt3pg81EI8jdB2Qge8k2cPGgBJtOXeGGIPYGmkUiB5q6Gum
bmQNkBxozfyZVSNsOcXRh+YJttedTzLqCulS7OHTh5Gy6zaq9vV2pNIirdKVepe+sQFem7P5mG9r
VHt8wQtO+7T0VypbWshJQHt63BSv79kJhjczcJ+3eXI7AVLfjSCL6DzUSPEYpHN2ByxjNtHNRbMh
ucapil8+NBqdKNekmp+nhw/6BtNR9qRjD0CCwPHLsa/SpvhXkipOWUwFYPQLWdVzOhtqF3EKgjSl
OrhWeuVbvtSMR1KwRE9sOpwyeHV7nyopxG2sILeDEtGHZX07pceQE4kBnqnbN4G195Cm9XEesQxJ
wm6Z3tq/Y2Lb30KxnSR1DCK4iLKjkf9dcFBYkiWuh/4iYMGYyrSS7keooN09q+WFyPKvvIyYqex5
TgiCMYy0855+w2/mWoqrLLLIIVqfOYyxl4dfp2UyqiisKHxk6I8+7vSDoQS9BREAPcem1qXsN+NS
hoeuH6mHR6aXjBsuYu46/284bmJyP0E/YT6mkXGHf6HU+xUaFTiYu0Gd70L/bWj/1lRbRk0lfTAQ
/YA1hLOsjuZn10P0Y2EKcWDZotxMESq5j4gwcBQhEjrktwaNPBuSN/63+f+u/qbcii37t8JSl2gQ
FJQuacvWQO8CtvgQMpmXVgrC0+bfcR4tUPjOFfEUlLr2uFChDxLTZKtAl/cGgth+avfFkng5y3Na
aPuP0yq2BuI+hMy8mgEeRq7Qvm3/XnF3r+4IO3dGANIh83icXsQkysGgfu1jzowsaQD6sC1q1p5U
b7yyFCvSV71z/atpu2VHL3H4GEVrbu3h7U8lqG1uZYESKsECut9jsnCowO7GrgBV5PmxWmWF/olL
ZstbgqKIs9lgRdzA027j1pq3A0tTh5R6ShlLuvQMlC/PBz32RE33g4vcyejkZGWBFnpz/vQiqoKo
ASWOhvdAuKZ/3/JMnN7yDKKrAmCDfo0dtuusS5h7vSW9fhu3VHhV2Pdg2Z1+wCij0caET4BTmwMg
tRt2TrMjzP/GhTiqesqlZdDadS5sdy2tm3zFQ5pJ+bJOIHSlZMwP/2BVSUEFKmEdTcW4t/ZvhzF4
FFCBHCSX9cc+QkKcE6PSZGOPClCLmYKwJnQ6aLGjAmh22jBpRI6Y/cnlbnX1jy7M8cJkzLUbh9b/
LQEKUj6cbGXbTEbndXiBmpM1+FlvCGwaimgge8Fc5v0YoSKrjuA7+w5I6iA9PdjV8DcNZGuq9iaD
yrOpWQfjaRJmNpYgGU0WJ3Umn/Iyf8MRnGP8xWBBW7q6UtNltJCgWFHjh6YoM6ECUeboHzydxrZq
8ngt1G3EiiAaHdP+GQo0y62wfhNxUvy6B5fhZFt80KzzHP2j8lnA1VV+8uhWlX9kjc1tGMrBDdn6
SIaLG3tKQkm3rS8H5NonUN3MNeiP4nwy4HItmuogW7IYnri4cduRUnJywjhs/K7cSWlUuOMJKlOu
fPiXMhQADuXrVMA7+42PvUsCI2caeoOFct6wPFwa7myxbFnuRipPdcixdY9xzo30hr498hWfyiq4
u0nWo50QbS0E8gCSa4BT9gZkI4smPrY+hyb7LuSc3tePwIlh9AbmnkT7L6ANRHyd4WuAYpq4KqCM
vQGH2mEqSNkjx+rE8PYNKEdOLZphX9u4vXE2APjzrIi+zzgVTVy84Zql+MsanzlxvDg3se0sOOPJ
LQI2yatK0ly/9mM9YoTtrSivU0/BN/TSPQLkWgyCFml3UzE8WlkR09dUVe2B6+rQm/y67p6n3yaK
z4ih2nslBNwF4pxbYdU+MHv0StL0457rmANVvQ+8sY0lbXB0MOswfVS1r6l3ZauJspVt0ffalsgP
tJ0w6OEpm7gC5lsQDpPxOEXH+vbkOaBUm6iMofaLFffQ5YNvQvENtNiwZf8hnOkMqhYPOdjCpyhC
C/lyq3VF4gX/Bf9pYamBiZ/hiQMcHAz3ph2UgTbxezrq0vsCnsRGkei8aq2k5JYQWerrUuouim7s
Ki8GakwwdPdBUvU27Nelqiq++7lJrVPmZde60PSP14/GqtkB44iISnsRpruqteOT0iYcbGq7L5hV
6fMHY/Z5DlRH1ygGnmK2/VACAKIBSWgUOrMtsy1bT1tThkydg5bCWUg1o3HTFpXu5U16g7TRipWq
IUm9bSEZEwld+MkwwCvWB/HofcnTkxA1ztMLq38FV7VMkKp1GEYO1zG8zUp9uBIgDLkd083j28FA
hlTSJSU4tYSP99eK+m8OqWnJ+8NJgo+wnwdUrnHNyzdp/bX8OD9AfPMEIyqs8VUQ8hlHhf80GB5Z
h7+W/2NYcGr0Gu+lpwqDtrQU/LrOQ4ppvjUc9nYBsQqlrjxqgEpj8KOhliqmJ/anMDat+TkpxPbL
qYlHZ6KZP7vc1JsEds3ejPH/4w3Y5UN0DwhWhmCLL5vhBfAQdfK61ziqz6I9cjhoM7aShOu0hEOG
p4yNOkTOdp6VCLBR+1E18XOrBJUhjsNZCn92Acuvf5B4cMFQoZkIx9T7yo0ofNIN3AeXHGr9tNlj
PG3T+pVR4MQX+qDFWXqWGX8iXctigEqjASfuy1iqBWUX9vXWCtibm+Y3BkpFXq3v5/TNLO34nz0+
NtH9quKEgEEc4Ug19naPDacuecoAXQp0Om9FJ/XO87fW6B3spt2BOfM52jtWatSXhY0hAhJQWEcs
ooHuLL1JT9fhQMU1qS4yzNwq0A5H1Rh3PVKguiNSeSrZG7o7iDaKt4T2gbwWO1hjExZhoi3+6zCz
oZlIY+wsNHZYF59YvVmhOzGxNCdFT5Lt+Zfm8ayDfx4OEuMny3pMhtv/Fl0lMWvbT7BF2ooi1gQZ
yOo21ypcR7wTJ1KGJRWA/quVMn0zw17+QSqfYJrHpKwCSw/wFwnLdiNenL3WYChgQLy1a3WxlraF
rzGrlA497aKpiwqoc0boO76awhONrY/4bB/f6/nM+7JycqqX3OXK9LlYOpqlklFo32QpsPpSqZly
S7s3BgnUhxP7ib+gHSp6iyPFnwpvJuh8hItaQxZsn46GxvRWx43Y4NcNqv6Ds+DfPymII8sbY4TN
rxNCuR3GEyBZ+WFbGbJlJwCiDi+JE/TtzCiZh6P88Xmm7/On6svIoMY9xcuPrToxuGE/AdP5RuLX
HvaSiSMTAYqF+vPvyWqduVju5u1d3RZwsjqZqZRFskWaStnBQxY6w1WcWiW0Ud22kB2A3DR3Nb4i
qsbfxxMQtkj04JyyaIeNbRVPU09kkjn/Q2BL/67KyDFzYk5/DMiNlPk1i1yf7yVyUBQAQc+InGgW
AH7sRL/cy/GXqzYFciQI2Lsb8S4bBVdqTgZ1DRz/myYR+ABjIRqEyh38ovraU1fIgXO/Db95BGgA
Emk4vT5t0s+rik1qrVjmXo+dues9BV9gzFH5RpDBQERH0DnbPnCe7NWrb6WGhmerc6fBYQdK7fmT
9y8nYjF2e4aNNYTb6qdqgz0llawAy8dzpi2UAylQJNv5EeSU8fMWD9rnGQeVhc4FN6zY7WrNcVjq
azIPfiD4S2+YSWzo71IzVRrWXmTw6E5HYa6RES+ifqmOW5lJNyjmgMYjbQCTh7gmbPs6wWdrbDBY
th9SuvzS5a7YWw67OY/VC55qNE7u925CO706Ej0KOen7e7X4xGwSB5HH1acJxPKxPWqxxDpLx6TN
VKopFLUKWtIuYX/zNrbwmAAjIVFiFK4qklr9y4zxKiitxZqpgTKAgjyq/pi7T35ibQhU7td4btJ8
ba4r7AW1mbdU0cwLvE1WRgoP56QnAfIy42D9QcCeA9jFsjfOVRiFeRy5f6z2RVzXtp0df7huMj+g
dSnnH8RPJvQ6Kwkq6I9MhLLdYoZ6XohP+KjdhiuBOmklJbdVl/uRjZvIJHeCQzmpobxfrY/L6qod
js7RxwKxaRe8ES+3ubHDlCwF5C1I39lDgwe0OEjm78+egb2W4C5nYzPWIv84hsGejQ24rPckBRbm
Ok8wCEqRY82eoGVZgRQ5xmuCvf5mtuJMszJow9bW1eQa2MXLI/5J+8feKkU2PCZ5q/c7xBZ45u9o
nH+Swy91PTua5pgHcf5FoYUqL/5kSSGIsAPIQzWiausVG8NlX2Sz12y1OK06eKvxij7L3UdCqKCy
Rl/+gF/WPtrxqi+J4DH2/9DY5Hn0Yp5eYiq0asm4K4bIDghlwNjqHyrIa7SkK5lFQoeFJO6EjVFy
iuxn9blPVnqec3papjBNg7Qktx5zwiRMaQoIDtbA7/vSFc3uNbmiAgItsnvliThEz9TK6gKapT+2
SOvkinC1kOGQYwP2kPIQIae1Ink0Okr+u4DpjnhOcxjN+TG5dNpY0aq8+55APoTCaNJtKLaWs6a3
59By1v3Bdde/jH+zZlfBH7PlXd/vxVYKEdhDgqKllyfIk+cOSwAxddjnxz+yY2zl4Qf+LzEZP6XU
CC9gdsO4tnY1hw1alKyF/oAw356mQ1ou6dVNshGkQrNH4vV1bkPnKJXyeowKKFaHCG3l8lQq7pEx
ENvJeYZd0wdisLvMfnDs8LZlw1e8bmrTePAU1caBf3whWmEeBtTCKhrDquFbn9uEcMPQgkzU8WL3
DhR5cqUQdCmaWGSQV+3zYvS+2y3WsIgUOHJcnslXmCCeN1Zel1mYoYLhmlxM3KaQcfgkE4Xa7eMx
XlYPlgbCQfdOZTiFJxzwCgDcDHFGQEDR9wkHJ8hCczmUn6MGCdfrXPWFx/fEbE99e5Q4kMUiKqsj
Ozt/5bgBy8+ggL/wiWw0FuSJNSo8Vs7YUGuIlbghJCULcF2S/q5i6wgL18Mf7pYa7dzN1z4t4va/
VcQwPW5mCivE5xc+JihHtyronoX59FhmQhUL8BH3MaCH2Y1egmDHEOMTpcpO0FELpRyYTd95DMA0
t+VYDhzhxV52P6qC9KySFQok4lCdhh8bV8vr5LUEiTh/bJsfYhHb1yqWapPF9Gl9zHAJ/6OMx0W7
4NTNRoKEoXDwg33Vgd0tHqxliMTcputh0OKdcyVRr0haEdravCBHIvGTbjnNgYAcDxXYRxQfXztT
uzb6DJZSXxAClQ1pJ2s56vStp1bMuKFWF7TihMXD9RLFQ8oxNYGSj86gocRgDNppcdpxJwkf0nXv
rQajiHHQ0tS3pBufEouOfCmfYx56gCF8c0vKJKHL1SPG1dC5/LmlS39jZKVX7tGvgUwbu/x+MPKe
zfHjSYCEGfdInArJdUECQ2QyQprrea+XRkL9ehQc+pxmTtbiZH/ktzj2cj1M1Om8kxVF8DpAzrNM
zRxw/Zx/WPWYqPBXJOETC8/qnJCv7RMynXYHmFHOrg68wx4QMzt0u+ifn7BdRFrjcQS6Q+44aZ2v
7WP8k+4VZMRVccfo71ipqP5SfkYHXhX7z+rlRFsAwFtIq7mHrxhb1ka3INCg/GKd4SMufuRwqnoi
pJzJVPuDOP+vLlRUHIbnxZAcUN8pVsOR/ZjHfbLhKIQ44iQaO/2CMhcQjrWkXWS8V6DAES8qzu0e
gCdsLBFU1Zzb4fW93IYSEXNFFSf6kvGtT+tKz8EsTACu2gEYQxcH25kBsjr65ErvEbOYzIogJnx6
H8I2MPn6yO7Yja8s1cwljTMo6RNq47LPRQqUnPFcgWU1QChdI6RDYwbltA4c+KAU+pxMKtc4+THd
XxiBhZjWkGduS4lc6VxSpVDZw20GEo25SkK6CUE1lhvBX53KEUlHEW/9w+9Zw1H3/c/GMRAehv3r
6CiQfvPVn29YvlvC4yIaYV0VVsDKp1LdWNitqgl/wIHslhg9Qd9km0kw0DP9eRK0RtMHKmGuY92b
H47JJcYaW0Bn4qtIbxxDfovxJQJUL1gVk5bggdePw0xPe7tnlcvLfAy0+XxNpSCreEPrazJoBBx/
NsajbPJt9vj3KvFiFvOSqrH+p9K8yn+/VyNWfYTNdL266Y41TJBEYO1rwSMmKM6Tmn72pMBGvQGZ
ZNQ7SDMnDvEg2N1XYWxfMwaQg8RGJWH7EForW2K5jIY+YEqCPXkWFKawXHyOeR2/ZnhHz+Mbf4R0
NmpvIURgP4lOfHiWiJ/p/SLmjTOQgLufW4EB2FJLCz9lXQDIGkl9R99VDGHJdNbk50K4XXhev4g8
EqETIcjW8sq+YoHmLbUDylR6pBdixrwEnFfY05LalUjs5A3h/xkEcU1oK0Cm2Jaxg7xQ3pwRTRXR
BYRa/FqNJM0Vg1wKXuWZjVjksII5Zgsys8ODqH7b66E2z4qB9bZn2oAxHMXTIu85pGpB/cbVMsfU
3yzLOub/x5c2vSG8hQSYKlT1JiTqX7X3/BC+V8zG1KbfDXv1doHpxrM/0AXr7WcNRP5RVsGN4CMJ
W8t8p5iA4eFnPyM98kyEEDNgft+TVf7NNfDUHz0s9HaFmYYMWmmT+K2TS2aVf6MZLuBriDAjSF1N
E2t63cddJFteCodDUKetPdvEQeHB2mW282taNsN4GHweqqP7jMKft1dVLWEZc+cBPxDspvz/IWjT
AL3t6HIA4LZCr2ZXA5KlRBxB8BvuYKAiC6j3JaRYxjKUY1R0KY6nd+ayHPhnPqDMEY6+EahBhkc2
WKbbcoj3Y7+eK8MFeuQfNzvSieSY6jk5syQ4h+vSOQJC/4Djop034owGwuo+xjF8jDoNG+P13Bto
L8m0pdCf8Yyc1WVq/nPZYv9KFwP8vC2bVDpxwH7zFVpcP4qgzdeyJtmE0FMtb94cQXt1pQwMlXcf
INIowV4tYheQRBr+2oluf7vAMMO6OGlMFKjw5uz0QGYXrzvpeOb5LMFvpS7HHSwYZkStdyva67wz
aPWveYNlSU5HQL5VwIYBdOf0kJ3td7KccsU+mBkWqcT3ecc5IHRxGXdrYHGQ8FZ8E9IgRTOvvIJP
UQi/UYb3vKT3jXM29rZsahOq1bucMVJqYxXrMICVlL9183HQR5nDgOSENoqjU0jpWBrqWaw1Tl0n
eoXzQuXU4l9EQ82bG+mJJ4Kue4iZdpVqAEaxXGvTprR6XtAPapwzMSub8RJSnqwh20SgsPnKHfK+
tW0b7SBwj1vHfM3qQSE6Ba0N/1WCxF7XeONwLlAb+uO8cB02OeoDL/PI5TtxzpHdAKqge8Og1HGI
Hmkt/aNrBAYXI638LxTd57VrQ2e06fHB6Lt5gi+XGq4HjQH9O1u1v7ZI634pFQBIxvfhQSiyZPRy
nj4f4TD5DeC4SNggWld/xCsG/4IiKDUK91iW1RKmqTB4BZQCV4SkkLWRUsDeDEpxFCVcSfb6NaBw
47+zDQ4hKwGBBG0mzXjbr+JRkO4L17YdvBqmnGTFv3pbcFUGVnqIqH9qJMY5WP6SYqRZRLPsHQYg
AulTRncmMBSo2pEXQnj5jpV/TCIFY4mNOO53+Rcb6/pSq8Xir3Zm478nNfOmORVwpY6GX9BP7GA+
HSbsZdNe2X1XFeyVYuBQo0G4yuutIiYUSVM84D2Le/UN+av5eymThuuRhyrqBxK5i23TPG6cFji5
SG9oM0t0wofZDR+Auj9pK5VOJJEGvksqXwEmxaFYceMkyHXfWo+Z6DvaLnUavmGIOzweKtJIWOz+
4ABxGDajnlsOTxRGBMNr05EUQj7uyvAlmQn1Sc2oABrVUS/BfM303feaEEMdWbbU5lZBdwL//6+R
UAH5EJldHmmXPgmN+B6r6+f+cx7+PzkHXyI2M4ekykxkrPH0u43ortldHtNCx25f8KOiN1SvJ9Gm
OjrOe55j/7ntWwo0gQIu+FXoFbq7PDj2OvY/miQ2Jb+AU6Lg58e34k+jWEXtO/3Bqni+Z5Swlr+Y
qttVE4BmLmzqgGI7xEwab4f6TiN4jgZm7TMvvYedN7Fjn/R9fPwSU/SJODmw2W1//NB+k26Rnq89
w8ErIi1QJAmDxdo0P/DNTC8hilV0rOpq4wO4qXfh6jGzC7XEjjHH5I0aRm7pugXh0JJRZlgWTigG
5F+no4kB4MUi91Vbw3UALKYmMUkG9l/TJu77Wkna2DxlS0P4sFK2bkRyjZd51lgdb5eJq2jvpKol
PDpAEqEQ+EHVkTu6jD1PfZoz7ai9T3QiLCgSbUnFxcmGVNq7c1fNApJRM+MnYoJNK4brBGy+hL8t
59DVBNElnWEin267ObGaL0YNoo0uNIaLEuSvXjaBuH7gGfIM9bjHsFHcfmU8bIFSBdP9vM9M4lnx
lw/+VxrscWn5vdopDK1Bvp4Vkn/TQThOcuLaBoCvNzaJ8qaj5wTgiAPj/FF4swUqqtaRpNR4ryXL
WF0eh8Jd1JWMyOKG9okjWg/5QgSK4FDLwqdxpfQRyfIyNppYZxfqyS85Krk10nbO3WNeSCpPsGE5
xkQorh6EQXm+gWpGZ8k2KqT6yRUN7zwkPoGzjIFW7SLMgs+eJBcFazF56WIMvCc9aiKQOJ7dKRqD
y+lOLvtJ49g+VNtfPK3rNWbiFuihJruiefFmwMqgHtXl9xXrYJPc7fdsjdSPvZGLcAuNl8ZkE3E0
fV//ndzKhV9AHxoNbZHP8iktV1QYpbiHqCfj/EyU29/3NJaFxhknQHMSTwZdoXcxg0twHGBsn3wi
nW+8qeDI1esbFJsrR6r8hERIzunI11oz7siuLiBKNX/jUGSgTGmUJhAraId0yAvMCr2hHMBWpyk5
47E269vXEE9/ldI6ATROFfQpyV765mNz4jH9jErkCubT6G7NVzMYqvrSZxLIE7Qz2vXTi2msHl7r
/wN05T4Rwrkze40Os5oEQHCO3QqDy2GJL3bY80/wPneQwiOScaHJ7lkWEBJ2yBqlFeSSJcSEMp97
hG5fFKZONzCAtbsFQ4a0H1hiM0uwYMMv8zApWQsLcS/iRg57Vw+WWcnl/s9Vb4PMC2m2WqJinjv0
2e3fUOjK4DsmxqIHkVud0cuexDU5N5smi7zlYyBn9H+qeIBbGdrwXnmlrRM+49/OCccgKAldyFTO
3pC2PYmeMgmmP0U6tRLOrCUEKXD7xf8wxy1PHbtKEwQ6jAXEIJddrKIlmZsMX1VO1DBuPI8kGiIS
w5uODSLFf67SZGrwPqRNFPwYaBypB2AwxUH+7F6UxAEJaUEty073+pvDt7tPjWCPJMFcxYX/5Cqi
oleeoeIB26fpqTHhL67er76AgPvJy+LSvZvSy79IC/V0vyBtsbwcCucu0iEzf8K40ac1AkJom+Tc
7P65yVcS5emSIIJ2XzBvFqlFmlfhiGf0RVBJGs0yl+x4PpoJX+5jLHDOs1HLXgwtFFH/BpvI6lgL
UY6J0aygMJjDNWUD1tvJpEzfPXcQwBuew0b21b3HCedTc5qzameS+aTztvJuiKghODtsApyg2z4Q
J/DdVxpoDmH7/MERv+E5nUhcI+VnXNYUZDX2dmFQd76e4dVh+CFoTMioUVCyq8b++CGOzdDN1STZ
UncR6BJSJuV3dunwvbw1ZUzIc9r/vUFkVvuXftz312o3ou1r8t0kuDQU18xPre+c7DYCnUWxmsW+
tJPzEa2ohb9QOqb0JZfc3y+UAWqf72lkUY8KSlRulnc7mYSBBPTauDdVYcGFgIOmbPEvtK7Jcsid
RZ9NwSXKpGBx4uC+Bi8jbjWnUu4Ot14AtwbHuQAbhlC6T/3RWOxLkbhT+41AnDJGYVl0R9cvYc2d
gg/3c3A0dpOmwXsaBiNTTZgwx4w6HFmf8vqbltO2evH6WaumUJuWuvBCUTyDI59Z+aRroZlykhiV
/Po29bqo238o9otdWysqJXqVYxf5HHgD3KPs0Nf533TqwGNboqwoGl355ga+gyZmhJIrURfDerau
7uvAbrYisYCg6Xpa9ZJVXS9XVEEHxmmIVDKNeQy6aK9KvS92ieehDd00KAwfVG2m81w7kFTzlJlR
s69LJVKIsgF9tN4ckc1Y1RjWbQ1v5YEbdDY6ax3DjiljDFelwCbuJLyGo6wIU+vD6jVGjJKWtTog
miw6xKTfgZdVwJh36O4xSciM+c08bhc3pDYcdXC0H5nQCJqnLvuUzazs5Q/B04Y3f8ZwIsywyjWp
epv/JoBlwcv2Aq2izwIO4W0SNabH3x6u1A8JVh+UgYLwYtb8Hws4ZuOaO4keJrvNa4V9W+pMZZ0+
4bejzAcHYi560iSyuFJ54Pi2oMxrt6Wp6y2Zx7QywJfvHOZgAItkjTpGK0A7zLldIdIyeampjkDh
HgjpvOOnvkt3ZUjnQnDTsQBpzDE4fQo4JkhLdSj8fy3fEmtQWP5Bsdbi3kbM6wfjT/UCAKr3Zg0D
h+TXf8TQLK+u+pb/mqtNdUeatm/tuv8x97hbpyuQBCZj3piFsGo2qFVLajxTxiD/BIGZAekT/Gi7
8Y+pGgndnBBFhyLW3J9tu6kbOphfVvegeQfv1HnIVWFtb3ipU22COG4+DqBKz9maHJ1FI40JMa1i
6ikJu9CD1LVGvFEwyWnRbe/VWHhALtbSP0UdyCEqq1N+eO0dKFV+J9rpGWa/JuA07RNlKTjyHgq+
zUq1jZtRC8LrL+EYrD2QsKKC40ohkzhs2A8QRDEKGf/BsHkPO6C4YuGvOqP6xIuN16q+LCLSx0GJ
YF2+BJOr6O2ny5uTrgMOUZARzdEJHv+LhoDAsz+t5Q0CIcfo4xKMYUB7XmqGYRISFWVm9QuYoRGc
1B9PtdfmalfBncfm/EPQ94pnGvWnKP8Foh9/LW2bzbLTUpUxAerXo/8ThyM81rdn5/037F/UsuKi
+0zK6ZYqnxBq/fIlRyczoOMIVGWlHry+lLeipCMWQx2516X7HQqLAgt/ynw1nVTFd8BjdTwxuI5l
IQ/opgvv/+H6FXBL+MHzXkU5FVznoyYvtN5+6+MBLfhV2Dl8no3IBRjYC7yinyA9abSGv7RERl9N
pl4DMkaZq30voQ2Ije0E9IPY4yM/1936sqmcdeCGmWc9kc1HZY+HFhvFLIVgEj2vwD+gDnH1at/+
VXyQHL1v2f5yosFKvi4O4TZTR5+4mu/TSnRUp7/GChhxK4vdIMeKamv4qvTHKkK54e/7h6fgmnuG
pfCtWxFtmHl+lk7660q/rnMddcVE97kXloi8geSnvs86ZqhTK4/oI5Yijr1od21JJt7ktlaYX5De
/CfMmRdh2FWHeYX8WdD4sz30P9URLKZ24CBSMmDZpG5QInOZOI7/YFbyLPIJFr4sDwQzSunSBmqh
q9hMqKzy4w7VI5FgErbxfjI18gyM3gSA4xWh9h/+leeqba45Z4FlsywBzYFslrhqvrWk0BgNFRrD
PEA+RLI1NL444qpBUjBFwHTbZAwihnIjj/VOh8tkSWKVQv5dmLuKHeD5zkPZZNR0Z+i6PU54j5pN
csNUVQvw6PuQbI1tLViKEl95RV6QdWm0b04m92f6gseFZ6wPPXNcB25Tt+so6C/YoTIzbiIO062I
xSy2jUTGsjQMIrGGnbZQ57fBRnVi8+mGUECf4WabEv9jBQCJdeAHuIlD0FX9bYG1t2omojOJAtjV
9Jevu9Ldu98tRnjMOkW0XL5tK7Mu6uUkjc14ylQ9MxR9F658q8xjp3WaH9FeDIp2Bx+QgBtjFy6Y
j9YDBl1XkFgxrz0u4lQY1SWBo68aV7bFFX3yLe4iq3mqTIgZjwLsCTqwatcpU8v+APD8GzEDERMv
inFMYnS60ezyTPJ+tH4O26l0Nw7w+dO9xIEoTWXMz4kzaa0dnOCBpRI//2eoXx5ZsZJgjbubXfWP
oCmFxYJIeWiCaSt6mSvGcJi2fsSOWsyExMolMLpv5jklOaklMrypjpQ+3EaL4Z31OcTvoHLM5Pj1
rV/S46hrnxCa4uNFrcvWo0Dk10nUTPdjMf+o/Hoy2h1VmCqEuUIEd14lrK+aXdBJh39zxhIxrt6T
o8p4QEXLXERV6CxLLt+7SOKse4o3LnZL90pgU3OfSKjyRjGibd397cK0TSEPMCKfSy/8ro0ltvvc
zrmlawMq/8ouqaKKOP4HLWeBZMbEjkGJVsK6Zrg8/a4Hlfx6thPOQ0SpGA4L39rUKQhO6K5luZOa
KU/4Aw7yW8myhhv/piVScCpxAsWuqZvPzc1Cr+pVth5K+uX352+kE+pvkY+1uPc0m1u/mZsTISBx
eP3HqsNTcfTkha4UTAfdLrJca2t1DzhuIzokLroF5toMTlO+VTyxmtX/4K4MRhYLyysAADJs1GR9
bLKsUZI0J13nIXbL/nIPHAo2Cno/cXiYcaaCI4Hes0w/M9QgDG5IxP/K7HpPBysOd0qZnwt9YmZq
vynx3ViHEvpKR2/Z0RLeRPBP4qOVYMXnxYTgk9uuW/yY/aBfaSmlKpnHTeilQop7FgUc4wOxtjp1
WwPM28yFeUxFaziql1kLp+lcALw88ogZ/EvW7Lrq14NPzu0KnCfADb8m8XYuruasYLfcQ9bFNqTx
wOX/w02hHi8E6ZDEtRaVmtmOOuEt0DVt+AbRGRkihE1bDn3NJC4XKK0iaDSSvk9Q7vE+WcVhPMx8
bsnfHtK/rHHLZvQNndXbHbUFzBwSSbf8EwNYwPTV5PY7lIaU4gY7TvN3P05wHpz5Bwk4uWtcrxxT
bbQaYHBGVapy3a3nAadHuLkzkINmNTnkiH6N/wxjUlCruvSOcivMYaUAaYw4JO/d8YiD+0naT23L
8ar5MnH2Y6uvqvHN2xP5P96P+NdVpSNupq5txcqedhso9rJurTL5sF1fFzyx7MzlQPnWpHN8/65Q
eB5Xd03/q32HeVejplSaxAFkEjzZy9mtR7l+0Fy+o0zIeTZgmR5mA3UdqsHUCr30obEemIHgKlXz
8SRrCIjSG6sGkrT8IBH8luS67KovP5MkBRO7Q3rMxXHhklqcE3pzLY7x4FJm1uTj2IM5VvSBrRID
pWe+fAd/HGSNkcbv040OblrYhzlS8oCwLETK89nyazmN0NY6QKxOYXrx3a0hvNkr+pj9n+M8zckv
n2rp5MAeGMurjkaUaMLhTWpPsUWfgEYexii1Z0byrVCe855j0LlqJMIP+qR3AL3HaDT8lwgh4nhi
3kPYs3ws33HvRf62IxHDgfM+OGxqc7+yC5ZV0eS8EObLdwsfIieZgDYFT3o464RQN3Q9pDp3JVhV
Su3oOInNxzbwvMVgYZyqgN3/eifL/5w8drQdFyy7bbUOBiP+Mc5uSOBcvezLo/JZPCo8Xpmyq3S0
25TNGtk6YjUfXcdxTE9EfNBpmDfpKa/oMtNQi7NQns69oLf01VhdrXVa6aSkkFAy453DZ8ZfFMZA
timZWYLwCjR/1aH2GNSgaLCuzMXk+wkvjIZ2cVC37qEHEpqyMk/Uri9EbZbEm7S340KrP9R47M/l
OC+S2BlFY4+DEStx70hkNmBbfnouxX06SSD23hYKXbN0theW2+0TyDD5bhy12VSNIdeqJdBuJGdf
NSg/QYJSchH4syyaNvH2crKHpVW7nYPs+YUTvwrg9oJj+nYnIWFYWGw0PIaEL1KYJicp9dd9OLmW
LJTnIaTKBmkln9HJwv1lwnXOEtito9mcMDS5zMTpxUR+2CNlzjTzhGPA15OJKMwyfnuzXutJA+nH
IzxnT/8oqEbW0rCCYxlzLeHXt03Oa6PRBtkBxc9agZ47yk5Zjun+jdmSAXQH1Rxz/SS5ijwh0pqK
62MIqtCUswcl5X+PuGyi4DgVYctKLij25Nq5+Ourr2RLDwS2g/jxWUAd/z0DZeNRcaPVK+c0Uxc7
W5eYXZk0gMtU5UNOGQtg8ySeOCsqfoKCdGcX6hIgdnAaPe9LFs8oXs1AQ7MxZwbU63AY3m20KTNb
GzLSOrnBvcOuwpoP6tRVDB0cQ20RXfXRDsjT2n/kZkN6esZ+d42zZkcQ9YU8l98xaUn9fhPALsEc
YZUzh7JJOQzHyqLrXPVh9HvNabs6Ok8/3d1s1xb/BLJD9lZOyTofurP4CsczIkQtnef05wS4jhzR
tSF4bybVRAgFOlqLHFaRZ9/Rl9k7vg4WvNrhlx3qe5V90lk3VQjg5czwEIzm1/M5fzebv3Hnrv5w
rHkn52wF33D+R9dKARt2K6FWVtC7DfI9TPhSc6/yN+eeA8mK8aidzwJ5j0JMobmHkEvEWiuSPfdl
pDOdcMhIfdoEiPa9o4ZDwUYZeCSV1FwBX/lwdp8OxxR2EtB6kehYZy1vOZVPKLlISdkIqMsoiWvX
D06ZPxhLpuynlXIbTG50C3BiCKLm3WDKo+ZNA72QtsIPW+VTZfd73VCFwknxkxSTaslHsX3n9LCv
XYavJ2+VZ3A8jO3mvCSPcXgzruq/G+4v+BBQEd77nYSt6Oe0+RNSPquc5C25uByqU0oOO0HsrsXz
9vkv9zf4i+D0KTcBxBMGAmjds1FpbbrEHwSEWky67dfAMxK0MjQUzGkBSxunTJk6gt09N3aMPd4d
4+YhDPZDhRhzp2ZkSC0JEXDsWx7VZbjrSWYGSP8gJVWcl7eDhUGKsK5BYffy5EoPfpHbQwrNtjfe
vLfllsIJ9COtpLppM5svVblv02kbxTh6uyTYkUkNNIC8OLIjiWSujU6rh6swnrIrLM9EojVhPkHx
hI781/zJXRbLnQFErTzWV/47+t5jZMuUFzL0lIaRqolcVAjMlZPZ6PLCAFhs2QDG94u84PWonM9k
dVNvK75s1Wtzg/Ex5iYtK9WyN/v5bP4qVGgNTmVP0RL2P5orsSry9UUeE1K9tTXVdvaS2U9PWKt8
ehO1safVcSau0OToXFMDkJhT5NHy38597l2aJCfQhitmud+bM8CMD4Ex8KmvPmFQRrT/dyHqLQt/
+cHcfd3913vo4Z4wxpNrHrtE1wIMhDPAJBBinpdtUoCHIcj468m4RdqtzJsjoEtUZQHZQrSdHco+
5vQD6HFS3ENw/8ik4DmsbZcImKyEYDeecodby/UeL9gwID6++6q2qHBkgStvydcMybiMiRoY1xVk
r3CBmi9agEUxPPSaC9BC8pm3UwfhlP4TZ0Wtw0Y14Ia2gnBwcqYcehmRAF0yrC+bVJf/9LFmgtwP
8+NOKN8qy7Tcr4p12f8WCFBxLizkvNru0vxL5TsTnnI2S19ysVpQA7SsaPb7bJ2/dTXt7i19g+Sj
MTAD9rIGEyxJ3XWh3DfJ8LeJXauIBoenljRXVeJg4Vmmt9hCs4aJyzdPZk9x8DqBXji/iSPUpgYh
pDYjoMLi8GaT9WkbSFCV6EuZJEz8eritTRCWhdPimn+o+SykX47IKGZ4vMT/anSlRBjAaHEpzgGF
ccOvJKf98oyuIDnv7g1BmT05lJYp8JBhMSPPBVN760Rf5u+d7jdgA0PLAsUrYuTpAtEbrQZpTpe/
6sYnC4NlH63YzLFT4gFmW0IEBuIaeuy//OkVDWsjwq6jo9VmtNCoTCkw+9sl68jv7EzHk4SngVa0
tv20j0rvYn6wIjYi/QxA9NCWGZi5O1Q+yfqZvm1R8E697LThfMDK9mCfLbAG+eIDlL1hb/h2YZeM
qMKwHnj4a6Ykvi7iLyxMUnrBnyP/V8Fg6+FgCG6MSBa2GyfcniJHxBlM9490GY3L6sWIuTgJlO8C
eZJrPMNKoIL8WVoQyDk1X+ZwZeVV15T4mgkZ+j8zTZrgzRxGxU3dpAiFBodKgKdxHQSrxNPWmbZK
I+/AJbnntvnWF5G3Q/JTaZpoaARuMpNo8jSwUYoVHf2VQMKeadH9e/HVj2jLkxOQvJz12b1hNIaM
UCp/PZ1DI1NK/iqG5X8yaQe0tovjWGFCKCARKFqPglJIQ7W05g7eCEe7DlHyjWEMBFTywEzPZaSm
/clnqjD9NgOtOvr20cEw9zlTt1Hvyr/qV8LdRLtsU/wm7oNz9K5IcpwBDCPCqlt1J+y72TykVI3w
SN6cfdKQDrdFMQhUgvUydzC2RFCCkY0tc8DapYEdt4UpLzxMoMBeUuMNO/5UfbdaFrBuZRZsHCig
vYgJX/AIsJY5ShhUJEa3L3bVD95UczZrY1WnPsgKOOZJNTDIkLg8fLk7VYII4J0kfQPsrFNs64Cw
xgQILTf60GCEyLAGNgtuYD2o+ByuuYnclw+udQGJeAb79fgPhVlYb7rvJDZd773GYcFNAOz/gZ7o
n0VHi99gUrJ7M5bAZhWC1e2aPYqTRjFWiIa9+hgJEbX4V8omdzwlEypsBqn8R6nA6A0plRjn6Pvt
+f6+CoQ0yH1Q8BcOxThC5aCZYJIGIo5SmHnEYDKOMLb4/O4WCTgQa8KSV++CpnLLkZUMWfFZDvlL
DBbXtjLxPZmoBLKNlaTrdWaCVcONJoJYz2wAGumBq2iDuY7/VpmQv5w3Vc9nZ/zeNCT+Ckf31ejt
cUAf/4ui/awMS4q/H4+9bxmYSOhoYpS8kTmzlECy2FpSBsFV4ykoafJkVa2GBTy+ot9p2kElY3pS
yl33YXaJ6DHYdp4NmwgCCNevbpKynbdJOa/vzkbXQuQPCkDJgMOG/2JhE/E6XEbpezB9x87hyc3F
NQDpbrW41p/aHiqEIk2UR380dOKK7k+QG5fwUlW8VzDucXonOptSXbQ5CWTb12VcnEpQZMIGXr6I
teDiJenLJHtZHvhNBx9Pz8yuXf7SPvp7vPnJRNBaWCvHPuoI9B2Qu6Fj6AJ0FlqyawsVNR8LkfdS
ulZqi8FhdF7Hu8tdmTu6ESmo/nw9dSTfNH5sJOy7wyEYuiCesKF/rMYTWoAXhon6OTKLRo6cFE8u
ZcOwu/6yS4MyD5CygfwrsPJY2k5aoS41nr5jxFIB4r5XsMpEo93Nq8ahVjVdliqMnx+wDWE+062X
5EEupmHVGjAJaZaJ5aJrKGjVlAvkGJ0rr1E7UfdyToX+jXxaproEXHFtKnivLuvQK0VXwTwu3rMl
g26+cCv8zU7SUHoA2CzDhSZqXtMM4SCsAmKDtdgbCvphIudXFT9KAnYsn/0eJXmoLArdtS1M7DJq
SZVIUkOcqurUc6EzwfSI5HqveiJrToyVIKPlXHGTk4tFlPd5qE218JuaQn+KeKot/0dOHUDaS0W/
M1mRPisjd8qsvXMrm8YMjKoUcMSEuO3BwvkD6MQCWh+zaTUR3j4l4yRc8nkJGRw9YdSiA1Nxfqr/
gJhyPfmabNSi5iBiBqeCwVGOlk2YNK4pTYUzZru3s+GVSL8B9zufQ5WnFyyz72s1DkfLoj35u/XN
JUGNjFOXfXOzdwcX5IuX6mM2y2jYz0D4RNmGp0/0REfqmiWi39gzKO0bGj/LVkHxtcCQ1GpGFih4
KH24lA9gYG+27qQDMo/Z61HChsBSh6VBiZw08DXtuY/6+3Bjam2wWSQz8hyA/D0Pq4VaguwfR6JC
qa6wijjixF0WNwitwwgfjH7ZedT9TV59ZH/uWZXeq2GYW8oniS8Rnedm3+qZRO9sRtXU/QNG5xpR
ttOFxNhX+aU3hHnPlnfb71F5+h8R0KfkNUXsTdDqboaExvPkidk85qHFQ8hawMHZ+MRTcfposPBy
/d5RYQIsm/2fGqU8znvGpf+5d8yMpwVb1PPxE6IVc3LCxQvgJLnfyrAoHCKh4r7iKzrlrPFc6kuA
BqQJB6y8GC2fZMxc7onmnP+VQ6kQmUb1mqTzxRdYFgf7Dv1lhPE5YDIh4+7+ScNKXFbZZVDYXL1l
YHunmi8adynot+TElRrBylcYFGQKO93skWh7TewQtpUYX70+jdtkBcCoDvounJplK6f4EtZUQ/08
IbiIE8QujS8PrJeUb/XI0vGgXyVzfWibFqcAO2+keeHdu3yLKBlmEnKTdzbY87BreTgeXKiB7n/9
i7R/toCbdiAay4hE/8Jy0s86VFe1meZpqwdtVhOHmkHZXdZIKUoFO25CIckh5c+59RMe0aW7FZDE
yrhPa4QUEi6Q9LXgr9WNdMYYbojiIv67IEIyOA8539JhiYHPx530i6twZxhVS1z9P4FmyEPE5OwP
2MGfacPzH1BngWYksm/TIZNoLjBAKbwaHQKOXjOHDE3Uo8eCSqWc83oVHCm8VjJm4Q3ZzykbvowZ
pq02hDp7AeKoTSXP4A/oYkFzd9WzlNi+Tpb3Zv2A82VBAOEermvdrheUaq54HgH1tQ8UIf2z8pry
3u17zbPgFT0sKEGKeFqp8Tjsz5QizL/TaYGC00ZpER4Espk0HGvefFau5kEHp4Jx1ynhXmYiRNI7
DhyccisofpmY9wT2kvB5i6l08CBVv8JULXB8o/0yjfIZhrEM80JZT0TeQGOllT3tOQaHtNjQjMk4
EmQHSJBoG8nL4JB0wsrdrKmcaMecHa6f9GSxeeLHmyz5x4cmEQzZ1Y4J8Rcgoaj4eEb+7KApVR/j
wgaJCO+YELqC8I5u1oMU82C1vaQaEauvyadTGrMRBv+CSyealu7brnCe5H3WZfiYFsKgfnsuPrna
wcibzInA5RpDAxz8hRFhiZW/HWTRrwFDRMW5QNhPz52C7cO3ondrxu+mxox9UEyjmi1w0OdjpkEP
fp518KwtY2b8FbCk496I5IL8LzxJodero2JZti3cBK0IDNYxq6B/+AXk1G8JPwLxDj/RklGm4CzW
7ZrMj0q1fgIQPpZhKQlGvJmSYsSKUUUMmqRRpamnmvc9Qxg4ciRRaQy0It5VrgGkXzx/aqJaXaZ2
Dkn6CNIOF54WFp28kvKgo3aBLSl3m7RVktp6BZ3s3rlPf7+fIPhcpnbMVomkbt7HwnLOCZRWiGta
zef/bQ8L6F/1f70ApIIMdq3YWWoKL7wvLypxyRRLH1hzh+yHZ7eanCEJUKRrekSKFcf/516NPhBn
9LDk/aVANpmKMdmOotMjCloBsaOCKBnNeVrBwHwfLQU7EP4rXqDB8HNUTs84fK5wtMxxg4JS7g+n
zqoVznm1Uw0JoHtgd5IqPISsEBdf3RD3yiB3M0UIyPAQmctzBkXOp762xSc3a8EximPMba4Ef8dF
w+tig9EIPDaasXNGIVSsu6sqhBLLCMUb267uy0f/jLKIUVnd7c/oXNE9HDAjouq1Y0/d0L9d1egb
onWgcdyft0VcqeI7X1AkZ7kVGgrjFIwiYnvzVmmejD2FX2IX0FS9/VZcrqaDfT214IE7jLM9RKtn
d1dq711YmPr6kw1HYY5zbszgOVtBeqoo3a3XkCKQucwjGFGHOiLcD1895x+6WF1y4FFlWoyRV1tK
yqG3VLcVsNz8tLCi0MEhg3fCq1ufVsO2J1Nvs86Ksf9uHBq9tXoAeSzc//WHlfxzbR8WjN5X/OBT
bk+eLNLmAdRsAP68gzn2Y51/5rSN0Oj+QH4qDmHcNNmzOaSGWnfi3meu8O8gq5U7IjMTPjujKDFL
A6w9merSoM48zQSKp+Jkeb6wui0yIX0NhEyo85zos51VW7tHuz/9H9K+9ZR+o7rlMo5YrvzPwBdI
4QWF0g96FkQ8FwXysf7RnOGvAuVj8Rz7ShS/BrUvAqy2yecFgeRTXASLoDFdTjjEcyq9kn3g1RTH
PsI7GYeuqggVZllvw2i6/Bn48gQrqToLirtW1kqmfssJZdfGY1dzgzzu+2Cdtu+/u9fCqxHGlIv2
uL4oppYBk7NcHAtlls2CKnu4Rh3V+luQnLfYkLBvY+5VpYsxzGHXV5cgTzKI7G2JIUIQDkdMCTMd
A76kmgVhOm2kqO87BqzQyE9GGWuk2rY6tdkrD93y+SMA4LH5efRBZwsvBXaGyeaUxDxM7H3qC/xd
TdhnQRQ/b7saCxnZ4OHRSYWTIRV/uYyKWgiOM+2m0qBKC6cRB/6AbvxFffoR+kb/unXFt011XWVl
GlaRBL4jXQnm+DtEE+fIjlM0TwaJMqM9KuBwm65SIVNgKQV7kqPa7K+F/R0BqvDVl59t9pcG8Yey
N//Bd0BnvXx7CACWsqLJRWrLzNVbSNcvlZ8o2EZddFh7eNyci9q8Tvjyv7pHBoikllikQ85fod44
L1+voYc+Vc+2SE0uGOPcgEVodar+06dGINkghy9mIfEfnlIjvTMQlLSuCxGjeuRHSspmr5m8p7fN
KxZpPhINCZpSBTVt4c8x0Pz61y12SyTr++ehsLa6qgHVII7ZD6ra2U7QnVD6rZwn1DwUB5hi7Jnc
dvIzaMWkb1JBR4U/uqgwwGERlDeVPa8BH1eCoWtqlFwVDjF1LasFR8sOHtWYqjwxnbs3XEbETE9j
IwxNEFgAUut56DqwtTxRdkbM/9/hU0UcFQ12tfg+q14sWl4NTr7gb2CgvJmGE+2jtz2rYqlCdTiu
Sx3fdB6Lja+FZtse/5xGeCqktuez58H3ocrIjEOgVirF6k1Fz2ArEGzDOyA55ni90xprTroSElj4
9wMrvj6xL659jF/Xc9pJFAw71uTQVwmJRQ1nedyb+IUPxdON2Ih6eBpJPa+WwcrlwON7vK1hFUn+
eGRZhBlPy25A26GYh4yHs5NwAMkaoBcYxA7FD/wSP3TMGzpR7Wx2khxQZqr+4GO9wHDDh6KJ9b5H
nD7WNAwwRHrdR/XRCEbNM0n69+x1GIhWNEkefJicOXoYNV7DqELeEIh4HOR0nWYRVbMXOHwZwQ78
i/78xp+KNSYmOUeJkTOOGiQ1U2d8eEKqru81CWgrlo8sz3dopxDoGhUw+lk40CsIzDzxYsQ0W2W2
JAguiYqJHz6EC/ZGACY5485BwE07Z6nv76ZM6pafdlbCLb9aza/7qPWgm9ITkDAnL0TOBb6OIOfy
bFthi/jbbL96+nmvYvWeg0+/21ZO0UBDtN5MFaJCdnlzXbTQ2HqWkmEHkxSCubrcyD0I1O6Bl4mR
H9kgCD+qOw5Q9idgiN6tW5NZVNigr8aywxQASWvcgDJ/dKZgL5v1AZZV344Ek05ebsW7ekWYtbXC
Ax71/B60pYElXfYSKkHN5M4fvRnFdul/El2en5sdS0C2ea/S4LMk0X/OItcMm4nqoqRzXCW4EfqF
F4iVY5WVUUXSU+gcZi7/gNQeTrY/6S9SNcuRKeil/r6W5MXjdphHI6rJ9gSXzqOS/ZOUvwRopTWE
dvEY3qEjyvahGJsGUlpfBpV0MJgafFdEPRzRwNoKMplJjCDrUi8OIAg9LIALvycePjwWW0TNvRey
RtKleUnLC3RXUyiD0g9+Gtic4iXc01Fhky08rsGml/4cXa446YS9uj9zaP4ttvcS5Z9IaQHi2mS3
jxDiFdQmgZEjbo2HAMToIYF94i3y49rV5P6VfvXjJtJQ2XNrUjFtBk3CfFfuMEvxYJHa0R6Vcryo
8ZDmN2pV0awyASa9Tu56JG+nR4N0BER8CodOTq9WHISPvm+v7JDiz/Vm0iSQzvoVbRlC3rktTAv/
eIrwJKXmW22n9iPfxpQ2ZjgwsMl1F08MciQ6Ah9ZvmlNl43JpdqVLsmGDhFyzetpRxDsFt4hqDNu
IbSodSt+g346iJjtbqcipPAfTDmW31BuErSq9Cid4wbnH0/q7ShYATiG0xE44LCCZV8suVNXvsy5
klkuQ7QdFohoLrRivjTIlUEOrrMfeJMGsdCYw0bTC8oYhD4AO4dbBd0DIjICKuJiY/rjz/m2+bFK
k+GlZft7SvqII460ecue82qw/bD2Y7+X3Hnpknl8NATHTfr8ndRPuaZAACAIemk3IyMMvObmn2rH
epTlzxqVSy3zvr2VeGmIjHjNVdhfvvViYKyUXfQwh/5Krxaa5WBNp2z4EwgachoNKdw/N9mNdYEa
Lo1JhRbId8/iUpoyxmzVtNlYaZRZv+E88BwzNVnyLZi2I8DjpP/ym6IqUy95DNDVNZjmtrvtzmNp
ZQPCTiqSliJwYxlVCbXoxTFvkxThhKiWp6rPReK4/L3LL2Buw+yRNliyQgjowzunhduDT21qIvFm
MCvIjM0VNQHN2E1jVSeeFFRGqLT5D8DFahpTWDELeTMwb2vgafy83mZikIYVQWHXlenc9DRdwmq/
VOKeoWZUmD9YqvjsWDkUMqV3VWJYFv0YvhdkIuRta1acpE7CUIUb473oJwT0BplIRajHwf+1tRS/
zp7qsnn9ZiAuWgUw1t/WSxKbN9GH3TAj9C4RUwyNUUJBSW4L5ceFTER608IlF0FkolnsyKf2PPiN
Ss4FYdUjz8NbdVOtV4iFXBNpkA3Ria66HszBwUKHUlRsLbFgqbp/cp4MoBKJRtRBf28vuuBDE7kI
LnD5WtzPrExpVHeAqSVKqk0ztWefCcPUE/PkK27uUVSixdThuo8cd7TdmxJjQaSQ43ZnCHqw65VZ
WEGCH8DkHJWiQlNvRwQ+owOD9lthBbfCPngi6LfZAltmn+q1kVp0KDKafMFIEXk1OSKJz3AT+jX+
PAEzmFlSuz0cnBSdn7EgNePqhmg1wyuHzCGsq0IQgJ0zqSTt4ySF52xNh3ZT3442qau7kQI4AfbH
zmCvTF4CU3Berse5PJtjhVtMXKWxALD2GytKNKJ8lp12jih9ZGvDMX6aMfFnLvF2wfhpAi3X0OXk
hbtn5iAo/yL0fsiDuSg8448/vtfZMFcxsA4Laxika/vgESI+HKS17IW/wqBeOUUr7e2IJxVEQu50
1KJTT6NLSMAG9dV0j5WJnORbZAZi7qxd8xQ2cQ+GuEfE6gXSmNHoSwPyL+d1GQCcDRGzRLpyaoL3
Jw7zp7PVUJppyFEqkpr1eTFrijw6W9dj4V4DxI5Vzwi7URYalnNW0Rf9aJOm214OGfLRcc1ZzpiZ
JWbnSR6mLeyST6n54tQuXXmkVEcApMyxmzQmEzWm6kyJ7QPAskWzPiYGTt9C2Ps4KWHP4VyEnVHf
pnucZoGF2vlhWtH+fx3+cX/pnSZ/iJBBYm52UJP1j3iI0v0wQsOZMpY3jcrLGcCUTEdbFxHb+G+B
q8JPPkRVGli/3JN27adsM+N/UDItf1HMha3AyPj9U0j6AbxB/SF9mDnXqU4bwcgEMCNtTLCxcWpC
/T2JFTF5Em1B5+k4adPAAX7lsuRAb6MK8OY3Ir5OTs2tGDbvVJlMi0otR34rjMizCKuzU4kgYFTj
3tQNKPvobqFuWLteNrP3De2rQWlhxPBaabtLlB9aeES4Zl0vb1xVM/HikGEi/v0XY1uP5ireqVVZ
0397rZSI2DxuKXHcskiGsA8gib5a8GUKNfYI6rEE+Ec7ssuz2lCUOD5dhrQLstibj8xJqUxNJRaG
MpeQqxY8sd7gjJVlOkegXlD6RrjlNjUE3EGqNmKu5YwPDcf4e0akCUVmTQWNZhoXIJeFE75NEXPM
VtrKJpv9ZU9t5XmcXh74dzvZlj22E/5CAbLOeRma1yPuzWjwOJ6KzXH604eCh1E1FproyTQQ82NR
5Zg/9Geg7pLuKEk/38Igj3RaZ6ni5CTXmJeUBcWiWkcSuyjuabvVt56ea0VYEpGrspaQzPrlj0NF
jEaWRia6xQAxQK9r8YVyEdqxw5fD/A9SDiyMRYZLJgd6bQ0nrzL8kPq8aPnyfxKSBsZIVT2m33NQ
QDk2hfbvAAS6hjC9l9Xavnp3n9cO10/v6kLB1+5adW+SEomumu1TjDxfnBnEdotHTOETMiIm+ZTQ
YNkOEWMhQwAlZlV0uC+T7IaEpRVCY9Bnqmo7MxcpMFinUZYyZ5eH9LCEdDT44XQWqmdDvXiBjADw
z+GjkRt+kU4HFJrwSAGS5YP2oJdhcm7f4BconFkjp5LoNVclK7gQL2f3eT1HcfI3B1Mc9ifCWS78
mXp5hj0Fu8cjsCDPwk3DoZZRX2VSByWSQKcwWOGJB9eVZN0GnJNYyshMlXyaGWBGs+hcKNLc8Eik
yXWkryZU2+j1iv30d5F97zm3x3YT0Al2NrE6XZFzQNSqSNZQ7m2ABa/KlWkHLx3GZ0yb07qjMtJq
pRVVUlqnBpXR+ZSsoR1wRC4GhX3XzGTzgGQtLRKJJL6sB6o5DDFBa0M/sGZ+ldtgnJlMt4yGR/QG
s8WSlWznayCMnXZyE/qiiIQW5FAzg/E5yIRPT49ENVX3SE7tb6Vd7+A+y/aof12zyvsoWbet8EBr
F1LSsKkR2820vCNbBbVIkmRHO29qev0LVNyIt6ohIc5FYaoNuQn+MDv7PaNIg5czyubRAF/AtIfv
rE1ZV8fB8yB5MSRrTJtx/R8nkLdzhdP06gAfYV1JC6Arvt7gfOV+kL0uXqj9iK/1/HloDPPujDOv
OUoBeyC6Mw9vCAeWrNL0nKnrIkKyX719qb8/Ixx1y459aD92yLlPZ5fwpuZZQYzvfaxAZtaXpoXx
wCDuOb3ys/vJF2tfj+DBWdELkvPqtxz7940w2Tt86RNy3nIYWGwh8lVqGUlXCkjpozUGG5P9oZPT
eIbDYwi6D4zhQmHJYjFpZyacOIXJ9DB+YjG2yvY+KvV9mNNT3UNnZ+SI3+j2lyayS5zVL2viQ70t
aiW1g5HB6rDAmfwmLJeysXEMwgMf5rgq/cbTV53P4RU/YEXww/swBAA/eGd6rPTg2Qxa6L08G3Bq
dAscjgAQNvCT70fuse6ILcJZTHzxFCf7HXu4JAkHYkNMpysTmEN+eh390+Lg4MG9Vl0XrPsZ5xXB
d+zSge3UgpQ9Zt/GNCuv71tgDnb//m9M5+w5sva3bUP1iJ2XWnxzY0AcS0kU56rf4pG62iZ/AuaO
ny69s1isLt2r6acmTNG+wlwdk/Z4OTd4Z9l6aB7inF0V/9tIF2eo7Xz0/MdBo2ZkroIKR2Px6hTI
rb00TjbirXW2OYdRc3/hB48utSq5soNQjO9tMIh7GAwEV3HI18eCCXtXztdYXvRI4m/bhtBiyNCE
VsxwnT1ovzWWcvSUO07cMctMEEd3sRxs+TAifp1ntnkxLc0jR2KF7xx6eQzmIr2NQUQliH2ViFge
kVDH08leaPdmM9H7sj+3G+mZY92BNEYzl02BzEReALr6EItC6KbCFwhkvhsU+s4JkcFFoAWZ3ikJ
bgRhGQL/mpXeUI+vynoSLRqP6vyeEu7RdBA2N2j5pSnC7tvv8XbYrF2JdNSOrP0dXpLiZqfopsJQ
ekxvAqoRBuWQGS5P4ZLtwAAvfxwUIhTy23F+rCkY6Gz285TeVWpgr+RkODyFgYVfqhcItjWmimqJ
+v8DbyRzBo49dMH8xe0O+mwLkxNa7ARuOW8t7yYzm10JksqzRazkBnNV9yQDfawRFrz/C1jDbxeY
2kmfq1WyIgLEeez6vloOgvO77ENYZTTQoBN5H7ZV+0N7F6WmUHxMrBliHmWg8OrK26aeFcCZ7qqR
rlLG4GG88IfbHnXN00BvOHCU1zHugOAbCn3Ce2v2KpXCszZ9TIPNJnVEaLZr2RApDh/0tKm7TphX
HWf62CPQ5VGD9zYHViLowUOZO2TD8qMwl5XQ2cWkB9t8+N4xTGmPlFQTSYqLLGZ5TRoACL3G1fr/
7TWxs0bjwgzsN2fje6f7hQV4mBhPL+jbQMzu2FxGSEQ4VKCrGPwbaoOeZSNP2mncOMDYuDtsP17o
sd8+F1AMriEgfWRVs2g5NrQ7cIT/HH1hJ1O7Z/SNCXc09EsAf/K5B8YWgV7g5S9VFtmnnRbHAKH5
jJbZNJyOivvDX9OxnK7HKPNAga3z1T6V6uUvp8uNlzIof8N3n5B0aJ8Dn0BRKIAtwxGeX/TuzWNp
+ZO+mi+YXClGk9VofAw3sxX7rF0DEyTSWH9wuKth7CVZXobxKARO57x8FVd5nPDo+clxxXY1P3Tl
sj5XlW8zxhgnrq9NJk6uj473VGy8sJDwQq1T4E9oroFhQqNrtyuzb0zB9BPBiiNvcA8jJmrUOgKU
rDxlMEB6SIH35mjJ977OkhCst2RgyNjsXAwSLQ3FmGqYc+qsix8AKJme7+w+ezW1QTUpc97tnf/S
SAjrQG8Ur3ED+UUje4nimPND4FU+NVjnJ2svXO9aCNy6crkdLohf4lBrbgBtjlf1mfGCu2uWw3LD
IB6we1xOe+lfNphlToAlfZz16jbMCzxmLWJgT99fOxh84/CLzvb26WEs8n2Et6j2B+Iqf/s0Larb
9++2TiGJOVt/5u5wL9ui8jWFZ9/fj0Oq9AYpwerV+raiGTGn81C/uHAcyzjIWJ8WCpew8/9WA2Zr
N4EHLb6ZNtfJYjD7Wc1tIpzDkIpWAuMEVlnA3LMjMENhoFv+sMoY+wKBKHOYKs40MvxygQBKcWLZ
CitBC8r+gI+9ZJ3n2WRqbsbPioz6mqYAdDIksXxsgrbw+rGsYU3Pr0aj/XOr9YE/0h2QC9+1Zc4b
7LfCgyMSD5E4h88GFWdsZ78IQFGpirx5CdiMedDXkoQIa95YR+nrCQzaJoYBJXnl2FqgEKdPR6ug
iWpAFmUTrsqonkRo2JkVqjZEzy6uYkq1VIXbfD1tn+dBJJbFhhBDY3Fwb7lS0fLYi+KARp+XFlLZ
N0h7T5CnEDt65F/1IylJmBH7gyRzZaNirCrC9mrFxi/Vde8xs8ovKN8pYUXNWSVQFoHwnHQcsMTh
RRs2dJGMex1W+FzWJfDAnjYzDkJZKRqdLWJzE4zPUo17mpAM5H9PIX24+89kLndjk4WMTN7XmgVl
+iJ6xrRhz3axud+x3wW6RrINk7N65D5M2ipOxtV5lAxi5zE5knwAO8YKGHQc2Xqe85TmZ3psVdEE
FDsroPhqOkaQXOE107NvgvjWZnIj5o2Uvrlla7bnGgs6IJZxNKLzXxJ2QeFUCCIfiNpzHPBVg4hZ
2rxNqt7V2EuvEIFvxwGowJDEcApOFu1IpAnNKwyQWWdzyXZRpKfAcKWUSVr2AalzY9gAhlYtSA/R
RRuqiqjGEI2DUz/cnBk+qT5P277P0JYCddGyQKvII4KIdmQWoxBHjZXzYl6bbcoyCxhzDFHxaU5G
cQ/98zQFKTsroEWVq+px8antnB2MVc5hFMz2ORk9uBVYmPNPOJF9Ogw6z5BLYb96saIeU3mUrPx9
+QboMqA2wx/4npV0I3+Le4QZ/7MprfZVn2jkb0GJwbGDDgyRF5ObWIL/vnO0BCLCHn5GoxKGfbeh
gLZpNxUn8b7vuluMlSOj4Qll1fAc7BnqEc0A8+ZRHfR7Sn+C2jn3QsYKcetnaj99FUppy06cZX6F
+sAo0JEoYrgVxFffswm20gG+ZgFO/GWJn2+3hPTfgWopMn1DpIteTzXTAe87WkSxXseiryma+Kwv
mNWg8DHhweXRc1Bg3BIh6Ak68TMgio1O7QVbHUsfdHt8uV4p45ZfkQFSLL78mcMvJyADfizqjCr3
bz/3W+QrCSu6gIIV0sxXyVZhQ7p5sgKScZ2nDb1elQlgapdVcYhQE39MGPcHosXmcJvDwzgvR1+L
tZMyi/73eDp6TxSDly/o3XinUS8vHAWHB9eaGU4aFQeaW1kQ4/v6O2PpmIvHQpON96AZxBzI4oQr
RQyXnYC95wrTm9p+x8OUon7Jh2Mzez3z591ojMLLPP0jxhzKjtSi+CIPajjUhnKbchwxUrvVlgQA
0guDuM1gAiE0B8SDEm6+2RhBSm7+i7l1Qh2NO+75GDfTSzrCfDdVMq1Vx60hXxGCnFaELb5h0L9v
EhZLWLrHjKEwEcNOlUcDcW5g5Dpgu7lI+6umyYtl8Vgo9DUIpRro72nmLwbfhpUdFMNC5oY/pNlD
stdvg0Xeth+mDFgPbdviV6VrcrUDhOAwqQ3yevnn6JJFYhnb52OPmc+DhBdt6mN0GqjGKT/K7iWj
UuJ1A45j/bWYR7xqlS/4kfCHvSj2ARTGqWJoslyBehjjmMhW88b0d7wC7WNHZeN5kjGjZVNm6bgT
IimUVwo8UdnUkOAtXiYPd5Oo0TVKyro254kV7Qg4eseETS7KWQonCkV58buofsGb+CWdXIQ4Z1U+
6/FOeP/ZHXMVHUyu0cqJbipmkDZbZ/xg2aEu3ShDxfPpeNkrCAPocvdDyXcFsM6X6b9vd4FrVWP5
JVht5gbvGoO5yt0cQ8iNyAX6ZCK1CzBDM5gX6EuIp8cH2J+nGah7lByfdX8N4qFmQV9PEf7jmOJZ
PUC0x3LGQO/iyikW9NiTM4gWiCnFjppgxe5ivwJ2WdxMbxKr4xV+8kS/vpr9OxQ4Y3yu0OJAHQI/
XZwkRR+rdj5arJ9ikBEr069Aqo1HFcb4sev3I3z9CdKKCGl8he4FFDwtaYOfwEhxhC8lsgQ/TEgH
N8uVUm3wC6bgzPNnT/Q0ixvPn1lxyTcqSNLB4BCAAgUF5wfeVQv559ES/zUPdQf8vIeIx0cuRuos
iquGxEuN7zDdx8uBrEiIWmrxJzUOaxaf+Vpp1nQS+4nRpUzifkE0fRjeX1WuEbp8IywJZxqSksqs
FHWN0PBgKpApfjMBP9/9ZJgPbb9O61AG1gjI0b7KKkxW0e+5r4PPeTTl+isFNJ/An/oMEopLiDbM
xQcZMzOXAZfKYyPavtrTDL5My5gvRs5sVmkjyx257CJyeBwVSmUT+rx51Gz12P8Wsl4tHee4P19Y
QMDsfESyRMKWT0UjCBJKeyqeO6Ph2Lmn4p1fMvQuKSAuH2bOv4KcZG+Y4G88kOKeqeN6GmsSYmWl
Ky0ZmG/dvwX/lHiq1jdyWvsnXx2jPpo/AJcmoQeA1S9OWAi5NTBroqqlyStA4/nPVozJIXaPx1Ac
A74w8qXNfMkXU9rtskoLFHzhWp45JywlCQ1QPKaWKAtGCFIFnmGMtOaYTpH0yAjUeFfD8yfT7ILM
7wPNxbcBth9yDx4dUF/nA8qwFqgNcwKy/OlGHKQjX511CGlTu4bZTx5eQwBhfaQfNozMBQ9FkNrL
vcRDyxf+V3L/piOPZ5X+x2nFEOj7YEeGMUEVHntdh4QyizxZH+r/Nh8Ny+l6sYS5CFjEJAE7QypD
dmbvZ3lVACe5l7OpaK199iE4gPtydqfqVsbVPyvzpNWDPetWVc6B6jYMZEPDpxaA/3gSwrWEqKk3
UTvKaISqjn33j7/hK7yACvLbxB1zJOyAROq7HMjFcciQ1BMXFmBx/Bo1Hc6j5QMIvrg2i8IX6Y5B
iRK+7/EHZvPMspOg1AqcgUTqurzh44rNIGRJEMPcMHGFGzqKjc0pQopCkMlLsoLmStAE8QUFLZZR
k7rdTFd0bXYOWQfhoqa8tLV+Pbt2Bf3lOxIjme1wiJFNb9qpv2AwwgD61vrRs3SLX3aynvhysp9A
n5GXAtsxb6Jg3rlOA/r0EAtGhz9L0hYxqVlX9U4dqJmJ0+/pXxitqVtip7S9k/q1j1wg/ShIVZgz
knfyzPIaqaMYyrln5eOWkywVOBrzKoEoeNJULgLlrzbwmUy6wmlojamlJTv5lBv3fgeCb2DYXdeE
crja8q1qVAbsatYtaacShNLRJ6/XmeM46n0bKrD4RpBUeWZeuEJ5hyI1H28V0RrefZrTKtqi4sbi
by4PJrhXpyokHLUy1vdL7F+/xo5wfhE1CZDinZZ9XxvHyW6BzljJrmkyiTR6Y1e8hnIjzdFoBckW
ANr5HKazvBF/tLqagFAOiCvSixup52cnRNoVywdMWcUkHDDwo93aaOsnuAmDfZ4cQhxyJnbzN1Ns
q+Td5JcmXdZ8IuO4NaHrc3SixJ9o62BySqcmsn9AKu9r4M1FSReKL/TuFvnBN9XdCdMSTqEPNOtt
SAzWYc5DaSdF4vApN0mNfhy1OAsumZc5e8M1WojhDUH69/yAT+jBnHjmYnm+V6iUUCoc/kbyBdMR
rU/JAxBuZgSG1E6pKNnmQLUh6UVFFuoRMhfJh5EQMcn5jp2Y2ZHo2Y+IuR7YDeZwWLrU5cYwmAaa
v9tXq4xyUj3BPJfr4Ct1eUhH/kvZKcA5K6r3MypolZ0+1WpF6HGXKlkFrImvbFk0cZ5VHB7AsGBP
Pkdn21+jl1VM8emrBMUg0ULefssEnqjQrbBTLqbw/WfEDYdUZXAAlhBapzIauvVAK4uMMW45aF6I
4nmL+CG+gG8ZAqM6h3aC4o8lgKpBEgxOeRNGwWzUWLswP6haw0Udp6ZTrOakGnNroiQBwku7o+rP
XBKwv/8qJHLG/fQfWOgAHFNQx1m30kvx3lmQ0jTGYFzB9srRPSzkjEZxP+nZElZ1g50k+0uTkY1y
dAtsZCzfmoA4AMPBc43Mu8+dRbFHVK5l4od0DjlQHgxRIScCRReZ+KYpCcJ2gubgVTfs2QCFXA2o
KFjt1f678dzq0UzQN7l6Lv2+cSJvS/S2/liCVQw8Xgi4qgX7lwVh0pOBhJYkZpl65+4PLgVc7yps
UEAKHPiPqntVxjWEIFcDIL1mN3ADdB1emH4gQljFpKjlAkUJsA4WxfAVQ2C4awj1nIqlufV9PMIs
4bUETOgjTMChjtq5fczHwuL13SBR3MhzssuaRWr/TeVQN2zJFP7uqf6dwXjBQ+gkNzRUtnYZbbvG
oXIwTUfQf5WDYlvGTthPgOmdUaucIJr0xIoBQdgnDrd5GaqN9sTAPwaDiKQxIC240+cz/wDTFswh
Tk/VA21vj6wJc5kSgxRQ/aEUM1u8KGN4gvYT5h4BFH/rw+FLMA253SRXfRQXK/WWNcB5MWIT1Vtc
pO1+htFPhqu0N5oYsdB+Mhr+0pdeuKFxlYq9Rlk8ykU3+rg4u6Inr5b7+HO/fqWgPovnlPspR5l7
BY5vtW1czTl3b/BfiD+05ACG5YLRAlMvKXgoDtYchAiNCK9r3sI1Yy0ykW9hXmxhsbO1ky6nYLsd
PeqpVAHTxgLPem65neB8AF0d8e463XPH0qZ3fWQddvW8J+EOK6r1rx0E8PaXzhCPtWfu6CGbAGov
11sT6sEHCaOOTKoHS0oZTcTHg5hshJCIW+sm1VDsnaI069+2XX7E50bqLS6XPjZXSwttjOnzxfiI
vcKT1bLPL8lcvy3PJbFecWA0Jew/D0R2xoud9IHKdeBpq67jP0FJ/y9twErC2qgFIpCsxhPFp2OL
aYpxs6yfrkNOssjdY5+wW9JfgZD94roVbn6IPiLIzxOu45DF4ePViF8TRoq7h2NJQhSbHjV7PDTO
vIx7qr+OIRJ/7px5wW/VG1TxFZK285P7Od8oXIuGuAAl4ubUMIPHevWMRPmEpYHVt3REsOqm69KA
CfyBgTAZg6gCwPyGRITM5mj0T6qHphc5p+hIfatTQCMbqOsRXcziMrviyeguFLr3lkGGZ7QWUtDH
QJqBUlcIXoN1tfnezpYJ4Ci06xkkPUIlErw75zQS7BcdBz0cfB1hXkdFotBFQCAHdQKsJzMdqstZ
h8Cs0PCaoyFMK8jftILA5iqSxTRZ2ZVlil+ciCxFPIFzdyzEbxbsLIkr6huf+0N4JN2mRtH+gQ2A
vTybHtJaqOdzHQYtcFD4XVwIeKqX0hW1Mayl+pU1OSp+UTRKwwlfN43deBW10VV8NJV36xBxOCoR
dKmnuSKhlvkk61reuSPC6fOyfzDdm0wx0ccCbFAQ//1C28JJOXTR3lq0Yrq1EdIBxSHgAJ/JKn2L
wA1oMRG/Vh3zwV7d0DzJHCy4evp+IZAM7mukckADhcj6azfGXpDaJs6Q5BpJxgK8X2+YIFaNBCOC
bImZeqRFGrf15IK+X5BrkCElPCkpU2nUBZN5kZAwp1YDXNFfcih7spa+cScGy5qFjcsV4jca6Y9u
Au+wURddKqw7d4vC1SP6Z/7CaX8Q9Qco/dz7rKKy/9ReqwecsdNATbI1gpZ/d4aYC134lPSnYkRd
lW22vp7nsRSjGITescDNKtzXdZu0jBX6LvB2YaxFagJvNSaZC8YgD27SbGXS4ZaYcqYoG4PiCsvP
NhBIonL+xdzK4HpiMWYiXMZC69NLsjVW2CiepsUbDuvhWNliA9aDe1k11bDUU/u/aeBFw2qE/PYG
5gzrPDi/1KH6hcw9hx7EoO3sqSliDYZnCu943nWxD7fCeys2O5gBxgv9DZgN66Y9/LKkJlGIruXT
n8JPHlsCLVV5PXXZUkVSzw6hxg64WwxS8HY0TI659SddpivxktRIs+qDOn+wOzWyuflSnJTKZ045
dwvlsKPOvu+fTG+/+lz3yZLB/ahE3GC1+INcdcbMG7duXCXlJN7O44ReBgMQIPeMgBZ4hTGuo9Sw
Gjvvb7nMWlqLh4+P6meKtQfNrejaRvqERFSob8zXGAXUJPGqR77FZITKeVvVk9KOpp1VtdINurMj
68iJOpfrJmdMgv7tFYmrtEgPW77edNBm/Lxb4JBmqd0rBK68iPHCJx/BilgiuWKtsI6IXdeVnsgK
PV2kxCdIkWCyivOvdcrMwM2kOoTXLRj5GxKtTHgp0hJ1ziVJ8mH420srI7NZ9QRX6CpOwzaJYA/K
Cuyn4I7N70IkyMV1HXthWkFtlyszo1TFZjBt3gAOGcJA7vvJ4QP3hgqo0xDvJqDwUbliG3h/3l6t
OsZLpi/Qk5R6Deo/x3MkJiKiEH8FW/3o6Z0HIoKv6LrTXK3+JLf9+BMCtwxx+eEcKc7CR4smMyyu
bq4Y9fM+Zk18ct6Q4jXH5B6bkO8LbpkaervsAoE7kB+ZxndA/ulJTm5j8ZRRj6cNhb/gC7bOLxcH
Q2wIL87nVPOj5XL1otnhZ4sIVxmGgWSAFCNLwxhImf7LuNpJor1WfeOiGzd/vWQXwWrtPmzHN7eE
iU3j6nhSEA3RkXlBJ3RYMEmpeRMtTqGE77J2gcCqK7JbOX/mdecNZm9aT7A3b/s53oqPNiqEqBlR
xyk2poTbY9/u4T/Oyx9GCtpx9LbofESgoIhx4g4WZ3BZiTInE5jBMU2yxvB5UuC4OOwLIy88Qtxg
TA+zjAGcpBGLztVnK9np9Vryw2sVeetB96CwRTnCksQcAKqEr7XBYPezYPuR+mOw60XRzsDzoJt6
8pfJ1CCcmZckIFtP3oZr9n+Tddm7IgxEVxQQdXTZL+9WIRzCR8JjRi/Ye66P/FZ5Wqyj8xHNlYlX
iVSgcyQFxgv6Mspfy8TpWDZY0LZzgJyES8/ExokpZjZvz1oXhA8BgSGJtZ0smi/GBbgAlEIHxuGE
CaOY1s7e+0x1OYZas9M3RNbRUcaKdGDK1JKu7Mu3XuXzCEpiYQeugcq29jOAm9g3ak1YrOBjrYrh
VDkoTVOG+13fxwUA09MN3jgFpkcYftOioVWDZUX8D+MinL8n0UUi0auPLgkXc6B+esaxZfp1h9ht
iJWq9Nolh+Fv+gXu5fjaXP+0+B1n4V8Dm0xYJ4vRB6VkTDC4SCAMoVsjwmCfKZSyMSFVtqvu+YNF
rR3uBT5VywJWx8L8qyuqP1lBxrhAPsh1ZZBv4XLoEd16oyu2SqVW6hTTfukVLO2FJEp4MaDJIlH+
MUkM2BUNhG/xH6ZbpBfqLF7nti6m50VKMT2jzmEGrhsycMrnkCgKANE/IPYUZEg6xxVVYmFRTqO2
MUCkecdvWfzEQiygRMgTok3v4DGrMhSdKUiXWfecVJIdHd/oePuR6CVtBPJIiizLk3Sa3QhjBBRv
Vtu8c5kkpWduKI2LW3EtcaQ5JeravrMfBBXKwr8bx3Zwtr1P29KGT0rgacs8y+HrDwnfyMYSEUp/
X/1fhBBmBE+x3wSNCILRr+uOoHNQCnYyyBRVkTuzd9u3LYXWzSg/K4jFNVxS8X/SaMUGDuziN5dY
1YcX2V+bODSn7ab5lgfWJRrkHffSXor5FF4wdH1/RL5+GlqQsUgqhrfqKGHSsmFJXzjw/LBWAXJF
PWUHe/gbBKyefHucuof2Op7vX0VxjCkaoiOhLq0JyMOeONj2MaylJtepjgQyYmu8nMUgW4zYrTv5
ltE8ZmRkZHBVFPCbpoGs+TajJq2WkNw6OENNtuXG1FRG+x63m/wCXJB946wBYVelo3HeNKsA/pAU
OU4Oq17jS+TBFl/g0376+sy/KAiWbTCSvurseabTQrYhcjl/Gnie9Gho4h1Fg2+xODMB0/gj6B5n
h8JZNn7HMuT2qkyhdOr2M+1W5xO1bsk6NOyE3CPv1OtEbVRWI01v3lwrw0yH1m8G1tA/x/OyIGCJ
XxORWbL89Y9WgM1Z03LYiWa7pvoRtkoivA8FO0wXVXfI+dxQbkC4lcVNOb9ZV3TLCeciGp/iG94b
QXtylPFCGsDyv71adkizQDLSUD0WedNQT7bOY89xfeF0nT0tBqO6ZAqRv1h+buhyJQZJqKME9Tbp
55fd5oOVhZKXIiwfBEqZrtln5eI92URyheLm1HBq4nMuSX74N2ijqjW0SH1Y05h07QJfCK60IGWC
T+XyaElys1utdXcvjKdBqWAI8EKSac+n+Mxr3bq6GZTTM6a9uejk3lxCP/OKKf5/8J7sWnUQPL0m
q52tvJA00fbrpYpFl7CMDxHRKzrgSCFZECYNE35BCpJrFHVt6km6G4jyqh3lps/48Rby396f/qog
INgXUdgoBsTfMioAweXemoXtVrHIX57Hi7oTsyyZjsJ/TajLQLjEDsCpHmVF8gTmwlF4cfDLLvNO
gTA7d68HJhQZOaBcfo10Lnh3w0LT/tGTlrhbzPzPhnvbr0+ew24WWQN58959DT/BOrzpEhN3VfBE
D3KxqiT2VVPtbLrnf9tG4XW+vrvoq+ZIZxOltxCDi3smYucd78Wa2BByYAQDVMqnzumZ3FWaWDA1
j96CqODWCGsgbvn9Q5MGT43GHB3/TXb1dQM1aTsz+Q5dyhhCMZlxA8KMuZNl3LSrZtvX81fezjYY
AkrOZvV0rEFoM4yQMkB6ZQt88G/0HGNYbRly9F5DGMOL2vM6d6UQllgHnf8vAgUEYpOR0EXrHPAu
74mIAxH6OvrtsKwK+hyDCI1sspefteNCKFKEmyryy5ARphzgMjenByAPOfO00NaQucuAdl3IBRjR
+4hChG0yJqfvJ5KMkvkNpXlA2sTnmJxi+br1Ylm3VlFIzMJ+JjeCv/HZNOG7vj+cyFiCun9/GIWp
gabp9/yrY9L1enanWOzAk5dwegbsTTL0uKb/7ASGhYa2CRgj+hfCD6FIwkXa84A6PZZI72aOn0/e
U52L36eFD/EDldunKRZ0NVG15f6xLwkapyB3LyrlOA8m68Ku7m0pX+7rjalN71GbVFLAgvVTxDYZ
Hp9uMHjY3Ohz/c9kAakzDkbGFBVZmhLcywfImh32KmnUPFR+qM0edRFSrHLbNXeyJxAq4HfWjgBq
bMf1oL+j7njy4HNuJxNHIecJxKT3/Uj7lUQk1L1CG64WICt2/1oMRGkGnQ7Apae9WmfFoWyf+CMW
5fl2wlBNFY7XdaCmwysg91Cy7IWgGoZnKoeXWeJKn4ZATtwLAxZraVdCRL4zCgsRyzNvcZUboS2g
qONY0OY1lcvm4tWhkP0i6m1mhjHCi50KzNF528JlGA9beEOrodb4xAiYHmpelr1dm4ofBVmFZky1
1w0uGj2RR1ht1Qnx9OFfy9MZMX+NfvX2jb/unYH6V3n4a9m0IPZXgfpXt6H4LfEtn3RN+E6j0SVv
ZSw69m5dpdl9m8nDeBv0xp4Vp7sPMy9w1evitd90QjX2xoNJrFSlB6IrkuUz2JK1BXf+s81cbCdO
Ne8/jJKpbbjFh9ijJqRoOMK2RZ/81tcqQh//GkFWhUQOJ+9+nAn77Y+g/WVlfw8OJ+qk6ziQWVuI
dlV1r+NvIX8wi8XMqBlvbj89az/gG91Fmtgj557IbU3+iin/n4G51cCZKwHfWekzwkjC+ZAsViTS
UXwe8ES0/PwGpV4/KqP42s+rJNkbJHZooNgVcJ3GIZZ5uXs3EZA5F3JHaqrBuL63xHQuoZvG4x2R
zLG8cevEAxkARPpHTRmhH2uqimRknwJ3DfQ2iUV3s0hsDXkkw0LlKKS9Dc/U9I60ha/Vc4lIK6cc
9jdkladbw4xVWhPJ+DXFKmkiQC3dOoWYPITUqWJW43uX2yE9vbtsAmmqOPf9ZDmu7/J3MNObimdY
J9jLzOsGHhyd6w0Yn6xPLgo2UFL0c2cW/Lwp1evZk/pkRaM5AXvbTe1nDi76SKrUaMA8MvKrBbgo
DqzmJgGteqjQ59D25vP8tr9MKXvAbbqhtKM7fygDuxNtIJL+nGiH+EWfCal+rfGQe9bDKOETRA58
4yLqOknK3nldkCrOEEjwrGoR/qjSVMy0rV8Fp9rfTz+Gh3oabG8zVNBLpimj+ncZENxeDo7PVddk
0yr1wpdh2SGwhW67R4Yk+VOd5n9NuaFLshORSO8JoaovPMazhFTPZWULf5ItpisVh9yUTelpDpac
htG9NqFtC6rL1LqRP/mIRdyWwL1sNUX90CW0fUoptAJse9ObuRE+CW5XBcTe/jv/BB3/x5SL9arU
lv5vjEUkxLH0hUd6OY202qUc1dqZNHSrJx+mRxXKamwiXjpufY+mbpGwLLzX4g8T16/7+H+77Hpq
SNuFXSuhKC/pURJ7hUmIAnfPwGO2oWcq9cBBCdMRHdiD+8OIA/hDjKIrxlstefmRu3gp7qHR7Mj2
vwSLRMWBT3tL3x0YqTRB+ld/KvGufpZ+r4UW1LHFPadrICeq+QUP1TO8dvaN+zg5RkjAwKNqtrts
GaNXpM96KeYF7MrgaZxADGSAJvh7weiLRVkN3PT9tjhgBAnqiVvNXCNvflnH87gm/pJK5EK4rEWz
B91A0J/O/SalpS0dtT8EKHQdaqoMt57RKOZBz4vluy8f07hxSXusCK+4maSEtlfb3Dad/suCJ6jC
2yTxfllf7XiNoCq6U7sfI/FZfTzAYUgzToqoLER1AmTtfXl5DK9Q+H5yWaQ9oRI4ns/Vj6Gpv2S4
NgM89Lhg8WwWRx6U1F1wAkuulH5ntGYnejjqpDavEJevTgIyMVKPqGzCec4Y3m2sOMpmBvKzcNQn
6CPqZMShjXQsi+4aCJKlpaPCA/e6f5/pMYqVhR35chVzGEPgx9aJ/cezwDBXiKGLUTqhlOUPp3nt
/eZND81l1NRoqazpOmMhqnjyUjvD6GKlHWc855kdiQlONw3BU6NO1P3vdwlULmwQh8aMtDcNvhTv
L8edW1nc9fLrSrnYR1vRgVktk1iU8mtIm0xNM+cqk3byo3/VC8c26yuPa3ouRHQp5OfdCeA9PKSX
Emk9PnGVBjunfxqeo9Uw4Zir5EFOysaQILtYoBKDhQlgTvEfT9hAjX3RtPMiMfygYM0ZZM3gYtRc
3nFMhq1o344JtNHUJ4zb9TvjRGWGYbhgo6+8INRnjoofnnOcRUIqbdOvD4FhN3JkXncUHU8NdV0w
+8FjNVKNueH3PP3M7NIYOwe6lO8s4O2qyfJVjZACq03BOkQpxLpL4SG0dXJ7+U7+obbaRDoE8Q6p
bW23KvSX+kVXJIyRx4OSdmkAZqYATjiw1svHDvdDzno8l6xl11G5TX5OYZhpmvdFcvuvV5OYgEWL
dClh+dotwo0PH9J07jLm4DDMWTYac11WBBwHlmEpYJ6G8ccSHsSXsfDCSLgndHjX+Xy4EintS/7j
1RdSHsYUu/08jOLhsyRN0E/pLm4vXyg4E5Pt/3GeeZQEIKgiBg8bgi6RQVwdU9cluDGcuA32S7er
OQ7/SHlB4M1asYWRa2yYgYnvhwEsnqpryEgXzai44C3vpIOsiKmU2zigykcKk692n+EGlErr+Z+R
GIbeRt3KYBtp8ykDFp/1agMwWrgKX1u36IiUaRhOXpq/3x8WoVs/uKrvQOYjHHGiN3Y6uPwyfpYG
v81qWF2sIdviBqcm6WWzRrOLEP/lE6HcE83/tvCzRnhtiLHnwJh8xurRexcI50183O/Z6HFLfbBX
qEGQPvBuiC4brNhII6jUXk+vg1AMuKTFOnjyQ+huGAzq+isLiPSh+/wE024x4xp7dkz7as0nEjj6
+YjP3WhZnXVAYG0xCFEd3Bw9FPSIb1c0Ybr0oo+zRmVRmX75n7jWRfepWel3Gjioi7acFg9tJQ7j
tbvZr2/B70whh3+5faP5qVGUMYlUvejtvpar7X7zHXEGbG3sJnAOchY9nFqygGrUDe7j/IrB/Qf+
db/QBGbacmJq2wVdsxYTUzUJUkYoGV/FtgBm+vwKN0dbxBxTTMAD+lGt8snhSdQ35FYi+wOtUm9G
xOAlt9wx6HEllHcnB0KTGw2OunGkX2jKZH1uyoH6c9gZtZ9MOY+xRBMXhkTwTIoOCGQer44QTBjw
PcLsAimjYKxmZ/w/nX0lw9gQsJwyJKVHOoTmGJj1WXCwVEoeNgbYHqiWsUFLIQ6NC1YwbDv1KuBN
x0lygPzsbWxJN1ffyCqkIW+bSSU28lwU0Gmcqh8IPwmTcyng0MJRz7zrKKNI/3nBPkTiTPh0j33S
nwg+lWosB/xC7ZWJWGtXhoQ28e9Ewa4XvpgMgslF+m11ldf4QjgvKWlS/cDJ94yrPZdSNkDZPgfx
EYQPSrVDPW4QVDsg+dzhBqDR+9uws11ELnv1QvLVSGWF1zZzFfDwMjXGiHRAeMKOwCxjqDwWHA5q
Czoou19XF4my29GAruaxapclvDpbul5s1wduhUsPaSOroj6+MkCi4x64QC3NYZ1eLR6rUi7gRb+s
oxWWlHUue9138uM+GyPWvtVMEmnswbE4QyHPa0EtBpbyQWRLyb6N4FZN9JI2gMeNmYLHtsxgIAuS
fNMxPtMDvx6quMDeoETCj+LPtaUiSYK0dwcCEoQmZ/pKPF2Y12V6jatt/zWt5i+/G58+94zydm9+
CauxzXp/qu5fWJawVEtLoM2WGU9qlvVnKJXmK+eKmp7gcEBML0nDNflhBEiu+kSojiTOZNIxUkoy
ffolBRLxNoF31PfEiFT6ZJRR4ihSYQfgpRZyM+2CaMZcN1ZaoW43y+pNj5CMBJSbvCmW1HIXnAuv
lGLg3OYAEvDfAXv5fFF0szgtqZq/Tl5aVS/bLw1DD+WzpO69x1358OmPxlz9Obat7MAvyscUKiG2
6ZMaLHsfU87xF+FRMTB79HExo+H8tJGRO0Ho7NSN/zfhC/dpYDMlEFy9G5MFmwR5Hzqrhfg4ZF29
yflhdY7ekQX2xeOP4+Ie6r8tR/6vydcsMvt3G6hXviVb96YGNHevFNHE4dfBJDFSPcNDWbDsHr0f
ei1l9P/12N48twOhW+vXije8XsTlqAnYYugxhl5tuX/AvA+z5GvkVfsjQ2twrYydk1rVxNJTRuj9
Lm9OhrFim155znyP0NnBJbzKcX176zn/4uk4u0ug3FRUlJCBalTZQq6l5BVQNHXzUzAIAegrudep
VzMOwIPtASpGEKT1AlncmGXzuarTHGjGDnQlwI/qGWnk8FvG4JfkxHStDscTA8d4hDnTslH1DSAh
SC+8G8SZ6pC2PwexlI/PisqSbmq7SonC4U+gPIxpEAd3hDct4iLDjRzH/sUc5FcsdVfAkb8woDy4
c92rgDYBG2AyNmzCUtI5LKn1PmtGk/pkhVPlwX8kztf5vv8XK3cHh1eAAI9Ak6nCQnoTQ6pYipnf
f14uAL3kNpaaPnddIUgrsQW7QmOewPcueVvIIRZTQZ37aIIK+qwjeAa4gWqy1E+1DDpezGJBjbmb
tUM2NAP7S+pzgMIjlkARGtiMSUfRnoRrcKWnh9CY0lBBrHg8coiP4BKkhI3+2iFGCUg/NnQeQry8
9nyJK0mFOLQLT+w+DusleLRtnwBXu7y5+aDnTBE1TGnxX6iliMW0D9HUJcLRDIvsJBxNJBD0ammj
IGadMGMUV/rrichol9RbT/vQwabhHdNGPCkZ9kz9IH5AL2AuM9DFP1byphuynC4LoPnnwpY/ZfdG
nMRTXwrNHgzQHjeVd7STjfLUm2pKCuL0QeiR28RCjiaHSYE/Gvh9wO0i1ud/nlWjTqNmuekg3b1m
iz2f/ijrBRdy8F93jL1XHuEfNyw8ogS/WILpsLW58Cj6jNaacJ5KzxMCe1QfJw85HHHt8greDYye
neOI1q/CVur6/08cHRU1AGpzSIoPd9WAHhmhHIn4/eTzfk/v8QtIBB33yvjD6r0F96t49WelJGSK
jlfrX5UZY5s3fOhVO08lG6N0x+E4A4ODZzgB/9aKRfOyziFKoYugRwPbFV0LrP4oyi4NFRo02CqD
9Kh+NGkehDvHSfO5Dyhx5ZgPlk3CI4TSJae/jtE2RZ6XNhQmaOk5v2ywn+uZ8Ou6/kLNuwlYbFxz
GdRI0JssxSWArn+bcIX/5H4Hq/d7fCGpY5Kr533XnzNGovSeTGKtjTYJtUtEz5IYpbbB1L4RJVav
Wj+dKVUcfnsX18xC7tL9YUFdE9SA9EhSL2rVC4noWxxEeVUyjhtIqo1MnOH3gra6JYIhGunpl7QC
c+LL0Ai6ZCJBqaOXENqKyRoyRshSVV6E8tNU7iPAYsJRwyETVDjQYJv/UjOkf3RbwCsskT7Rlmfj
f3b8KR2MiTx9SXdmc4JQ/P4B7Vd64jT8iu0t/2whpz+Fg/CycolKi3aSqC5+LqqVayMBittxH979
zqzGkjLmUATG456I5GRtoleSq2n4DzcsCHzLsnB+EBLoEdNF8yCl7Dh4IADh20JEqVDmFFdiwnVd
cyOqKax1ybzlnlN+6yPVj2ziTr0m4hnqbjkFdadFhZgPC56aWBZV0G3VNwxcNbqpn8peZ/QS2jV/
k2ocbLcWshw01GK4074BusGOxUnbhegtaDZ88fhAxJcoe5KiqTTZwXofMsANmZWEvM+j3v+ghRGl
05Wc/fQlc0+4+T/Omadf7LCvSF6nGdgLCAwUFPBOLfG5vROisV7BxM8BfB1Tex3AzoAXBV4AfWBX
11ghMtZgC0nD8YAy23Ab85m1wsWh6A/LD4Dp7DHZ91TGByzrjfXdgMm4uzMrKC5x7P7ZSOqRhdkC
reXe93tsuvxsADdeV/P9Ldm3l1F6AWA028XORymOtvUDzotg0AkLoZChX+f6Mnm7nRdI3AGdG0l1
pJmpFwtIRL8B6bgTWeHSCKm2pk6m3YITn1Ooxox4F7jqc21jXkgCb5d8uMaWMMRyq/gabIv622UT
TF1+UkcS2a8rnhuZqG9i/n3H9OlcgkkObHLiHgpVhn74mnDmLN4VnljCoCzkgiLz6QvJT4S7fglY
OI26u+samdOXGKWd9s+7VqcM1lO804Hvdnm0eCOYjfRVcOOisdZAmHsIzbD7by2foZDUG158riDF
rKNUAkWTQSDlrNZU04hC7wnBNHDqJsN7LY8ONsLLM+KIy/w5hTr4OIt2t0BiTqk0lvL6l/0fkslo
D7CsFUHK95x8pDSd16o+vbEvS4XDnUv1KTyShoNgrjW54BcyJASu/oN0lJQhe+mktOiabnovgE6k
16OO3Oll0CjKrHKHkOM6PofbjIcxUqyhZJVp3/W6smk4kDmTovk8656ld5dJaZgmLZf/CK77Nl4z
4MS8/ZxrL+VhcDS+lzN/VMJJnwy9S3o1tEojeyrui3nxvFk9jt0zs+SHJZ6x3q+PbsnlEJztMMw8
wlfN55sxNOwN9EH8dxgqhKZqvCT6eVCqgyxsjyVpPBAxlC1B+kCA8yRXFCpvjxTRhkWCg54qgeaK
o5wSn2jmmUmh7z+ePHtWjExvwdIaHRSFwCQg/rlDH0SeyFZdk2NbuZD27ZdUScq1tTVYHQIl05Ai
RyZqDrLeN6wTr9Nejf1zoRHINpL9stFXbMEPIKArLGrHL7DBxJ8Tvy1Qx1i3RElKozcubB79wQn3
SetPkTDhicXCzeh4UyXIK6l2GBsHutcIgPyeIV6wztzFCGfwolJUqSit78uQG3XpVB+DSMzqy/Qa
aosWFhTJblZGrsnlOkeEg6Zk0fy2emfRPYih0KHsYx6xmRAMrwSuKwrbZBumT7W3RoyYLsjD4cM8
oF121yTDgSvIze7LlcpaWdn+ypklfNzdEs1Up4ZITSKORvYDULHcWVXhDwq/SMN6CDAhnHnSt3Ls
FuVM0zYMwxqa+63mKJuyfLpUafnV+yV6tOlBPVyMa3vHHam2nCvjHyUk2cEYZ+mDDp47oofc/eA4
79gZQZ4f4/WqAig3qK/m752+XLoSGRmrieUt5MFqEnRE8yo2938le2/nX5PM7BiWfSsZ2Pd3gROT
sgtn472Dgws64uJYioFMs4Bk08/EbvYzSCnfQQTDP4+SVejd/Hh7g3FM/6I6Gpqxf4GtOhPNJYWF
mv34bpmEVAHG1V44S/i1Tt5bPz48yFRWl0isve+vvSInvjhF9cR6ViCrq+EkZiGuDfCnVESGU0dx
BNz7tOpuNm5+A11HzXE7bhQxgMGSxnf/Vws4RCm2uRmGmGXfETAyIz2Vbhp5k81skDZ/Sn5nauFf
Z1Jou8z6jq6BaDqu1UsSig5M9ldMmVR7lphLmod80cge/VwUhmTB5woJ5np1S8/EjMU60wj0n4JC
3w/3cd7+vcpbtgYVXqCOMfJ2fAris0Ur2TKBoB/xLEv19lA+HMXLhmCoj0dcEm0iJm2x8dh32gt3
rqJDoMk1Hq2599obfJOWq4ycg4jTi0xhOMjc9kiWHD+U81pHIbtYiUsWZqZz8wLRYHKmqbYIf1PA
kqGJjJz6aRThUP4lS6DYzI058pQxon3q1asvs87nUZcXYZppvpwh9YeOokdB60o6VZwcT1rKUgPT
WbZAfMoAWbhA4U8y2jKMBt6yUy0gb2jaqXg2K1Aew+mXA0UKDUxyNVMirIS6nCFpKwS1kdYeM6Qe
2De1KwbN8/n52sJbksazb68yWLSzWVzIfb7FJFBmnX+E6FOU+A72aHHNpvU3/xmgLDn8ocA//zoH
g/RbI5dDDeZnehXqoXYiUg1yIIkJck4DY9JCZQ8YKoRPVhyn1zlOniO5Gp1GRfpL+aTlMzak8+2A
jj1SE1kr7kTa11QObIbe1Pk3gFHRor2U7K1QxALotA3Pk5sj8YX6ImB1fp0cQgNbF88ent0PC/YQ
Eu+F0OGXRGObXMZ6C/BJ5czqUAho4sRUj4h5+W3Jm70ALbglS5XuUHD+RJyI1EJSmy+5vWk2EHNo
LsTFZqw+4CxlrEzRzAWjkZTevTx1+M6Pq0eVOgNuGzqZjCGb3buHDJy6dZOXcYZOq6QA1hbpw+AT
VVNcyHiGzTs78zeoyWPs+dqgt6L/d60AI8EWZC2tCdlCW5v1ual7lpeKsw7BmmxIPRZQ0duEefPy
kAZRkUXJyOhpJDcly/yX4UJgGbWMmKHeQfhe4UmInEAU7EhFVuvx/xaTXQXx42ahF+YgNy1EWab4
/FVWLwELlYi4hHOSKtJ9KoJp0Z6m/FLoqNbvMMmWBXlT7voxBCr95kpzZeW6UA2fjb53ZKTFPLBQ
vHsRLfxtCh9bkklkavOmqNNKpKQiCMjpCv+2nyBtV+abmpdxyQ7c5dU6eC4rREh9OjOfNEoy/Qxy
kJSU8KaUt6qCha+CTCEiEmDH71Na7lh7o+tiH+EWf1WiNMvIQVYtSJAX58+05flO6N6D32P4KV7e
kQ+iV4z2Zr+vr19RSzvIbXij3k0llRGnm0H5saAFG+Ud7Ea4WpzvvBiL7B+U47l6DbiioLB2bdvk
vzp/HxugPRdO3VzJMef48sNiBLCF8isg93M0QpEeBY+46COXxfs+Oy/nqkk4TImMB+KU4on5u6S2
b9qCcw/eRb2K0N0SpDyTjarodccVwEyIrUbxmB4kdtMpvCFuuV7o8G2pfCO1e4Z4g0J7Pwguhlr8
d6g4TGTml+5V4U1aPW9yomqo2bfW8eQjz18JjW22sF/Unn3bzU47s9gNByRoYKWuq8GyP7D5n/eF
lwtBI/Kxm8SptmymuHBXe/UHxu+UmAvHeAvc3XuZ18wuSaB7/aAute46hLENKT0lc7DzSolpizpo
6wTfAYmak2Yo007FPCxZ2vRATpE6DL8kYkmFylqqxpA4yTL05Kzoybjq0BZZ7TDMGnhOrL5HfQR9
f1uCMOmv+8RD3aL6kKAbugT7DH76A8YFqt2YVp22hUoVZzV0x4TcAOsa1S/8E/Ohneyfmi+KX2o0
9np1GUEiGa1dRbQGN6GR2dMaDGCmZSwkWI8Pa4/5O/mHboGtZZm1BQENvjsSFRgij9M9dxYm3rAh
F5sVO9/riDygrLQRN7wJ95eLtIQK2JgshYWCTC2IHlza0Esd2VBx2kc9a8Z1mno//fSBMFJ8TmMK
U0yz7z2hVRm2juyQRkbxklUmaMgu+JB9CEnw1beykWwSKkD3aSyjd44RKsWz7lpNAdLkz9JEpNGY
/h4vGXezl2Kr7S6A2euFcwqlPoS3xo4qyoIHAwRpevxu+0yWGSk/tLKOJiyln/OAKKkO9TPSioFi
2Y6HUAMETdhFpR1X01iSB6vugXqEV7XVlh7dbJNHk5nrYA9fJ/z/GhiGzcGsDrLIb9K4yb3HKUkW
byPy/i0+OKRbEvP6vbUK9bhH6mro1RyHtpUFo8ZgKGwf8P43fYWwQCyQmEZXsuFJjbu/YDpFsVEX
fQobbuiiizJIWfMZHEjbmkJiU2sDVTe1TpRvFOJNm7nkhGnN1SJVu0scjkBXGP1KLNwgOwkDByjb
kEwIfVcI3/n3395kDrP2oMd6holZB5eC1iZbh0VAGN/zaYfB2r4SF5dNkOw2vYFEaEQPea/+RxwI
qk0q7GgWZC3juVhRfUxiapTxVuTqVk23C+ORzeOlK9lSjs4MbOuLvoS/zUiDrIlJsjLPg6V+PT2b
IxVWreExzwfLPmJGxTG7y30KnGr1pn5pIQRmnY3RhGk/sR0Ofz/72X1shQp+Jdj+E619yuLttoYi
La87u7838q3Jvo+Qw6URVgxm4Il80KQFOKi1gC5A3NNkzNqT+Kc+BZNotMydE4rMVEyxGje9OewO
nY86b+Clw963pe5e0IFiBWZAAkrt8IYS1JNZsmu0zLmz4u91j3bH+ooQYpuHSMw7+K4hxSHzP3Sx
rnen3IZpNfFFm1Iri0JHTvq2rpdGqwSeWwcF1S8BCni6CYZh9uLGlyePdM3Gw4bnOfVetFfXSXsX
5MCBV88Y87h9hHuGa3omSG4fnT1CKwzfCcRlmtJ5hIE1dO/Ndj1w2x7OH7nxlatiFIS6m1UKUOIR
ovywKlqo1z/iKEyn9347Md/Hu/wC0oLXxf+RTK1IWh7SMYPi+fSBSa/HpXeqyPg4+tzsn+Rli9OX
ybeOyWMDl7HqiIkEZu1GI/BkkZONcPK3IWz10vCPGnDP9qD3OZcWvx4v1+/ZX32dlzV8XRt9Wd3p
omzXX2TTpvYXfVFIfZeDWDHTQXzntofIoWzH8UosjdCewaU5EoQgQIm2/B7az2s4Yev0N6F48gz/
VSA6pYRVmdQX4iQhl8KrN+focEmMdu6e3VI5aPUcPIzdUhSGmeS03nIX1Fy3IDxvIva5YnQC+IYy
UEot3ysW/E9o23GwpRFPxWUo1tXa548YkqLuwyrcmvEduy5CubIim/Ph97qDOT7odWEKyVS4DgaD
7H3rPLU/tjbmhqJSFQaKTiPs/j2l65gD/vgk04ywQzY5RS3dCFRO2i6YWCIFfD8CTI230DW+mbLW
Ku86Vbn6a2SxjObL5h1+uW0QOSRjhhFg3CwZN+y6AXUj271qL2b/LiFx5YTD5FVeYRz3yjMalLMf
rES48tu2qHx4704vl+IM6GgVngR6uZC+o0PAlxnjqSDl3arKSPqogC/JtAWmc8xLQWYYxWuwnFBq
W76nzqpIAj24owj2q1Znzqz///6Zyh7A+g5hvvpb8ZFx9dmLGQ3NZp48uvH/PCy14SFH9EoVrQQK
0t/wH2Ua786ny0O41haLX3Gjyh3ymptexYzqYX7vevuMObfNQMCZeAoKx6rw5vL37EQAMOmRBAIK
WtEUHD2vrznIXm3xtBWgBkfuhuEDXZ74IWyjSU5V8pa4TMijVrvupce/6S0bOwJvvMl+joxRGKdo
xK1cwen9stMkaWa2RrtlsDP19PpChoY3lQ81o8+SnTeahN3riIaVfybmScRqdqwtFlAmx01S2W/e
UqVTpVeLycri7Xzc2B+kus6DXqjQjjbI6Jeg7e1R14U82OWctbnMMhTWypzk7Yh2tXVqJpKnOfWI
SHAYNzpiIefCqAn1YyE3xQl4HqoYZgmSyorH6icCBMSqjuvd1Fdt/7UhIcfK6suIJW6EHzxGNytG
6IXgDDY8gmkHlpeyvnv+H8LsPb/RjqOiVsbaqcp2ypDqA/zjnggl0wCC3YleDY9UWIzFOuJ+TbPI
0vtCiQNmuh0HIkSXmW3QzW1Z3SARK0JWMBrc30FqT+B64zKgNasuwnKRw5pQkfHSLcRW4TTpIRqQ
WixfjYjoUaDy4QxcP+AqhKlEUL5G968mAj6kRWUbSwbRmo4BPs9DHbWJe27XN9Ed+I2/FpztpKAy
jdF7rG+HPR+fK+8L04fw7UHTQEK5SuxL14YOVuU0NoI5iDxX7gBDU10Quc1dwN9Y8Ab+Z1JXSwfx
QDN+Vyh9h8XduB1w3vePdvt7ELzWu9KNZqAcYVhn4+/NrUrpdJt5wbW2S3OBeDXZqm+m2g13IRL+
9lsjsFzR1938f8+mzA5ZudsiCIQnurVUWZvLgPXXwXGb5MNyRwZ6B1yKl8tm7A90/5Gr3XC7WA7P
/+uFqWv9YmU5fKnOr3rz79HPDWMJEDuKrKT1wj8cyVkYNc/1CE/uSSFDTshzXHVpjUl65lQJqOoC
sJm6TF0P5kAa5Vf9H71DkJm9grDBywhxWkgvA3/yGfEi4fNGDCH+EfaAt5T0ipjNs7WPHFmzKLbe
9XEeT2KgIc2ZeJFArVYKExnUu4FrBmER6TiE2dNj9yx1cd8oo2bal8JVIfcPPYnDfxjmSyAwGWxL
FhHu129FWUdTIbDicSb0zCEpVujmFVsDhdolGa+Txpz6/cXXHcZZnjVafVBzlKNSF7zl0CL9sEOo
8/7rKpLwBAFl1eZW9lw3OhueblXL7ZIb65aLYv4GDf5sZNAjm5fmEtot1i9bQamWcqZljbGnZuSt
NOd+iyT8BiyDP7nYkS1/d34vyc8BLD4LuWnl6BkdyUZQN7SvDp1FoKfFHA4xrZeAlTyUloOGYMUw
Yc5huNLUHb9Q3IZQAx7R+EZy6qp+UJbTkPA3DPiIIVsgBAS6PJavvahBPn/vR1CWOcoAqCkTyXBj
vctcxRK70ittPnrZaTsuCZ2Vil8GD2+SbPAgdU/GrVfxvH4lc8b1ryW6kvmzmnwX9PjRx3MXJICd
MOx7Oam4FOLi7mawTR2TyIb14zOAOkq9E3qr870ZEOptNPbIDM8n3DBtgoLKTdpE0xFZK7n3E1Bw
5Uh7MMerrsCsqmynQmfyQeBJu2NJ/+NqKDZ6twEGE6gkNQt8T8NvfmEMdzfl3cU99waerzXXj0eK
j45iUP6QAgINkr5fUt3VCNLZSM9++8MT3IoKg74cVAE1+gl1ILaZmvc4ekbz3HBKwR8XYKId73Li
yEzm+fUolZlGbu4LiDKrDh37k5katWL3NXD1SZRnHWzpce35y6joXWzmGkelnucsOS3o2Kwr2n3A
r9uyfJvYVJZZcP4MPbn++THKn2nEuRiOYy42iwphkNaA6GvvnKMSAR1DvCswmAFjdO172AcgsQ7A
DkIl9Ncn6tAZDBablc1EOiXm19yvhibwgN3ootMiwYgpEcGotvBBtd+cvzjsOab0MqKErUVemDij
LlvO1DlyWLl8IT6NfGwDW4t66atQN+JXhvb5n3kxY39ivyti4xgU8tzClE7Nr5hl1RQeOCvvHcs1
AcJjddzCV/Nb2F22vAHzoiyjaK7RhTXCD+5Og8kg4BfnCMscavIiK2R0h/1YqT6YBXaPZEMJKcs5
VZnIPXve10EliB3nl/YyijuotnFjuiQ2dcPCCdPxsd6eB4Cbm/zKXRy4wfkE1mApisKFb26t0RKI
OFabFajEmnl3m8AULK6vfKHdMfdqbiNTVjhqVzw5XutYJK5Dml/EUP2q1CP0pT3tZ7cH8w3XBIoy
gL5ibRalHA72wgREofo3kLmo4m1VxT78B1VTXWaHE55WDsv8H3JH20/gBpmxEHPAeg5/m/Fj/uBQ
Mc80dr+H3tvhXIn6et8ewXBeynhhmEEO4NJW14PzHbYoZpouXoiersisYdvuWoa6V0EuNacTaLVn
KcPAOTwGm+4fAAhGk7VFlrXxp/V/was7cqW9fq+OsySY+GIoIhpTJGvjQF9ULiZ/VGvThrz8uOYP
FLpIXWUb3lDPe6t09H7hO0oBXPqKNDQtVJ1I2HSNe+pJxMp0p5VIbZnq7AcRXZpqBfbF6TKqs7Ar
I7NdgeiS9MVMQVLF02uq/j+9RGpQUFVvFMnYf2PlkM3wXmv2mrLNByeLe30WUKMrK6lf5hAq+gie
0OK+Kk6dtkmGcu33+84i2PsaF17EeV0dmoAJeW2S32kktU9TD/dBvNYflk1j/tY0uZliPnm9oNfm
JKny0sncthljR9g1HcmN4YIPsshod7lKkXR7bPcxYKy/yDxCktx/XxYDWfZNpGkDd696uY5g64y8
JWOUdVJ4qdKw+pes+w3vJUyNoRfSVDqOl4kUGOFLadBOrjnK9MXkyNLnzfgnfsT1JZWhM9z/kTdy
mhuBOtpaW0CfoqOLFf8gehm3i707UwSah4utanNB782QWGA1IQk8h53fjRDnLD+S7UWc7eh0TdQD
GNlvi1KbzV9bkVJIEbXiclthu3fMUx34G1+ATm5F18Rt5K7NX9PwHDLtuzEse1NLO5noTU8ehjJc
e9yjs0e307yy42LFlfOzZuWNVzPa7A7/JiFPPT0Uj9w87IDgQ7Sh4YIOjQ8yOYIFBpff2wlfEm/+
fZLpxcNv6mAHKOPE5DWxTEoGfmb9KLL7MEAZ3vPxEZS7zVa6PqmxzdDxHyRjmxSY7vO5DImNeyLn
bI9PqxgCMTmsNL+Bjmv/iJieVBfkxaxLZP0QNBIDWXA0lvRbMnhPANJRtDC0bWiGppcrG3/qLogr
iStwugTwgVIsoLOmd9R37g4xAhGmiLIZKhuHiQQMOtn98ZUT0Rlqvy2f/6qjQrl1QP3CjCyqy74f
1vnH8UNMpMckowSGHzr9KZjoSPksu42ctFMYwOT9VsTJ/CZYCHb+J4maL8RdoFxyOut7llIGiTIO
QGCkG2wcQl1RtslOHrAIfQ4jblIsA3CMhzr0ac9tQnx8aTENC8azEGkz2uNJWMvKE7h22+QJroAh
vIHJPvIV70VVVQPleo9xXdc3gQNDXbE5XfIEjItHfh0dwESJv5mR3uArko8a02gRMAnzdMixFw4q
EV0ypI/L55uMJSrbvYpBVaWgRnVE5EL04ewV7aQEMec2jAU7smXmj56TKEvMp+f/UDlLPN+Nyvjt
m38lW40WyLNkRlh0aS0Wla95nv8OvvRS0gefuU+UR88y9AAbAKIcGeOTzVeMOxYvNtS7WvZTlt0M
iG8RZkwbh4VrDiGPTcOXLxpVuwLxY4ya7fKnyIH4DKQuvTohCcuaFa8Ub+gdFhu1G5uyFOJLG6+6
xAUNssMl4Myeh9E3qBWRKI8zC+gdEfJ4WASTC0idkekHrCyV4I9qUG17BMr/s0VjTNu+80x60dbC
S8ZaEzr8qDAsORgBLoeGGOYPmIRXsgQI3Eu8orI5vx5SGxlqCNmz5bFI1/bpj2TaTMH8jCqiyXYU
/sSJt8ylbuy9XymsfavlVPP+QA2s/0w70/Nct7Mp8suq4OKyJaqyuALEocPtFrGRH2VF8zqS25gQ
x8SUVKk+FufAwOhqOI+YQu7sPHuVitjqJDaMoJlPlDLObfHPSFEBdTkHDk5qWa5dnd6p42dEaFzn
lVtVcJ+1+mmwWQmPl9hs0yWZaw/RFzrLycvYQPNYKlZ2PxvGbuOuP8FC13YPsFPD1fWNGNduZ8IG
TUdfRyh8WCH5+erGzKXt5KQjc/WClmn/r7FWPm0mTKuVnDcGDfPHVpDmRZa4Uuw15us/2R4RL2Ha
I0fY5GHV/Iy58mngJTse+JM7CiUGlY072XEL0mUJUFeMYt2N4bROHRn3ZHg1DPLPIFT5EfyyRerA
JcupohatNgnwA5KvEYWDK4mhJ99PFkvi00xYmgCCgI+IhMExBXJpYnOIqgsXdUlEXZZ2wXAxSNdM
R7tCOX7/QTvY1MGI8XsNrWmDgGx6HOdjuH77/rIDvMMIqMdjLGIaAaXiigJ6p/l2/o2XYfWxnA+y
QfyYqTZbxoWnVnJukEhNKDMjl+i4GxF8lbeVkTRvUFjlw8k3hfUbMjLZQzHxVUxBWm/TCy0oecJ1
gu8Zu6PYucTTN+TW+mBU/bIKx3VhEsC43jJabNqz8/n3Kwu5rpPBHHXnZHdsz4oDLX+cDuOCVWPr
zG8PlBpxWdHs0A/zqU7N5L9Cp8JL2FV4fRTEPIFdKueYDssAixqPIdTj/VPdEZGXF48dExifN8vU
uNR7wYIrMqxTV9vp9VAuiHDxOWzmYbHfVfNU5o8MY9sYAyMKOqJdhpgQEnRbpLnfiBYU6sPH18sH
wx9wJpXzFPa2hJM2DyQfPE91rFPuTMGid73mIF+6W6+1ncC/qvOcRrr/x/mibWxoPDYD/U1NZVnw
ThMk7M9jTGEsupp+j5gWiGLYTMlydaAQ5ZEGds6OHxOkxrfKsDGeE88Zvm4JF2caxV6SqyBaUZah
3v9XXuxLX/Gpf+xTZIkPLFfwC9lbfoKXFlgPPeCwTNyeA9ryMOu/tUseunjVHuyLPl/wfz8OP6BG
XzPMzTWWXmx9X2KNpLKoTm6f2xxnDMCmKGi3W5p1SlP2/g5zH3noi3HgO/p5Qp9Nkgbz+8DQONR5
TKZSv9alAFV0PMCFAfrUmxTZh6PNy4+dAgi0JxZHw6zOmMxoQpNPk6tICNsZ7CZHFkKE/LlC2azd
1H98klkPETdQI6fbVIoicjexVOW0UQmIhnRnl8I2TJ7uJc7bbACXQSVgaz15R76vxCXCeZJGqkCn
txkcLRdJwAaOJDrACYewG/nLAc4aIM6Nio04npW+8JWP/zq+TgNwjaA3/JrUWGE5J8jCibNtMUeO
ghoWCXh0jc/Zh0JmGCVfKdFCE0TEs9RujBiCLIRa/OHniXmQ1E8LDJn0DKB79tPLYuGwmTBGn0he
HQ8USD2lsqNajL20SdNl64vMOsN33rVahY1dXAxoytRPUUwcKBSnB65ght5TYmAgQ1bWKt0fcqNU
o5grug43vWi7XlfjNpYUue9RCHOxXuauA0523YywgjsUAt+l/rnPU3hai+3V8q4IPFG8k1lQmFob
iv2OwR41kgATYDBfWbjSaXDbxpGXfAyQqDu4AG2YqF6S8UpkJEsx4DLsFP7vg+3jFiaI22YQFDOV
UG87CnPDk9mJyA/ULDm0DtoAAucJeUYOnLsSfvSoHmXLemvQrexdGTJpl6Jvq/kAX+0lbC4FSdt2
Gh32tT6Se02nAVmXP6C9PwwRBLPNoOkrrEWj+5tW4+RZVahzwm9qqYFJRzR0G/VMPaDOu/7VM1wu
kAycal73jYy4ahUf6L/q6jYfHCQnM5//+Kcxgmok/aoZ1MXFY/k3m3thUFQ1D/t7CI401sZQB6mQ
hFAWLXwliS+YBEbD4XXNVMJBowQllORUW9maEpseLfarjwNCqL12efSgQ9jc15d7G9KOotTINBNU
nqBVtaUNL9RlhLwpOyfZ1HQHaSMdanCnxd34DScG9TyM3g9fRptybSZ6NEg4Cv9wAWYA22rqAOFV
rD+EA1DzXc495zS4SCtWnTXtannQw0D4vaQFdbBSVIaqEkKyGg9CzhxuVdtfRnCyfSOYmHwFgsEp
4kG7NLc17ueZIywPSK0svGKW8Tl46LPZdNiB7dxaFmsHxWIZznudcLEkOJR4ihWz5U0yqCi7v6zc
4Ey5k9cYQutdcOQ6VlfCyswkwQz3jDy3qOkukA4X9AxLjf0wTKxvFUpeaDAP67g3iJ/SQBXKaOuG
XSS6/vEUTaxZbqqllmGyvsM6PE2ozHW47XVQsRQ1PmT16igSKQZfkhi/IQqTDJ9Pb653Vz3DFKKE
unMfOcfPxX4BuQPTR0GaxNDMyff3JHeMefCVaEnIpKMi0Te8Bx29K3RbApRrHV1h7Z0j2UhqsScn
Cw5ACEz0trR37FMKvU1t0MvNAUwq1v7FOZa8YmhGXn0pysV3xGmMTfnZoiTvCdwB8aYjka3rlrcY
2On/6a6qlWqp592/eHn+XyY0ZnDbJkfwDA0Yo9B3r8WqGNTGIqb8m1qJzBQ7VrSFc6nmlSsr/ESh
VaReHdeEwGjBPOHocrUhoUo2SmNKHzkBYnoW+gnFO2fyeLyogR9j6KzwFUakmHanObGOeCYuvayi
TQw6EFrIKTFe7HTRtzzdZlXXUePxyNOxSavd4Q86IyO0Sc1ex3YgiEfn5k5zwDwjUxyLt4WDJ5ww
iPvsg5Ff/menBKajXRtz95yDYPP+l1UG8LV7heDX3GbwdN083zTowmV+Js9VkNUZcT3yK7NC3Eyv
8M7ob8RzX98AlaGzahSwudU9BOXq8hjf7cHErwiJAHAYZA4Qb3Inq3ohglxkkue2q3BZzc5qPrTQ
XFMXKVD06zIl8IOTWP/qLFKk7Six/O8St8VsdKjx1hZONrxW6rZOWX0G0zelognv8lLPIw53Kp6B
3wFIfOgOwWzCbcT+eqfNe6VXAAVsvZX8vHiXyLFsJkXFBIOGLCuycXbWXfuJHA0LiV8sK5Gj/nL1
seNTGUlOaEDuPrG0HSizsWW8C838zFwcA3VOUCgp7yjWXuvKUyRBDNAZ/3c6Afg/h+5e4ioBpQt4
L3d4LbhhNwo6imdUswg6s4c08iYIfa4wV698VxVt7fKHMiflFyV6MZ+vyBIRqGThQjyEZbeFCqsi
YzuL6DCo8iFFq3VhPz++P4ADmvS8IYatYv5FaILKHp9EOoHUX+BYNn64wZYLHpbBWTHl6RXBgMCg
335fCTe3TBa3RcWyEuTyPtPnDk1IEy4r2HvnvaEqytRj0PczOu4MPxW9UzQ4XnyBHr+2GW4iUcBm
Ewa1KIBHTbenFcEX3wHlbXjnRj6/rbSm/US08fWK/xR6V4NyjL9QZgikT6KZHu/Jfe5iAqCUdoaH
BOa1KMeIF63rAcx7VkbnmCY6APKU+UQj4PnHfdYJ77nlnPaHj0FrbrWNz2ExzDJZLnphclzj8zcX
s5x8JV/ywpbLSI7ZXm4Qq+31oV2Idf6E1YKkmV9DPLbJEcmcmklNcoUegVrwXBc19qSM6t6OiC6C
2285iGYewVDsmxJTnqrFIdMguB5u6hAOjBxOMLQB1FEx5ZVpeu1HpEFstJ59nsbSy0YB19w4+23M
NJyiMBI+vNJASZXWmkP8XqdNkXEVKg7s8mcBMSoVfN0GTU7dr8RBYgs4ps2jv90e8KoyvnjYCXi2
P2jGquc69Lli/MupkK2ZrZTbKLXBb682BOqU+t7aUPvJ58/DAtpE4WhUDZ+7xRWRDNsKYExFkahW
+T5Lx2IfoHckLoXGEJl9XeA0EnW6MnjQQ1BkY803N0Nnkll6sl71n+2pdo9QoCmRE1TTTmbF3gd5
LhkTM5F2UIV5RhHqyfgqrvyWPK4xXaYctWvr+2zwO0CHkwXdhxb45baYdQoCA81QL5KLJnlzwd0A
NfepA+/+AXabrRikHcGyI57NOfE5FrJfbL+hoWjUh+1kqK8Domt82X0ouNMzr6wRkFj/ZlPucczr
EoIW37Ut8bqSvLyFMsWUU/DMbMcbolRyLD6K7zdTUadwqDWEa/UGq9xCi6pd4K5i/2Igt09oIqqk
DN2W3NHriM97qk4zfFQqPdqtrkP11fkHcMVVYXOz69YejBwEWYTRyaox+VKwci0mQuqr6SEta3VF
ugAaF6h0UbtVHS8R7qUYvDEcZ+vkBHka5r9KOyD+6E9kLFSDaGfq/wrUJMc9OOs/DkjFxW1grJna
yTFUgHSJ8muC3gcR/QoHZlOxh+vnNlO7U5tWXf9O1A6CqaTA24MswJPGNtBy87tomuPHwI/ezS/w
ex+bZ2aSEy47CmRMq4ob4b6TkqPcmueTUcEBN5PyrE35mEl+Hy+wjYEfEVKdFlXGoHLwnplrezuD
3vYeO2d+tg4IQ4Jby4zlnWQbWdALfeE5rcQLlhAn9NmCRYuWyDcr3fFmAgRPS4gUkiUlvd91kq3c
OyjXXGxJ1+MY5LyB/y7aAcbz387iZlfJNdL1wTOvzZ+axtrdN0IQU4AeW5XUYSc2y3/AkoQmiBlw
pdclsbdMLnCrVpWA/bIyF1WXRptKpDhRX27gPOaIbTHjKU/ww6dK2MudHFhRtJJ6J1En9TxRVLCL
OByHZ3O41lqCStJtjuC8lEaW1HxojcDIAEjS7d9KjSYfakmYF9HSdgvnAkyTjW8oH0+iFoCXvBg+
QgqhuRuemYL2mCORIZ39veks8TSTRNenRqkHKJBF6oAWgbNtWNLU5yEEuuAw8Aaar3XVikOKODCq
wRp7GkYkoyg4lwhMCnRUQvkvgu6jFFh031NqmlX8SShMxYNgeXFXn3TXBj/LycZKQD4qwzokvkrR
GsOcY28w82PPx/SyE8XLtWBeG3hUBuYK1C3/a5DQSnrULkKybRtf1QRzJQa84Lv1s0irm3tcIagQ
TDYfGnu75ueqasBBi772hlAv8oZx6U7O1gfdstoppn5mKwaym925TOizvxoII20nMFzB9JUWnPnc
dwHWQ3Pi7ByhDvMSVV30ALCeOIc1WyBPTbteccuxje913iMm2XF631R+JeSgI1OO63OPj4KQ3+ya
cWG20KRU4A6Wz4ncS6SYfuDXeSVk5OxIUhQ6kOLUAByryy7qWpkeqJ16KmVYldyI+d6Hk9eLpOVL
LXUNQQHTD0AwuCX7iIrx2EhcHIoYQDhZDvBn2J5m4J17E1yniKZAA3nMWMliWhRk1VhwFg2sNBCr
X7hZgqf5eUQaCSinBlmxt9OmrDBz3z0tAanAKVJiJeoC40gPrD0ixW5/m2ULxot8nnmXTXfNLMFu
NhR1GSu5Hh0DwhchyWBYqeGcwdWnhFA/tiyfO3p5cDETjLmxlT8XZJmP/3e6sYiBRte2rUSsU7fL
WK25bLsoSzdarw0Wl49lnoejYLBz7pud8mCl14ABdTKRiL8NqGCAlsbTqxE9fjdFHTSHWj0pRObZ
AqcT9+HEf/UZePPYTdSeHnk7bKTFlWk3AniNUk83rGxRDTWyGdK6X0cpTKW+TXZn+URIRQfKDWQt
tielIBEL/eQssCrx8Cphr+A470q/92AqzmX/qJYPjoBQx24Q/v1N0XxH0aToN+Z4qC/EjkKVHxte
zoBzeqVtp9RWHyWvatK5lRK+wNWIMB9I9yPNzpr2+1dtTIVKgXTYlYLpOvFnCYEGud+kYkl7ST+o
WuUcmfQX52j22OqWSljnEcmiTVsLSdoJBqOQSJ5QlTFwEVf9fpZV3yi4MqjguG2GnYvuw7DYJ4a1
+zZBkxrUZ8I2+FewahMipOc4jldfbQILt4WnEl62BuZ9YswxBQdNVIKJJ3sV36a//SR1PbHUCMz4
cvlfbL/QnI/S959c9oYXmYq8YBJ0DDQkGYIIqGWNnAe4fp9Yip5Jq+HchOXyEDTXvP8ONl0jL3Mx
HYOqLV0MQYbx4q6oJoN+OAFuciDfsRQ7TGr11V+yaN9H5IM6mepda/PmpIcU0/wGj4hJuug5TfmV
iJrTqWEGWyag02zmtEBKemiF5HeC17AJskpYXac+qklG1PXF4qkM3i7ymCNS13isbxSH13FEFcLk
SAsezsv8bcAmq0UylQDRvPHuIuiFM5EQXd+ukxY4hMMOIGlIWPMCfVFxlo2S3y3XS8m90B7hI+ER
95sdlakJGyrfRY5jscJMgIB3aEBzsDvDNjne2QIQnML0pYJuuFzZU2ruSSl/8EIUpugeBKBwZeYY
5XLVy3Ul+cO2h+tzRZUmlixMenrXhglLhv6dbIokJQWJlmTJFdCCRwBnvhe7Q8QTwFqBjZZOeDRl
asuVu4MXS51w3CRrqbe05Otyfknf2AI0Z9lOj/uTOpRj+wjPMsDk7C/tCA1micVRkWA5JBGH9z8M
pGdTmnZpVFlCmmYC/MjZCAkoil2IOJvr/egZ6t6+drH7Y4f/2kSG7LHxBBLKTVq/0Tg9lbGW0fZD
f839OR5J6KzO+3Y8Bmo5wVRPtbc3hIjD7LO6SWuccPEPmkn+ndreOeGPTF6VVeEsvVjdnuuQxsdh
giN+YBoYmNsJiRZzNkYmBWWCSbShWH7UzUfCdyWFybJXHI0uy5puABhRqPGQX3/6I0cBMeXlg3yv
Fr6VoAb+LqcSsskhZhgWPeg1T+I20Yvxb7gGFLCduWzfOif+Ii/L50vGeP2rohlxqvahrnaALjnm
u+xppIvu/lxPMXGccFGXgeLRY/Ti6k4ynEt1nD/HIQBhQQLZxUZp+Cni9Vn/vGDSGF+KsQPFhyAT
eS4SCu0eVh5cBef0lrpWmSObvDJLaphRzNwFPE17lFCBCDtfNytdEVnpg6pSz6gQOQH4a2YTSkiq
6vLJILBolgun/JcelJsXVkDM0lfEuJ7Ch4I1Yh3K/0ekyQJNZmmt/+ypuPs9ODxxMjqqr6YpOSG0
rc1NlkOa1PC+23/IHtdISKj9pRJCy3GUSZmb4dojSclG7+9C4H8nsHB3Vf7X6zxwcvirUPbd0he3
zAkU2rgiRJKaNNqEvmBB/OR6mtfpdzhnitLCGy1HkgXXefYO6Gw3esl3MuxWXWIee181E8YGyRcm
doBVZr/irKEaaybwkqeimHvgN4g6yOtuOpfWTGYZUUqnpQLbkeXw9T7WoutsGjlmmhMz7MZ583c6
gDW+aTXCCknmwvqdjAJjnWKN1kvwgfFVnZOP0tqUosSuNlTk/plqv3hTcgBJ7eCrtrSdJX+hfeQp
iOBQkXbxB+gRgkncmkthEdvB7wnbII+ANlVIsqR7SCVVO2iVB7mZviwBuXFXWv5zqfgD5jb8vpMI
Mou5NEqyeWRy8ZWirLoy7vqeUc2y+KXGxn88wkzFM6MUd8QxebG5qUcHezdtGNGL15inv/8wrsKe
NYyPGIKWo5wV8p4A+m0bs3KdL7hd4b2SefJ900DrUyPl0euQCWL/1bz92FlcoJD1WJWaTzCheETH
ZJB59lfByLtVnARfflJFDNH0v+3PbGlvCvFA4+3eH7p591VFx2ZeQLwJqj3sJ7FZrMlaVKFEXIBe
3Z6r+3OF8dPAd66jPP6v+PbiouA2hrx59a0/20+DVsetgITXgK0fQ70hhrjHOQDjJ3YKpAYjBYxJ
79H/QmJigWDqIrN+6cT2mUgioBvrx2SqisltU4pko5Vh7nPetapIjAKPKhZ2iBCghiOzF0gn7DvO
RYJS1eCpXTmCDOxofaaMh9Y2xMZpke9MzZou8QweUOeOKLIYORyemM9ZGCRrqMZfGCOmmaEDqWPv
pAdHFR/6YgdnqhbUSHg+kxKsyYSYPUz117cjlxOGtkMOKTQR3Z0oB7DjqIcYrsyzYuaswzg2m+bV
MwotpsL50S+IPu8pU1BBdgD6CcWEjbIsJZ8HIwtJ27Lczrx2km8zNl8WMRrPpOgYjsxD3kFk0+aC
FFn3f8z7R8LU7siI+lGX51xX78TmhOti0GjYApIzO/6SkoyF/GmKBR5dcliCSXTrcGzFTVnJvbHE
y0bXC9tlVo6V7pliy5zSwfXLoIVnw5g08VxeXzcfKwb0Y0GlOmXf/YNH/UcU25EFpMisGn/D9rHu
QoT/m0WhIRDQSV0oDFORRURhHtMfXCLXS29TuHCB3e814wJq/9aLfWZMsLQZihgKFGC2lZL0mMuy
8sAl3SI1on9/V6e3IiOXiH2vHAIYeiZi9bYpSlHoGQ7XZ+9bTsW7bzXfAWxLtMqze67iYQnVHJaw
1KBPFOcoWZbOJoALPFbvYukFk/3NZZu9NiPz1kiWjPqolbAeJo/Ik2ttmNywJRo3VBxMUnMcM43i
r+inKhGokJljr+3KxHZVzJM0WqzUv1TGAna0qBspqR1tyFlvI6LNkbS2Vykz66C6xjd23Wq56Ew2
FxNjk1mhoM4tqMf8yzljI6q3kTGspdG89oPjyDiPSG9sppiRmdNjXWYCuRTXJ41d4uu+6eEiXh4Q
w8mRSEZ+GaRjwn84OjNpvujtKaknZs7VRaZulYi1N7z69nZiVvifaJp/qS1Db3KopoovyIUFXg7c
TDbmXfILJRfhRm1paeVl19zrFdbB8WkcxZH0zJwV0NvfhiLY7di1itxlg7XWMUOCbc1Bb8k4efxC
80enpV+Wms81ZBfzHy90wbl9JK5LO/78JDTQgjYZECeDcDjPHhDn1ADYcfZiQ4i0lF2dHQtqSJn6
qkWl3asCanjPy5p29p3zaSvQ+Upe04yLCYoFbL194XUJJmxBSs6eKwq4sLivI3vm1PNOoEwNMzOw
WUMlKyfSEdedmbA2uVJP6q/j5bJjNjPasgHV640Q5Nf5ofz/WJbNMDJ21cwU9++A0hZvcnzgazF2
msGpJBoe0X2TbqyrUVJI0i987Sb+japrBIViE8g+BqIo9aH0tzLQReai3HvSOmDac6G2YxcSIKFP
VSFin/LKHFoj6za6tZW0y9szDyksgZJGqpfL0NUhz3sUOsebv0+h3SYslYKu9Gb9Rd8IKjOeuOiV
5xtvnvidpYOLce28M1u1dbAn5GpuXH2hISD/6PxSapFeeCsTnrT6MyJ/yOSHOmal4rBAA9ufpNHO
IvzzEh8X9QDOfgCO1qp7L/K81dXO9RFgpqSLL5eo7RFO6d4sMY8EH8dEcuMr57jWpvfXyG6xnITL
TJWAIpTCLhm7AhjZD4D4OMZUWqFO/A3uBQSxTjBgc/nvcToNjmPuS2rw5bWZXb15BlnC5nWjqDCl
xmFY1U/qwxUBafr+anVBbJpua93+qSwa/yDlCoUjbGfTfrNKPrWyGUyVX8L6s1MD8+RY3v3cUQ17
aTb2iJD73ar6vWcEjBrdMJU5zWib1JmmmFggfyOp9O2hs86oVgIS5p03r6pEzS47YMSeWE3jJ1Mu
LGlD6F+ss47h8uymuPO8W4k4V1y4XFybA8MkUAHWsuf3RxZWx4gzR9aIuLuoXLhL+RQ9G2kumjKc
G528AbVixUGI6F1iYQwlXHYmyUQJZldhGmUo9CwizadB89imYF4otNom577oxv6NtQ2BpGsMSZYm
+OveiH5Fcd1qYFhXJCXOXYBG3VMIIX7kOdo7CG+06YekJhotDKrUUkMn526P+HpP5Hm5oLaY/QRO
y92TI25j+T/0sclKJvJtoHkECmwxnjdpBlHjBjSb/cnwxl6vz8cs8R1Atd2DJ/efiIUrsJ0LYeag
Xigpq9ZvA7TXr/Ng0cyUa6FhxSrFyJcIaanS6BqEasejCsUnY437en62NIHwKemFbSALmyVsLeGq
RadbSslhzuD2vwzSsSiU8pSr68go5VKSQjrMGknjHJdWXe1LItz/iJzLBq3o9Cl3s9CcUzB3sOij
S5lERLIlOb0OPtHuh/dJGmIRBE6L9ZDG8v73U4+JD6kMzl0M5Awn+TUZ/XIFepGkZ1sGfqYFdADU
qtCYqkXzqwG4soLasAcD7Hm2mULvoGHFHyH9ixpMWcTVZ1E6LGCOzEzJWCLcsxmh0Q0NgKn43WsO
aVcFdM1fFJscpUxMziplayS+GbcNXOp87bM5H1IxyQ0G5cpINtoL5G4dn2zzTYJDuBYOeFieRIYi
wO4Mtk1H5gT1zZm4KyagsARbvYePInFrpxDdenBMOD7wEdAk+QMYWDpJTX9F4wCxJHP3HJViLUGD
TDKQYFXq5YFzVtcwPK2Mz1Njc33Na/IDlqRIVo6rN2Ts7GcGdtp7G24E8NHBIymC9sckfjrltkoA
theT2WqK7Nn/mjtWcJAQkdTzNjCtmRZn5y7NwQA4F3TGU0DRfW9ukXPEuwhb1ma9b4FBLI4lPofN
LS9c051dVphUsoeDnhyp31MpGxfCXyrMQk0+ObPt+bBy48SEzQrYIfT7/nkdUiadOd2+8rjtTWiz
UC5UraUhbuRx/fwMWAyP10+LfdFE+pRIJl3r2lKzyjkW31MdwuyVsutk4zdWT8a7XpoD4ek94JBx
nnowz5DUaxD/uYGpaI7cNxtb3qnq096TDgCrhaaKFopAzkCMltXLkSqBEDdsrT0rhf+TURFkZu+I
ayKnr50E+T4GjeGYPe9OGzTVARq+ARu915bPyxA1/4UGH332D9Ccp9VrX4BX3YTl3oyh3ZvolELg
G9DLRvHEq0Bm4j/RIHAjcelAJl5qh1YXmbc0BSDy1w2gtgJ0fRklIr4IRmoaaKJKBP8vvGFf0Jt8
Zeai5CBq2HQccPavgzkjgMNjsxnd1/8t/lcxNGjclcvDFhMDmwrgAdceRNrX7rT+bCWurN7vqGX4
f6GR4gF1OmVtG7zYe9WU7vhe9C1NAoZ4KUtNyUkU+wbzhd08ga3Gcq1ure6KXTIeCiyYgA5lUL8S
LwSO7pK4226Zucf/EVhCqohaTObl8b0ZbjM6g1oWHR17FxPf9bP6eAl1lrNM98LFwtmGC5DbZf2G
h3OoUP+RvZ1NB7ioW1O0XUMeuwCLKCTuAXexUR+6Ik7cE5g1QU693gH2hGUgQ8jPgnvv96JZeWsE
/84k6A6n4rnF8l1ti3IuTSCYS/Ig/Adb7NUJcujYgQ6YnBb0VFIpvejy9PVHPF2iRcnLRRYRIwNW
JLQO6ak6eHLLDYcG7jSbTL1qS52g6VYH51KnNgewR4DQXRqOrZVA1uHiLtxuMk7nhlKalcdsUevI
wDQFWAYi6Y5XwN5Mpx2z3jMG00UMl3iEyrJRCxwoSW3DV13yaBdYhhGeKt+Ri5tCUutXrSbkaZz6
QAK7QXvLAfUSdxSsG0v7gzRwqW6a/twDF0g+IHxcIj2/GcCE7EWbO8PWS3FHUZfvexD4yBGEgkao
+2L+wytCDHNUgqQcoEnzo/0dZAZgOu2SwCFpf4FivUUPFM7+SqyGqPzPlgWOuJVz5pi8hGQfBiNb
iHZEqag6xxX5PpeCIwiBOJhmmEwPGinkiC4ptk1sXn9vHWjLOxf1zyTnUNllQseAhUpzl4y7TVAa
HiHPBlAcA/rnsCs45YylWvsd3Pjo+WRzyNn1YyKE14WfP0Gi2yX72mBjsT2lArIkMtiyEIU6Z2Sl
NVFIq26vyU1EbIRzdjXwdh5JgjqzXsp8HX3VlHaZvGMV7Wy6x8HBHf9iFwI/UxaSZPZT+RxAYd36
yh79cdGDYkGHx6hrLG3uEdZFstMvqynqKTVVxGTh/sasN2/iS8y6ez87MHFPBLBJRO/eRbd16pIp
Y3DLMThI7y8yzmY2cT8BJjvE+7AASJ2G/RzsMy5F5OMkFcl99q4cv9Cy1Iw6pZazUuBcxFxsaIzN
KWKLyyAAKAcSJei6TxNTfqLJLCVRaAnbaRU3HCF8dkigg8pnhAOSeU7xYKh8g+m92mRXlojNdaHM
bqRxhp5Ad/ggusCKvcPeU6kBg8MEZWCq5Lx1eEb+SnL89xnB3WdzOdvR80lrcPFYG4ycP87hYiDv
lQ7QnW6/6MR4Er+6jL2hfZMfYLs838sU9D134qWVqBhygCWEmY7T8Jr2lc0jXO4tok65dbswvF9B
qkIHhMDC5RQVsqwIqwdrMTydkvajQLWrJRasC2LRw4qNHkuSzCjA8cOsECuG0kwl/pWplUfbhyHV
PfTLGLPEs6jwAGEY03/bN3/2HVXDPMvEjo6YUpcEZOyf6e1CECeHj5zVehLfKQcbLscEzGwmAheq
QlXuKpJ70AWwZPnXnWV/yQD2gS7wZd4j9hQ4o8hNunHZ06quMgDasg1vVyPol65Z5ng46nG9wiPT
DTo1oiq91b8pDrDMB9S/VRY2QPXuvrSGqU/uFgVtde9/R+PToI7EgtSVmG7CWjWOnQW1uKCfp3Hf
F4OBAW5op08WV/YN2OGyiKSsA7q94+DVkvJwlBXWRa5dewRRuZcQftiMM6G+M83mm3Fsi9fm5RF2
O8g8eH4+1fzd38IJqexeHKBNG+296FMoIVuqkk+8YfYw4WNy0b6K9FiLzZtbt0fNHt90vl1eTLYG
eE3J2aeWRlj5eedp5678vSvXh1VLja79e/unfl0huSdpEKKC08KKkCnRL5kojIm3PInY3y9aZXNM
WlrKCLy7jnefrHHf82UrsLWfrrQxUlidxE/ciYCV8TADeK3FmkvFuCIs/J+BhySZY29uThbh2sS1
0AhO9ZZmuWx2jmvmkey2bubCkzspsZWKu+cavIVFL5rawJdm5tbkTqrlGx4FDH/cxML3as32Isw/
MS8rVwy3VIx8dOhqd8DoU2firRpZ1mMkHSd/hKcL2QdDOLMHRrPMe2USg9CMICQycTguH6ioFwpy
Hs2iYFyrCVZh+XC8t0FhExVO4O8mlRUna7HhSzkktAx5y00GMYcrlFVUyDibZN/j9ziblgKnVO/l
UcKDtsO96MfkD+2Wr4ZwkV6moG5kuJEaqsWj+f6brdnbdPt5oW/zi1CtwblCN9Np71I2ECE35TaX
mH2BPyZ1upRozJ5IzmTiE8nCXZZDCIlnknN9YO1NVgoECRjbNFKuuZJRU3tgjsh2hANQ/2u1/E8p
gHsJo8Nbxurc8HAhVtWNRJa0PANxbpee1V6pHxDnPQD8Senyk8gk0qC6Na/j8lllNaROwdiTk4iJ
W3zoqzD3Y3nzn69FT177FefqYE/vLqYkhGFUI21Bq0zl0c+wesqWkQ+TuccHot6GtsoirFy6V/N2
3OVmyaMQZ091CDBY0vLculu/Z2dUZJyYC/zPSRiaRUuoY6L4Xc9H5J1IliWbneifrq24c+wIwEXW
iZSIQEq3UcudvYhlO+wKhQz8Yi9f4/ezaH1i3e7BQ6qQ4qwCdhJzx6KWWeGVCkEnzO5B19tdV6DM
K6oWycK86FhD1K91/f/dIIZzl+e6C+IDSfNBxiNh5OlM7MPj11iWm4CnUF3SNjbGbXWzLRgcPSQ3
T7zdF29x0fYkMZFv9fNf6Wl8cSqp37LUVofx/PD9o2QNQCTdxPjPgP+wrE0Vk47M6Bh0yBArkwus
vz45cbmsDubcoJhFl1kLseBpbuYAQHfJVHwOVAI4GWj/Fz0G+7eTtRWPz1qrHOQuFivZy/zygVvF
Ot0Bt8dDz67iR5ERUXUILv2f0eJfUjAUPsejSatzhyj0ielBioeeUIWuWrZUTH/6loUDvPwd9iQD
8JRKBSpZ9ORQKeKiXxQ84CP7XMu8CtQL/hjBELzq9MmlwtHPL8CHIQ6bJmrJMHgl35QOvSK+7v8w
xZduVmQFqjkmFIqvLEWd1s1B+HieJ/Sso8xoqRiV9SS5B7/ti1v04dADXSukwjrOCpse7XDruVia
2AGS0/LNxi0OkIT+kKGC1KARHMVqNX/9VMenLXUO867Ds39SonAK4YsMiQxJoliUyvkE27XTCOtW
UVqInocrK/BjVuA4LBJp4jx7oqkj+SvcfOtWlkbhel3tNxiW8pwc1IGGrV4A8yAXhFI7KAZwc39E
MvhUMhJ6HGxYMRb00v8OVfax9m9Z/ZVI4K8u6od94UTTt0aII1eC8WL3AOUlxNNz3WryhGaWX/yz
dW5Gp76hHkLc9SVENN2wUnc3/H4Tj+j/OjQkEgAtrRTCtKOtsEgK66+k814VrgT9UnNFvxyCB3cD
hkNscDKHyifryAhnrZ6XiiCAoW9MNMdQzEc/XCgabcBEAveVsY7v5U7+E9bdNZ7CDILcv/POnbNo
twK5tMaFN1l21nLWU3MFQVB7caPtQdfxKAo8MKqtsTuhxPTC+XEHGNSZJSLX5rXMcAPMG83ldELQ
fe8K5/+K/pu57jUH5VU78hUYBECp7kbu2drmqY/7XsiqXEAuaUrMViTOifTQ2NjkLIMOl3plOUPn
cr6aqWUbZfqBaXfp57A0cRV8M5xbXS84qQ7DSO87xZ3MZ9SPi265G9OgJtb5P7tByLsks43y3k7R
kENwCiiBwPO/VjIC9BulGFJxs0uiO7NHjvSG6iOSOyJGi8qeB26aCVnQs/2hzYX7FOyyu3RZm1p1
11I48lCp9UD3cBRC4q+h/+dFXNy+nlx1wc6wz8DZdCnkHS76xvUyuQIUoAVfGhqqFbXw8sxsQmVP
CsqxFZpkFahUDGdMo/eUDXUizCmpNkysXbJ3Wo+sQAdHsfF/KT4ApfZceiQ1810/GCBYOYrckz+C
SceFCcl5bLgz04m7nHf3BrdbWK2tD4hO6/1fpdJ4GT5EeHg2V9jC94Pn2d5G2d9QWb8SVT6E3hD6
Ntss3tLN50magGc4GxTHGNwE/tIsRkA2kwm1t2SpK7Uwnz7DNVF5P9xmsQ6xDQgxXm2cV9pJ1YOs
l47zpNNx0HJkp6WhEaQHKGfuQxKZeLWN+oOsx6qNfeaLOynfUk9wr3APOT9i9UbE6E7qtDLxDT0v
tyqRaSLSlKrFQjYvYY5Ayri6q8yyp4uIi0jwW4dYOZ4LFUI0K8aeu6BHMajebVT6OmcpftuKLBUh
0aE4inAthc+JozcdKptoJTwkTFnR2OjdIgPiZp8izQk2f0IGP9tZnJHWHUE5Fwjgu1RcUem5R43C
dyTDBYt2j7wVvngXHL99NKwEzLEMXo/dmZR1QlAThH6btcb7ZT90YHZ3g2BROFfMfz7ibRClPYPR
Xh2Ur7Na4TldT1ebk7TOgBcLiNkIyLVuaxgV/YJ3HpBhkry0bzBRKdv1gKmLAdjyW8bCIH2J9gsE
HrUbLGVf6xjE+N6JS7dSTR/wT3fSf0+kXh6s72FJIY9H9UAvufZ6KQqRLwtpG4MCz8H4Qdp+LuQD
lDiF6KYXbvy7yzDHc5A/p9fVsLNeTdQMt9LtuhkeJDFxfHJDvHKqi+cfOrIc7jsEb7HArzjFxETv
T2fAcN1BjrK7A+oJKeaU/Mu6cBzc9hauNSGDoP6taHjCmeFhZ7nvxYEYI0xjAU6l5PBits15mSIm
AKqsYntMOCzAChLPhQu83rL4ncmgUx2hmGj1EunA9cgIRa9g+BGqWZ24btmL9NiHGTMaPmwPG3qi
GkEBJo74orBUqIj7itsG6x+B2Y8QNOzWXDiBMDt/Ex1N4g7Ol14AcKshnM5P8BajIuJmweYG4Wov
ZdfTc9SrX/hGrC3toi3SnZj9WPKVklPihwqcsUvDJMA4NrqUJbnVQybk6ruCTtwiE4l/njw+cWAh
xqc2M5GS6hTIXxF4acIDSi9eKeGMx5emZqgeiKBc0wGo/pS9ps2UVjZYfbqVoAJwPirxxTPipnUk
Xmt7oMU6QScIif82t3wVlP4X13Dfp5frF3icxD6No9bYTbaFr1qfvDU+qQfb+wfXLrKCzF2j7WHz
JZUNVK3ivWqBJ4AwcLJKcgEtx93UrQ9REOkpNaNnjOo/QM5DEQepvyzIpbpeMwrNAZytvP+JCcRQ
uD7TlstkmMyQtSa1AJVTeZnLl+orFk95jMUKNEA+6nbf1IKUI7braPLUJJSy4l5aVLo/It4Wgd2R
n6r3xVQUP1bbmTnzdwN5O1BWkIDwySCueoW55HMlnLI76mhHtCPDgZvMoa1HEiOphXycvTMnVqIv
0fQE1dytjbN+JuCxOpEjgXFkWEeGGqroXLacKuIRPc+7CstDX2R9rRpGouatdQuwAym4+o5RVRfz
yUr63pfZeyl5Za2iOZiVDmnjtLcPiCkwEUpwzT6s6qNsO6g20vnrcKiEeYyB+K+x0b2SrSYyz/RZ
CZtTsli3NpGXVndtNvruM8YUj0zAZrngnoOAUod/jIMD+sB1chZhhcuyji1uYxh+XITR9zmI2AyZ
jmvzQ3trvZepihjJlWm4uzikpT9aZf+O5kkTJ/jFtLz6j6iGwzDwgleJV6XuNEY2CoEZJkTPcAs7
1stmiqS/QavtSTPJIkYxD8M32SC2mLoPyz4IJx3KhReFhFrtMJQUVLeAwD6NYnpqC2Vm+4mutXPC
y1KDmnBAUcbBZ8YriFkNMbrEH67OpsAxK8z8LGf9RfHzU2ABQHyQPx/1HZRH32hDt2NnydZq7R0d
opKKjofPzw4PxGoq6ZDepXb6bnxqriVVnCBsGxQ2//FSUU7KTcLx739Ds4fE5HbwVUGUtrixxOyF
o7cWL0z1MpnJ5vvmsnSqZ1FcffIdkuwk5SuSE6yDnlYei5K5QChkeQd0lgqjq3cAGb7nGKeFMinK
qSSUgtYuOL3cQKlsxwTFfV4Rt5DL9y66nB0wySxxUiU7uOTfCoPVtLe0AjAn6vNCeASrXvCk4xTp
HNTmjDB5Db6VVSNswh8kbcp3UEnW0RZKPfzmO30yQ8S7WmEAxHj6rURp1rI9Wioa/91O+1Of0z/8
WfUgJA8wLralbitcO99OkthE//f9dAMBxucbryHD0ILivikyAMhySfLrE8hlK6v5nQ93rEbPl+bB
y0+Q/jNLCiiB0B5rMA3nytcGiBGFqKhaG//trnVTuXKABCX6iFm1u3/+4Uh4miYsYsB2KizblmaC
CyGp1XBtKWjdLSOMIWJdEFqg0XHToybig1J3pCaRcr0yLJLc33S7kzk1UK5RNvQpy1lTYIUkXTYQ
JNg3L/uiQ9dvYqkpTZv+36R/a+GC/4fpQaVtyETfdo2ACc0TNuMBJ3JypBHfUmbW7WR81h9e9KXu
BGZ7x0MQoT48XOA7oqUFoGdjsbvuOnb5R1GrC3SfFSkne4cM9hlCwFqUoTgdB2+FqJQ5L252gu1i
PfMNYNSIDTjyPOZh53qQnM3LAKiRkMB3+AVcUNkr0PA5Y7ehhhu37SodrLD5iBBe+NeBv7lgsyHs
s+BqjaXDJJ2Ye/h6txIgMyaWM/NKrpqRMGs+JrKIwzz6KOvGoBZs3ce1VyAKpGR+cVlyfhH2WVjd
ZI9KOmEDm4qNX09uLSHkb+EkhPmajZYS5U6t+/54bzEq4/BNT+L7Acuey7mw16oI6LHt8i5+xAAD
0mhQDFTOJRxZ3TR6+PS9mrLqPQNLT6OBNmTz63CbaW3ksRLB3ROmuFyjTOjTkIgXp2dFWss0IuI9
bILTpBcF8WWtR9G12wPTA/bcGTfzi0TIByqM3UvmgBE+HvdUnclN0GjL2olWyoHeh+Ss82JbZbCP
6xDnwdAznXQsUUKkOM6wEw9mh+42Jo6sbyyT5r+2L2EmkSoQkDCPsv0GV9ZB2L4wRdfbPX28BIg8
k8bSW5sXyJZUnaiZYKguVSrv5sOXsZ5f9Mx9/YnlfnEC/qo5vUwKB7h7dP2NlqRwrhhL4jVIDayr
hNiUXxi36SMv8Q3tiVrZOo8+dCNN7OWRShOP9RXKUTC5K+rQVjBpy912wr4wo4Hhe+mfSRHuJCOk
RxUZQXudlHPloak7xFhZDZV872Z2uW3pXSydQQKrPfTqdUfC3mH1yKftYmlMf+pZ449d1Ab6YfWt
FJImcYHPa4ntq0RIW2gMCMPFwSDvXeY2QL2LzUGmDWFHzHk/ZepGNnAe4Z7n5GiYnUc+APw6v24i
kIzOlajnB//NivUKUY285jh1UGsP3l94PoEBa6ScGNy53rYFC4nand2P28bM3/aY6ShjfpHS/Sn2
jcKnZB0MskOW7MOVME7VKYWVHhVm9XDap9M0JYZSIZZLOUzJ+ZRXyQ7+R3IoQkIa9zxrND2nXsO9
ckyjF42r2rum+S/n1H+MaswgFuANYUFHy9RnVxGiyWng8iOWIK9YirC3xvMN1pwTNhNadsDij1X/
gpYdqJtfEAed95OdW4d1CjOCPoJmaXie/5rewGSoS0h+3Ih1VDpt9ya267rlXkmBJitGx6GQK5If
KO8lwqAXbM6MrohBoqVuzM4YncKO0tqYFModAmK65EjTYrW7Om/Fa25PqqKEgZP+a2Er8klu1z9T
kLQvQTgkRdiaLbDLDGeqpjAGOsB1/Srj6TwpJCTpn3S5ZUHVsD/6gqtkxN9Q9BsRjPgOdghzrqTr
2jg2Em0rtEo+LzKik7CP7XSRG4vmFqid+bGNtl0KRsG3ZJNGRmCCV8Az/ZS6BCjobXdlvdM6Oxc7
k/ATqZ/tsfNko63skZIQ4cVu81+m0eOABNeqK8287ovvWU7myxldvk0PExuK5itOY7mMLsOiIhYE
T1LGJogZrPXQOg35EvPMldtSBiIdI8Y8Us92X0LmqOu01swqnxNSZvNQ0ZlYuj7QIRXyq/RPZkMk
fyYdQOsfThlYUPJU9QiMWi+jLcTt28DCf0cNipRNGvvaVvbedehZhfPMVy/ftNcJCgvAGNq+lyr6
EkyCm+zARfi2omR7fgxn+fWefZ9kw6EULMt7WrD7fBK12BF4hhAJ7xFHBWH9J3gm5a8v64AyQNrU
4N+VoKbfsSU3xDh1FIP1Cuhxv4WWQ+owFuHR/kcjGBhRnRFl5ha3kOcID9D8jXB7FLiHUOExCoUL
ci2qirDv0u/Lpi7kExvaxuxXvTeBZCZMXHTGSG/OufQS/u6gKmrupZZGw7aWIQZtsnb+x4j9zUQM
ATNYWc/f9pTAL0Rob1lWSlgfkBkrY7f8nFy/+CEanbJavc2+7loUanTGJkIdKb7qEijh0bQIPQr0
hEqiv9VBWKmSAbV3UhWDuWuKcmJCMKouhHYQeS0Pty47YiokJO7qfaC6xzTVUpwBP4sD/MlqJATT
X83Gdy4f//HiOHqiO7MssJNTL8wcG9HV5gf9WjUv3MQSlRQXh1E4H1MCB5sF8aHSaWrHLNME+CSc
GlpfVaKimzv1KXvE4VnuVHaVPWoq9DzV086fsMBQYCRA74Sc9k8FlGcLZgsBrCAccY1KKcQRGdAK
9ITv1yOLa/uG62JJPaBMv4e2AV42oodWgFhhmvRTGtGJh+vVgbOvnicW8YPFltNkUbsZGtFG/U6p
wt0vV5176nsaBK5qLveZHW+cMfnobx8bhGnqZhHcg2405ZiLGWE/t/DrdL40FG2KmczhTb1vFdU3
kyWUIJJaTaAN/eIClsBTPL23/IxYTCFZZqch8/aNJrT6FFVqDMDovo1+AVpeD6HssfPgmziarpSn
B83DKNWM4leo7qg38D7RfrxkHV323BHGewrUPJWC/UvxU0WX2BHhK3rUgRXk1j43fomQEFKEeXkI
WY6q9nWnk+ciOVhgxblhbnYePY4BOz0EbmyTi4bZC6axrA+tuZ85xxFJ5KnxjuLLauJdgAl5lboL
2bn5TsI+8O6a3c0/WRIwU7XxHQcODEEbEW0FhSS//+coYH4bDQhB3kYmU+WZ8Q3CLOpEQnDLAS0l
onQIG4biMNIWDV2vH5e5en3FYWErGDuAd+Xxtuwtsz0RSe0l+uNcY8pAMRBxKRi300rCga0NHDaJ
UnN2uwu7jFtGXLJcAGPJyjyA04KjPa9z6HuoWOUJl/qmwHdJTSV1sVJP+dH5B3QuhW4atxPZ7p+v
/1bKX6UTakMnyKR3Vhh+Ko7uVoltYlo4/vpnQqXdPhx/ax0kwG2Vl9slK/3L2DrgtV/kVFnHDGRS
jv433y2URVmGOjWjTJVylzUhw43+o9nDlSt5aQdO/hLExPI0IgOHegopl7dueFINF84zGqnvR8YH
pGbD/e+p8CGpq02bNalAPb4xw3n7wXwoMRiMK1oTeH75pAcY0X0YOmXJLJDbB0cUMG8OFrgCe7TW
RWYEA9jy7CuUZ3J+Yzsk9lfcYR2Z1PSOQeGPhKTivam4oQ9F9pho1IZYJ68Gk9g8qNt8RJ9/jzk5
/uGqxNdXFe002Cyt0VrlppW8wlsKvWVzgp9NSzSdERaydbkZkqEpH/ESJKV1k9D4RrNQJIS9ualO
F3/dDJnmv+lgoSajKEHLryuwZrqfm22oHxa4XpqXSrhtwA9Q6/b3yNrPOKDsiSiS6AfAi9K+/8gz
J2fxjMjl7b6vEeBynW4tJxxfG/G/kleje+hsokMEiYGdul4TPx9nJjpSCZDEdNL6C/LDWFCUlrVy
ywEQ6RSZTSJb1iFh4cIMUSbBMmnfRZFudB2ZqjRVJMUh1b640NqNE+UQKAs8FLTObNXIVP711dLi
GXuYWc8s0zAtO5fhat/D8UjaEMvaoa8KQNiU+AQVN3hCtLc+ol9nda1l7jMqe/BKs04dhyEnlSKd
cWy4Y9HZfxFaxreY0rY/U+9y+m80T+dePgpk0yPhPW98opwKF/sQpAY3OXOv+r7DmDt1f2ma1qt7
vQ/Hs1qM1dDwQPfxnKmWbFaUn0EHgiI2BeutOuwGVQjqL/C0HoaV0RwWglrxJaGX456IWS7bKyzH
bMFNIlqjv3Uyg8WFmNz07CZ/x0o3dOLCOYeQ+X7N9QHGrp4p8qpPYqxgSwvRB8o8EBff9UsPqmwC
0n3efrNLR8D5fHklQcxMvVd5z+C6MO32sSwHO6lJYc6GzEQv1vWQEQ67vdKZCA9qJTEGktWDauTn
tEj/ULqWUGG4mf4wDc8hgtj7qb2cZF5PCz/SIqxDQHKGcH0FJXS5N2TPfy64um0+AUO5ioVJ5Mp8
x1m3XipauaWiO7UkGREgHjc5B4oOl1AJ5Yd2kvZ/4XemDZU/bfhvbO11kTrwgQCyUOxXvSNa4eZv
2OuFCjvrFTC74lSCTZP7aE573UjZa6MPT9iFJW05rsdpFmISKeCp31h6KeyZttXeRBk6xvTcwtSq
Bdi/kS7+JCcUujYI2CFMhKYlbnBRB4Eiwna8T6LFUAQfqk5ehp3DjTsd9kDCaMoU15afiR483mCg
5P0HYpA3HGUjI4YDVZKPdjuDLM7SLmP1l3RtfsPyu5FD2GUcSqlYyAncUavDzN4O2GD4aWhuMaRo
jmFDR2VlhkNffUCh5zDMSkbkFk5ktVfkzZ1Z1Onntv6STcn0d7o56iGElchSuraaPmGQqPa0OzbY
+RkeS/A53h575mEKoAZcZpkJ9C1yn0aC6uspU3nfIFlwNv0yU7dbrV4IfjUDe+skCtGATKITKk44
jbM9zP1M50qdnZdK9Fz6Ni0vO3MrsfUiSecP46qHjxsosHd6rvxE19Nj6QQy+zhBuluJsymSlkJI
ZU2lAlWdD5ChpRweqVhoQtqYoJt7PJvEJ/brPFKpBN15DiefPveO7m02mTft6Wph4scdKzUKAPzo
NJU1rqxW/2oSyuRjYnYUaTetIHxrYWC5OPnmsK3uqPo/eOf1VoGhZF3JUobBB3xMNLwyl4GiwRwG
y0mVxYAlwLkOh22a5yp3L3z+i94tNVr+JtCvRuFUInyobkP1K1bH/pRzbppnbqRHQzgLfOF2eNL2
yPfRs7BQPA0sOLUiyC84LDW/FaoYRoAKJEb9lNibDp11Caa1FPNHIf8WCRIY34ewkH/d8s5pTaJr
eYGoujrA/TW50VVjPKld+mkhutT0TP81FGurVwm/aekqCqMk6UfY+GqzyWi3pdKpAvdIGxbDxdOY
CQi07sz/b36y8aq+A8w61nrUeSlaTM9PINhTk6qkrPMh81WNvFfgGT8mFU65I52ZlA7vUNDiDMEu
fxFU6ECZW5pxTmTik3TwxxdzFiPpmlZfMOzHv3QLIohN3HWkw3ATN5Y23VpllK3wsKwtoNFUCcbK
JdpCOq/ImZ94YyAO1yctPb1ZdBCYYvV8PylPWTFO7aPMBOBi81GIerbPz2gbSDCHZMZ62DubTX9Y
5zgPBAz+KzthzhDU0KT8U4yKy0FU0YP0uR4UAdm1rPbaswG6zd9wrjId3Artz6cDyiaaGx2k94ga
gYzmHvv+8ppxtTLM9werbeeb+XrOXHgIYliGMFWftPWNg189yql6O7ZarG6iUFG7fPrj3reukqZS
jFkEMeGxTaiKObk68ZH0fZQyJ8+XDFVo0nXR6vou84ml8W0MWGgmBPMb7c1Ll/mKSND2nm8i9Hig
Fljk/rYDjXDrpp/IC6U4h2DyuNl/IPht6hOsXaN29v8MCQOIDEIPESMw42R99fxkt/BQ8Lvqj6Jm
hgLhljmPcRbffTp3w+MOojBRQqZhPoC6d7KiYSd5NhMP1DtImgCHVL5KBmnMSByqoRPKm2bmxMG3
58fTYItn3qDst6LrU7Ur7Z+/udyOoyDJfgHgXcPVBkVRR9g9q8p05q/bnG9ri2z5hcJTqkaxP+jD
gLN7y/6ieWnDZJhqcH4ai+5zVWFLFaX+25m9EKMm26eJCQrHjzAlyZLDfR+HApjaLHHkijcS/W4Z
DkC0tP3QZYM9Zid8R9enLHkjekFCA01Yn+c0H9qChSiD8DY0FbQ4sSqxdRzNdHD+vc80sJnvi466
aCyQNxKSFSRmRlXL521wGrIgEs6BuCWMajkb1OhjYR8oRnApM23XvsKwXr5GHiIjhLpbhX2CAt47
lD4V3SBmoaCoGz3Qj9pi9cGNmN6srDzxB0Wg6WW7Mpgu1lmLeHs5eCzbxwZgGwxtPXCZT8aKIlFa
S7Tp28Psjdr3Rbkej51d7cwl8SyMKDSET/R9uB3HC5ejOtJ2vpem9wtom7d9tzHH1Eqabekf6Em1
PmRvtW1Gc9Ko249k/qrf1vKjFKu08wyZu0x1uzqhiegohwN14pzoeUku6gAFVH0Iw0yMj1M8nPpl
FdU5PUKgo/qip3DhrWeLKWumdyoIj3JfhGsEwifX53bLF11IwJ/u2UQZtQCOB4ofAJX7wPBroXWW
z1Nj3KAHhBUMNRvF+oS+Pet/xHn14w1bzkev0DO/DlnP6RznDuzWE7bSCZr9pzAls/YsDjtIZv5r
09hW6ToeZXl5yMeEgpxT/8KwOFmIbNKuNY7dcPep2Bj9iE6WklJYgcy2btG9oaZ5wgFznHXWqWSP
iinzIgn5IAK+SI63iKFGAQoR/ZfJD2QXAnEej0tfNYBsj/CHFD5NBREG29SzEdPcMlWbolZUo0aH
6GOAQfh64Qh+kkBgSLcyqowgjtW7My6azIIpmW5j0XygRMJWx6fAnlaYkhD5ATFOChXVnyI18x6h
Sq1tSa0tWub6P4fBIBEqKxqMXQz+gUDaDw4xgrMH/cgHixXiIl6ExAHreuj5zxBM5GL54BPE6Eoa
J4mEhZgYEu5DrIhShFMQWyxVT3OVCiIO69PeY/1+a59cE0FXmyt73HCfYNneBQc9T5wpRAVKZeYR
8LnNqfCJ/m3J2p5N8kwhyPG5YE/Y003cvbeIL2jec8eTXEDjILLGaL8zdyHw8B3YBT8JlI+CS4EX
4eJ10qHzkUbiqyQ2BOz4SB8N09hG7LFZPG1oCeITk7gpmnWjpXkdqgXe+3g0+hs1ERCPSUrj5/ZF
q+ijuyxl3XaW8GNfQv5ayN9tAcQJxmyV3wFzUGo8kQIXc/f3nawaa72RpvVu3dI08ARyY+XS2Wbo
y+oxO+nGOZmyH5KVDCqqJ9zhEtuRdw7hJbk5h1kvX4v0C2EQHjPNIQGFSOUGw3Z18cmBFHgv1CNE
/h3iC/U/vR3qBKxwEbO1KjBIzLc06l4qtpXMSryjnchX+xZHl1naGRg9H0yBQhlANHkxi4MO9ngz
WrHq+EUf6qJz/LqOm+JbK1YpXn5VQxnzi90ttwouji/aMXNJgt/PffzMDP9e8UObbSg4JQTuh4QE
hprSm0i3wgKW+dYRa4bEj7SJ0fGorRb9fYL8tX+nmAwbEn3gZRgXjI3Q8pPZZhtm//gGGU+9EdH8
keWzVUTZqv4jMkvTZ69A7DNSJQxrqH8BXr5p/HjbJwmySQ9R3bV7zNuJs5M6qfyK0TVgUHyaeChx
7TJQY2nnIBWZRZHOpBfe5lYIVKRDYzU4wj3NrlQXt697m+MgegRsIZxoVEWkcEMqmTL8QP7Dfl9v
nNFkuTiCv+TEYCSPiacfFC+PLCU5j47qOvL6VYhLLurdQCq1Qy9Mpe/kpK124CziXZpjECPsygDC
frJjKu3MJKpLG1j1TnEt/TR35U0S+AFn9ZCNuiegHdIzv1uo2sNeXRNVmg/olEwxoA/0jtqnY7BS
pIla0INNaBmi+MBqEfd3OSCcFmfuosSMvWgK4PYMVZhQ8AS/2YPE5s563ms7PvdS4QNQGHsebUZA
iG2jAVA6AN2yUqI0Y8fH80l5+SJLJLZ/ne2vRtU8OONwgsXEZSHQiiZNCpIEpMsUyMQMWrNrBEqq
OBKkylUQylHaDDW0oDmalUPND0KaytXpoivNKVXACXc/ODnswOgQgXPZEP/GkyKZllKSBKay1Sy7
rgT7KlccHFyi1TLr6WKtfkUAMyzeNiSFhFJ7G75RZRqyx2XL1fMtK5Uj35RAbiufJpRsgs+uf/ua
iUY/iTgiZOCz3+/iMLxnAWOHQfoTdJQCSSWJv9mha9KAL5KvoT19X8Lp4PNje/JKORmpqnLfajCT
pc+GNHQnapp3+mnwgp1TxsWbqdQtTeP2hS6pAKs0qCYTVV3kOFeWyrJHz7Z87iAFt12yVPac1Sat
NJ/1eD2kuxeLNBboXJr0rH0Qc/bKIbczEpUyrSqOZxMAwH+r0kDGHRFCEvQAsGvYxptphuul/JIl
xvloebIiMf7nlsjGMCZbPA2nuddRNyuJsEPi3RqvVordfFm50qMCO4J/1lAL6nqDp6CqQiMUyPiK
iAPiQp1aTPnj3Zo7beSaSHw63Gp70IBkv8/prxqm+EkP0wKdjtoJj91UZOw2pevxxGo6Hvq5zv4c
nKTIOw6oxii9XmgRtAf9Wjj/w8P1QTYjrlMNthtswMXSLNCw0xgjlI7QRWnvqcn99clMSN+fvKnU
ZZF+cCqPDpVl1LIKt61SYc9CnuQ9UarYzJMb1g7ZFrW/19Np34TCuyhFamPJrhfebM868rFWm7ps
deE3+MtiOsXwIgXTdQlSrjIe7Lv6Q1xCJc502n0e6gFudmjicOBv4aTS80Wurt0skmqRiPoZNOfD
wOsNp6uQ2+WEQwRF2oNaAdUC8nhqdmtPo/mXJH57Vhw9AGcOU498cIK12EvTtwkGOuqQ6ZjzmuEo
/1FRRP53gG4W5dAC7SntAR9kOgrGF5kOEGbBLojb1IRVbRMTjGow3yG/IHUjZSC3gbr3j2cRO1wj
kaMx69AVAOiWlApgSWHFCrbnXVSogIP9qo/vI9GlZ6Mn6rkYtZjD+ASxLGDnRkP4TSNBGLTDVvDg
I8RMhgXCndqGksjC6pYydVAyYXCjkXyLWNeL+chC1tGg1prUDxFLvmaQfAJ69UaHyIthI9HIQsRs
Tyc40GM5INJN7kwiRsyQQLOZA86V7N4MJjDNST6HpZf28NzaxaffDWA7Ji+hdZvuoctxb7opOt0W
S2mYDpHrd6L49cd3sJHnbe/Og0XE2s4cHw7GCcqFd8U0Hh9yZdz8q7gRIYuiJGuPl25RKE5bziqv
Os4Ve1GxoenjYmOUBK0HywrqR/bMbeVpbwdqIfCgIaJjAfaAy8AoL94buksiHUsD/FdZGGmMwwcz
oTFjUvG3MOcgzwJqMhlj50f1o4IQ+u0z9N1DJGbjgYS7vrPT53qS5u/X3H4kdbdEvAeIPwg1Gt2k
aYDPSKFszF7DqFUI/JuvCdhK2kWBb5bM08hOpjDfHV6UZIfqOEQ2ri+nhvmlvsX1EOYnCIBKcgqm
oBIXZPKjyplT/V6ixDgRdvDxoypF1Jz4Rm7huc/0pN6Y4VBusyBsqlezj2OY5X4oVDxaZMHDk8AJ
cWORJnHUt57UHRarjq+c4H8uP0XuXcpJLqcSQb60OVACuGR4pmSwF1C4iY/w4PygyCbhkty53DLp
U94SvsW/8qevqOwo0ohNyGczKSj8mVPmKyYAQsMKUhr1ftDZRpWAzilgJ7I4ovYnpsq5tFBmz/2S
kczsERFE5+21SeO097gkoy2FiomwuBMxkdAumL932FIKtduXYSjKACh4S9d4XcCMdn8PNRybK3km
PXpgZPo8ltC8BUsKYseJnNQ8geELfnINee8WdvyP4bE5AstbhL+O/eLnc0cTdaYG2A036KqJA6ZT
/T/IKDgs+SA28sMtehzhBUk6w5xvJ7dtIWzVphYHRe1mIkQLLPLGddeJIay0v0fVNLdDAKFxjpXE
DSUbaKdfRTttl7CkbmNZ9ICvacz7uWv68bzL0KXBei3dMdSvUDw+b7iteTaAK85C4NRTk9odrfI0
uF8LIvUtyDR5vnl8gT+KJlxAabePQMb7n25p2ABNKpLQXiDeuRz00zLkQAzNvSu6GS9PNppwokF/
JZSInkdgxYkj/yhA6mCSz7fPsNST+2yY9AJhAmmDxtGJclpcToPLNuNrAivkvfsXTcwE6PFw+iJv
ssBM2e0WU0uZmRBXMQeloKqXSfDwgXFMLGXcYkoF1y7+Jym7ZnD3W+WyLM9GtNjIAr0RJJNb7gP6
RUsG7GXGluwahPhUXcYpwQCtZB66waHGnVcBECAhgy8P9oAyOfhCUjljCtGDOfAbqvszQDwJuBGW
ePTTkojhwVJNQ8uqNVnWtq6TN94CaTzTOBToT07Rrs3+eZ4q9Q4XrI/sIz2kkELQU4PaK/yt+ImT
fup+EfhlE2ckLw2JfZ6vPj6Jd2PJdO+zRzuPAWAebO4t4bEO2Wn4otMQJ6Bq3kAzfuAa/MdJS1mP
yS+gdJ/xSg7GErSOgXwAhTENiNInJBcdcDetthYm28r760agMLhUlRvQRbEeE7bKVToxol2Gmx8Q
YCc75dF5qjVwDAlD30U/WLhO2r2rW1cnjdi2mktEyAmcXenWNsUwoDmkodvv/z20nunmbDTU8/nU
d/YD9MvKN2JxrS7kylKJ8CgQTJOi+HntdPMV1TFEeSkFNUFuLkPTVQ+d0P1uNQrGK+zJsBs3ibg5
91C86+0j8AVsNBNA6Ce9iU2MeHxM1e9KjXbhLvMhfE6gBLG3JameFVx+ROjjimeAh67FRAIgRnLx
SbqdM/CxpqKA3vw0FicWGsyyQyo/8g2a9/BLhZdpzk+klgHUtteKtHt/WelpPQutA5QwMYcHqiJp
iSB1RtMtXTYY9Db6QyOBIvQw3G85Hm7e9bDJuEI+Tk4tvEwebGOsTYaHomTq9DadB1c+d/4lwgyF
8r8jogxn7YHRcP17/+aZTziYm6iuJwmAXkKrnZDQaydXzHXN6QPxUG6O6+veMnWCC0Xa3C+eKOyg
O6vg4CjgqTGfo1l4p0aDGoM08aGF0KKBOJxA0CF9K7PMeg0MoJB7kcZHanX4HSe/HJlKcA6bTA3d
GYLnh4gmJYgQluHP97KT/1PeBK8r4jOtzK3pUyXcgvgrjpjaEoopevZWbn/G7zXo41OI2skGPljo
aI5Db1S8jUUkKQE0sCZkOpDD8+C/H4MNNb/NEIIEIsA4HFY4WxMb3zF4r+E1HZWfqBjRvwD72cdi
cvSB4SV3KvEKK+ddcNG3RCNuburpd82zybyG+jfjnhuVtOSPAdKQ16tV4DR9KhLPQ2Ut2gNOfUn4
dyRNljILbmLgp/1xwN4HkYCfW4Fd11fTB7yUrkH67ohRMVnMNucqmVK3otXkx0E0V8skneRxg71y
wS1fryQMlcqFRzhwQKuBwusQW+dDnXMUkP+BytY3mJo62dIUJfzJPr0Y3qm3Xk8ITaI6gOZ4aWUf
jop15vIzmWsy/NN9ZEBw7kGp/5tAZxcgYpr70RBB2vYx60OFCdmPPOPTvFiGnnWHCD+5LcTfElET
oCxVzZvx9/i8XCfjvUyH9aehrBcRYnq+FQdMyabn2uF/jvafei7bEpKuvyW0YNllIMJ8sUYRuwS4
Y7uIaTTguGWmsyF1KABPMHG8aHGhwHuNbEGHi17+I5Vgx8zWDsAronQHrNM/DwtrHIeeNjr2RBX+
fMM0kbt77JLjlUM6ZkjC8OYqcGYuiAzsOMJKugBGE8VAbBnxb9qcwy2cXvR4sp/sfmxPuco9XsYF
7XfBW3iB24a/Ca3NXj0frNX2JEDsdX97eDlkJ06+DKg1O/NEYiFOfcDs6yOs0jDw2B159AFd2fth
qy8ivp9PsJl790/X0yDkufOnfriZdO7SCPh8K7Nnkdj9cz/6oEoA1nekRfkJGBVcBP5/mkhFYQtz
FdgnnzhqqbwQPFObpk3+1yk5xb8MvjlYVRcERyhrMztnTTuKHactOXVzv2OeizHrsFkjgqeQxkDQ
2d/SJTIzMGo9sSrP0OSMo90iZligPDEDMdr94A+oztEvV1aFoKLTcgK3KDiHG47ecydULsWGWfz0
0ztbr+aNp/XxojViM2d/d79CVULgLIR6tiTwH2Om2CDEhCfrgRZGjYwzH1CvL3mOaHKHxSgEjm1O
NDIr3dJNVA3MBS5YPeD7W+h9HhOCFnBVIL5v05nYTDeyycjeyvXwTeHFWozwwQEAG7PHXUkFp8YG
AwakZcdM2d26TPl0rmDKMsYv2L07487V4eEUZc0r6IGQw3kNv2rF7i4/6fuq+3K3WCB4/9LhQysn
83TXBiWQ2OOkFlitCcDSv3wPNzHeT/C0slQaAfWPCUJQXWx70IlN1tr8NKhjvfjeCjXO+Tt58VGC
K3yQtFwL375Mdcxn1Jo117eLEVYVkbPkZ63eRm1UFffBN/LiySursmkPXipWszmhhaahbqJZlltv
8MKBpuJJ65ufpxPJXV1sM41ASjCFkr2mvr0LpQbxwWT7PazF0Rzc+USirF3RUK6wZyckvxHLOpDh
t4SE01mttxZgz7e56NnP4YPsA+7McVNtetuaIa0sqezu4yHnJBudQpaXCHITa8l2u4gho04eYmmE
fZ12KIr9Fdc4XGx1Ug5LEBH+9FIpW3grcS0nXdlK8zP3P4MCSR0j7sOnP8/iwzH0I4372qt8jaEW
izkxbeAkhIrKwOr1Im1QE+DugUFga5G29t+8m0aw1GsgVDYYKmSSKFMw9TkNDWsVVTg0Tfp2I6m1
t3up+0uuxFKQ21tWMY9d0a/Ix5Wg3gqHKRIq73mY/jT5K03RDRz1e5+j0YsabH6Toeu0kWU3HUDP
aGJjgvUkqK3ikxIDU8GXQtWbuVmr4SiPHGYuiiRi7sWjFy74QGwsMouckWomS/7nXzm4qp+SPjOl
kSz8sKMEuMM5YjbnBZnMLjQB+WsHZAt7EMaUWtKU8G1/DlMK2no9hROaTFoIC+OKyVFyR0YUhetH
NbtHzP7BNd3Q4CE93ttEd2ghvXFTls6UVczH2iPmkwjnSpZRyUYz2PJFmV1WNtF17uC9Ic1fUjki
BlvGMOX8AcwgUtfv/bkeuwr88eVLkQAypYu6RagdJMBKOaBaL46etWF69hLGAxNzd/HBK3eiBDlq
KNbX6T4eY6gYH8tYIY58fNtHKNuLJlbif8kqAIKLAr4NGzZfuY+o4NrS8xeo8DXCy+kyVUhB/9vU
JGt1f5TRmUqNZ4XwfUZ2ZaXyNVU23ia0AOh0WiFt+zD+v77vkMk81vJEWCR6zoH5IJiywpxR/Eb6
3zi9weSrznr07lLPYwUDVCE6ZSjW/nrGTfwJZRPofHft70/FB8r+XuojR4Dyua8+rHJs2rPIgbSF
8IdI2zuZI718vg5/9IO+mmByV/+l8GJoxSJBfKug5Xb0RAnxQhO8oIINgUkk64K4dcKRP9tSCv+N
zixmN8h2tN8gwhvjqgGdBRjlgp/OJQi736UzLbaGhJNe4kl5w9otXPxj9ks0KJvfWvsJf8n9/oQk
7N2i0kzeJBS1zaY9RpOuMkZXwnD9CIl4rhMtJnYXlBP5+DTOY+X6szVqrXpBbXoZYquqakim5Jtj
rm0BRQaLN8pl3QdsQFpqILpOKdYvewwya+yTpPtoHJ3BIUxSmpOI0PJBkhwDWUr5lio+XH8rFRUo
PI8H/ukjd6xHZDCfg8iZ9lnmu32WzSb8EKcOmjwKJSp7VHfqSvaTqJypATiqm5GzA8CX02XhK5mD
onIU5cg9Bxz9iSsEZc6a2LjyoOlyy5TENHvbd3WVsEQ4Il02186YFpcJtZFYryk2IlW2j7Cadh7K
g5wjn5x7xdugt3RaxhwNkqtzSwkX7/KomMG+yYz/2XIwZU14B1EOzbrLwGQ/oJE8LVRBmj0d3AoT
pwNjwZeYRnEBzagNjIN1kPDw4Qclij/bLVmLZDgI66C9rvrOgrQX9wDGGAAwxgTavkZvB4mFuIso
VuwyxUl8W0hwEbnqArrFQVSuTwyGDvwWd1WnkG/GcAYvpJ0jR05j9mqFTucl0xOxsL9tKJ4Ue+Ci
L7RmZUB+gZfw+gKcM1a+XaAcjXw8JcToyPGDmOpm7rzWHEeDi8ytsRU+DyM8BdD63LNHbBb8Hrzn
1N3kd23+yQRfn+Orj6hEAyXHGsMG1beu+0rn/MEsFiG1Devo8RkVSiAv8OMvW7eLLLvnbJS9NZx8
tubZwEuJwJyQpsR7O62qtQI2mcEWPQq1WzgHoW6fHPdqhwh7zu6CMfL/HnwAaAuWrsy/CZEqAbV0
1yDCgHP2vLjzKSXsgv7+Nyo5ngsC32hk3s29EnkwF5rNDyi4xUEhPB353TDk6l14KZbs3D7S+Lnn
KmSa471OwXylPWhp05zcR//KUU87ezhMHmBeyjpQyPAhcVVg9FFoWHk6hZmSwl2Q2xIK560l7Zie
r8+FYnWtDyN8mhFxw3ruVPoq9X4iVSR3SBE2Wlx1hv+8DA8NYqQxPJtulXQvjHw70R0IO95p/+Gi
Q1R+ygc8idjWt1mR9UEpdUtM6EABSzEiqnCkUr3OqrzNAvHmdpZNpSYnjyLvad+OMS6Q35JtCcGm
PFvpYKQSRDXG23a0wf1jaCznrNbog7hU9gYAH/xMepV7455on40Mll23uwybvyDhvV3M9tXJtBRV
/zU4relbhsO76cc/cQBjs/8z+q3EIw3BGdG7g53qh842w3TN2PI5NJm+bYyzMYPvwbViunAkVsuK
h5RddwaGkwizu0nOLg58JMkeS+kwGWCk9CjShnD8+Tpwp5HZI2eAmRAvQ+GsjP/PAqRwog7233Nf
xJPQzlxW9u5Wg7iC3G282z4Rg+msTYdPCTazN9UcjXFztnPWVXlQA71HG3fm0nszgfrSlTM5WZqe
tRmB3YN5+yU+QNI5l6O+AhPT8lEp4hvAU4biu0ZwE52oMlpQ+krJ16P9IsNB/zxy3f9jsn0TB9DX
wzKcv+XDlLTSX+xUTyUiMJobsRvfpbC7LfqlmV9GNUKXJaTduxZwi883KylXuNkmKXmUlDIlQZy1
vb8kA7VVH5njO4QS1n6filD3n+mRG6VRtjmK3rJf7EMNTd4rqrttdq3wzjnnmuc/9t7UqvpIvSY6
G5mLCA6QzT8WY7Txvb8yJAtJDwzU5ZA7Ucwp3UtwsYkbcD/u5eIGtsYQ6g4BpYNPq3fbopxhDvF3
Xu47h7XtO/a7BQzuF4N/TVZLyUfwAJPFIJvMiCPp44irQnpA4GCX+KowzUZxRXJSXbV16dZxI4vT
45i6r7vthqVEaHcuIYHWO/GeI6oC+W15Bzoi7VnaxMc8tQ03yPULuttGT5v8FE1pBfElhHOWleQJ
4EfovI8A4Afkk8XTxohBeNZmcD6JUTOydtXjdxQvj6hwPM7liMWiyWOXir7zYRStlAsVXvbb9njP
LkAKJYj5/wNKm02c6H0Y+W4QP52BG92fFcr7VCGXOFuVjupMwGHksn8XfzeeD/nj5XOCWXWujso4
1swYsDSRFePGt/CWPC4hPR+QcfCCwZQPuvY7p38x1c71+HVZ09xoRFzeY5mjbz4M8W3OPQg2K+/4
C/SHu0IiVjEpKrxIyVAdZcv2nBLLKuhf0sXgI7V8Qk1ipmRHHn5qIXgf1PM9jWviFLfyGhEtJiPu
ZjcJL77yW57CBOSNY+QKAjcIhS8FaVL5maiFoV0JpSoImLwcfIRkE8NlRWDeFnd4G5y/HVC7X/ks
d2rHuDpy+AovRqHzcSq/1Fa3VyIbesFHaEOGdppnykCq2PJYFvtZWsLY/YmK3G7cZPiY+0xrYqQR
2+ltPUvxn6F6i8XWKOgwTFYVWccO9kWvqNom9PVqVPnb67cgGjzz6a8f6BlSOXcCJjoVll5o/6pp
EEmLgue/Sm9aBcFzDJImidbFKFJAOky7LGe0SQo2obYdCGnImbsgPR2lm4sbqQ6kRPLWm3vq3/4a
J9IO1HO5G+E5AjVoKnvVzBTmnh/8sI/iIT6ygUI4NvPLwTDNoXpahbcueZCGoteECTKGPb4DG7Hk
R5/6HX388NMkZGi+7UB4XeHCi/QZy6K1eyqBblT2rTlYwSo35c3wLJEK/A8gEmPSrUO/PTw3Vhn0
mtfuKPglC483kImrNAnhdBOHgYRbnyzZ2d/102GHTlzJW5D/lpCV5TCmW7ZMXxJsOF37B81M82Zl
+OuLHZ1SyBCU7hsDN1oiCjzn50c08i2fm8l4zJtlBmr6FmIEP3e/FiYLYCPJJFcoG+2JMh7zXAUz
uCZaUjr5pVC/M/tALzgZnG+qPkepfkQiteJTwOJ3tIcijPA9Xp+AVQHHrvf/Mx/PRcYYpGjvlKwk
5DnhAcOufd1liYj/K0qzD1lEkAcADNTTXhsfTyu1Y79BYi0Wo8y5eibBChk91vUxZgyHIBQnITOq
3BJ2FnM2bMRosuT3G3AsPKKDtcWKjoRWOa3V4YIlcS8ybxOJyAS5DAs5mwJEddvV06/kpuYOHzrx
4/3+MV9n6vvKAnYJevKzjWyb3rYKAR5l1WUJla7jM5wumjqT3fAZGuQmzik0qQoPSR3TDvf5oWBo
VG3m18Jah0/pqarTVMEib3R1mRIakbbVU/UihMqeR3Jv37j8qnVSDm6E6HDWBbsxZ6gCT4ZH7D1v
puYp9/TyUUCts0ptQBwyuWkyPXi/w2RUdowgBafzxnnSKlPxRE1mEeXeSAHgHp0UA3b9cOolhDI1
qcyL3/MV6nH279trss8btpWCLx8gwe87nPAm2KnBxejHQHStfdgMobrPw3v1BkPhF2ijTorIMqEl
eo3eoLRUPSIcE6R+B5sseXHiGl6T+0QxVHmhnZfwm/X5OzeXkmrHZRCOr9cyvDaiTcqZl+Wj8XWJ
DAoF708kC7R2844A5Rx2zVgEHs3Ma3flEoyY8qLRn7TK+q/jNFTpm44Kc5HQyEGFUGjfGtOZsbUx
nj7p0GUCYGo+HtyeJTbx9Ql6gp2j0MGaJhZlNM0V4PaJOxzkp4/DlnJWjlj4RdEAji50nL7f6Crh
2O75T2MJfqR2fDNpYG0Wzsqo4LRqTyC5wNTGcJL+1BlsJ+pZu05YjeZbzHvEEUAqDBmfDwO/8WZR
5efZOOPspmOkHHGCabHOn+bRgBDltjVtGxsIcQzghqOn6je/9YClPlxeDrdJiFLMD4//3QvsaZ+h
X50vi7B+NE2XXpZLDUtFKYHYRmu55H+jDKQWsQDCbuWTwNOfm+UM8NVx7mcDBQVIvJL9AFua5p0E
zXpe8Ce28bsUVZiRhqlUi61rRe113c9/BtHOhMnnbcJORKlsgh4jVo5rKdfDxb2TpuqoRgQvn6K5
ECjOQvMf1EVOMfhdjgWyxJKwnqDdblBDh/y/2ZuuYtOqqOTeXYKZqOZms+cn821qCehzAxmjxJbl
jMf/fTpm5/YDRtbYS1b8a3Trm9NCzvj4awaE/b2IwSQlcWO2qdSwjGALKdrzV2Q6XAymHEYhHNGL
X+dB0WoASPboPST+GPB+PsGztMIMLcrz3h6AUXMo3x3HC6MV8f6+WTXzmZiCf3zo7O9VyGWvhEk9
MVECz2gSZkEBdLn5eEbbErNWjMyIJjBYZ9w64GSVhagaMs8bwGEiNqKY44KvElx/aREdq5gM3mG3
2iwNz5UIeNOvQgt9PNnW4ygl/Yw+j3UNFxmkHe8F0JFooIuUbbswCbNI89J64JiJg4e/+D6E1rOw
WW5JbugEN1VXFUj6KsUBDX4SDYIVahXidtXWoZxrCP63gLi678a+5KSuvQU4PnxH6qwoCB4oB8bx
JtL+OeudBsmnO1neDX4W/CqilAQV6WE5qT3CHDbobHN20b4ibZJI2SmWJPao5JWic+UP7Ht8kN2X
D5XtAFbKItFJlOR44c2zle9uNwuWmZDdtyOXF+rgbf4Vm4Q5CvuxDODAttpKZD9Uowcu3n4FX/WF
0QZog/x+7dStY8xOOjgkmC68iCX65gOWMbWrYzTbFNs0e7TvpSeYb6CRo3qa/IKVDt1Wnpc86FY2
nl9oAogsdO6KVk+jSTa3UswaBJXNq2FoBUtCTRfzPy55z4d+Zmvb9sN4qWJmqdDF4VDggm6n0gc8
RoVSYgDOzUKNznjH1/xuqtnWOXYn4oxwV12Pc0bJX3ngto45d9jQm81wtXlUx27jQfOLAeqyG3Wj
qvZAwZr4tY9uhO/xA8OfP+ZMar+Qwp2QvxN3qYAmfgBT5QEiHD5uoCPIp+Bz3VkdgB3g+rW3m+6F
C7gxS97ymamzGFMvTVOiovKGH/+kRwaOwdY79djPkMTWsCXlN8s2jVbx8/++Wxs/jLhfBeBmBZ5f
MAaSQyqww5KV+nhOPVHHGvbzTfspTP6OnZXsiWjZqh8NwID0ah7P5zSxC4EFYMZxxr2qOBY3poK3
PbAhmfYp9aCYUZFhTkHVPMkBMG28TVd4ZuQGxR4s9/R/GXENQ43nRPxYn7ZdjeBdP0eLgldeBOdk
K7o3z3jBMsa7brklaXSHkksOECn05+/QWav6Fd6GeY5XxnU2Y2sUW6TmN9d9Wq2HVLyKpQRauiyP
FzHDYq07ubvPZ4BsUCMypPWfTr33a03gH7/ATElFLrEuf0QrVLzjNuCDG8GWd82R7ibuXgSnqj9x
mRfysYVFNQi4J+2w6J3KXnQz5SKUtFyvECHx35tZ761gLdJhZsyWcPDB4tTVM8yzpROmnMTEhvUY
Jul8CNoqkFa5dLJP8HlZKsii2gaL+ip11xA0NRPlXjLBRTB77pS1Di3g7O3/iMsMF5u9/uGJmST0
Lt4kcJhXOWKgECPid0yQOL/povShqUFlFXsGIC8YHjuxbf4536wnccWMTq1xe5LCjZDLQMBqZKE/
O8ItEYVJrpbE2ohptRpRmbeOlRg2tY9a+EG5nSgiMm9zjiwejiGlaetwQ532Yz95ryHu4VbZtSyq
1OB+GbslcU4rIVr71/kxtV/IYlxmRUS+DtUlOVl0tKf2tprI23tGQOZs4XLOTy54Qv0rgNS5ANGn
HZkcWX2k7bJ/T94YUrGb2mtIi9uqFBHwKySFcb6TRQLylRju/kR9e04U0Kzib0hQSR9PWFZS5ssV
shsw9UHGjXXhQD65lOK8EgpxVMo2rM99V5mI6p6EBwfqL/ptW6oHBX4RkcgstbodJIGW9hcm8+Ja
rA7CSZCBWNSfBAMXssRX+xA38CMQlJaElRcEjdTSlkRDLKxMCWMoLfzQCdi4T7LUnQRQ6Z+w9fI7
Xe0DWlYDzqGjseQt9/BCNZV59rV16u2YIqhGJK15Lp8zJdKXnNP1ZflaHM0Pax3Lu80z05HU9gFP
NQloRn7eiKKmr741tfYy10G1p8Hmfi+CBgvEFSRkcVhbPIZFHx7/auMYTCrm8VHiX5uYwF/D04to
hoaVz3ahe5CaGSWmXSOTKl04gr+br+zqUXxpkBvV+9wt2Wch8E5mD7vZQfJX36mEWFrvUEiFxTCh
xMT6hUZIdkCATG2RZdE8fecD8xwFIBSkku1L7uQdegAnpAIYUaJ3IcJppj1LgSV+B7FZ/v4XwDm5
UkezsUvfPLUwGfLBCQlpw/BduGh4YyDeTX3jemLFcNMRDVHPAQTIHAdk8zuBM4qYKNlE5VVKFW3s
W2sbFE8QBvAtlLXrJvLXNtonPwffNjBRntiZMTzR52zbKvxMG2AjlCTBiV85zF8Ipi1f1Lij3cwZ
Mv773eAnFdUqCZ1nCZSqOwPwD3n9ucoMUZHDitcPscIJivg/mo/eMLw1/6cC83XuUB5WytEVtPet
oIitNsqfhpTRu0c9YyXJyYFWfLZ/fVOjzzxsB9JlG68pRgrOV815Ypvje8PcRjo/qDpFxmMapWU1
mFR7nrVBEDF0vFKjX5O/61RWWYuOUE+dwW6pdkyr2XVn/RR8aHBfaJocB66v8HmCzU8ugz8Tv+3q
xt4ZKC2jzCFomeE5CjPAMyTnRVVaM/vJqLDNGVF5wMK93qjvXYxFwZ8GbXeIBVu7xuVa/Jc8AYMj
v//rbOLqdH+NvglkgfJNMQaPNRmxKn0bXhFA2TN+8vE76R8k9YxP0AJDGQZcolPJXG/Aiar3bdZ/
0Q/Iy4UkefVDgSsA8tC6XLNjzO45w/UxOVTuF9X3K5GlYyB0/3sSUKSLL+bGu/X7KLR31ZRv1h09
94p+yZDjF1kAXKMy2QkxgWrwgx7H4fEuetPHEq3qEA0TewRemNsATeT9P4Tcm4O9kwgbnWBCsvzA
WWU+PejpGzio40NhphtY1mzeh1gdqz8T2+fnBkDdPxwkYseCqp+Bqs2jW2+ZFfO3C7roQiRp4jji
YVD0BnEeZ7sOPNRTmwQsPD87cSV2xwxFswG7BC9p1IvjlkhwLaZzRDuDBUoxCWdMEvCMz92/zAox
LJc96ZK1iFMWaRsu2j7JHS2+3pdvDOTUFLU8EdaUUW4xyKsdPcUiLYbBo0nUGLOL6h9Mv1r2KVEJ
i2IiI4B3V8HPmUB4mPmSYSV6bF56Aa5cM15xSU1RVPkfE7pSTr4dBgoIQoCoOyQyp1X3w038axvG
oiexFW1/H4nzHggMgjg6jgdf3s+KXDOr6aN+zvu9pSLazyjBmHQ2Tya1nI8ypxsUl6MKZnAi/uuh
v/FhEI6wibca+O6KrAbx4tDRPqdOG52uCxi9QDqkSOMW9my/rHMAHkQSemDjAHdEeQlgEhcOuwUi
isClito43BIwKuAUnWxQrYSLOW4bDk+r/j/0S4l36yc6/GDgYZXVR4WKLzXNO7SAYY9doLytk/v8
AX6ttUAcVVjEqDr73m83Nj/T0bQ+KDb3uc472HnfS3sx3J49Oq/reZhNAl+fwAxG6F+abAOidGN2
h/HkgYh5fqtQIU+zJtvF91CBXBUj5jh/hQqKKAjjeWuX0kWztwkNTAnXkZiHTmMnL3DglkASUj3n
bA9IsIY2xqvGXNyZGnTjnLjPkwYhzibGLXB4BLK9B2LWshJX9baMjMlHoQIT35WMpxtdvrL5ZU0W
swet2o/bEmZrMOeDH3XgGSLQec47E7UyoqJmFwfdmNcHMgpFVwMidv7cIa+BVjxYYvbdqgp7bgaS
F+bKMj2RTztJ2a4ok4j3Vor2Ervb3Yy4jjUfkd7h+mkkPIohdqzveGCq5YdAfVOLjtQ85+USHBZy
6ZXo1zWD2m6uV/HaK5s5TdQo5SEfA9i99P5PPrElUTEEzzkN1sx18YIbY9E45ZEs7ZylAdHRmtSG
cLLy4OlKO1gmK9FF9G6PYbOjvkqAIfKmNnnAucM0tR2VL1tD+D8wTLvcdLHAoGPMlM879Pesc8Rg
99Yqk3LffrVxJ1OijHm0PshkIeruPpVjOe8pu011A7vY7aFUZLO3UahlsKQLRMEH8IP7c3Vc5pql
f/BjbM4loM2gm2cuJq8KNe3XtB8J4Uobl+Yml3Ar0rQ7Oq0NQIhuxYdaAzVtzplQ4uOpEsMgj0/S
Wevbewg+0iuiyi1RVLNKxVx2pfTzIm7Xzgr0i1VyXevTd59enwr2VnNVqFJpYjr2bnVZJ4gDxjXr
KEnzWyduuGawPZM7eeE1DkdgGu/8SNTHgfFUyqbDZPGT7dvLeBSvB2O7WrMW1IruJVvWSubaJvzf
nCVUzB9qXP6Sjz8R0e6ZCU2IyUFEH07r2LPnmDCBOQfwDoxKEzStHzR9D+ZjJIHm0tC+YvS2YjOA
MLWCsRdxsFFoG/8EmQuxOeWpiodt2oB/fAgT2WZgNdkCUAWOUlg/B2K6byefK4s0p+bh131qhUo1
fYe+dllzilx9lKDg3AfVwStZa/me9U8kXG1fPNFq53dkXXtLn/k/xox8+XZehQZNjvd9TNHMnnEv
aKJyy9BmJluV0oSdwXqEbf8x9iHKc/j+VQkmf/dpzzpyVLQZaEinIT+6Zdcch3KrmNIYgXKZuxAr
WM6o7+W3aOC4wtOW0BgatZWWK0EGkFBXijVbV43QutXNyJj9m3i06+k2GF1RL1nMT5OHmdXCtnlz
k/S4XMlkzymZVbBYe96KG4U9IQtMH1W8eCmv2chowC6+fNa4AJNDZ8N0kIHWj3kkTdttZaTBvcC4
kPPgFuK3rZHTglYZhSGe/QF1e/sDfD+1/dd5PdMmiXay09+3AJQ4ulU3OaE2lMl/VVsIuykAiMDC
dwvEbSiuB8TkXbST/ZpByuA2SX3WpCfCKcDBpgL0phxhUunNpNIt2TU4YzD8KT59vznYYz1XYqwH
SqupTUwhbENZDXTXi2UIOmI+qjpig0zJHTkw9lRUNr9fpBDnhwn1yvaxm8x8wKkkF9nXeQHLC84t
t8Prsip2QVQyygKmr05moHf5EZVl0TI5CqYTlvulkMiI/guzKJ9LyuSC5JXIhM/oUpUt66iniaCH
x9dkJdbaIfKibYgfWtKjhORVW4GP2ZB/PR7iJfDIP3dVsOIXXIrIpT2Y9nq51bCVXzQSTNu4U2vq
r3uS+vGjzI7BXtz6rVR0KbgksN0L3gJp2zCVQs7yyItYdUaZ7nUU561OTcn18ISXvFsQSrPIWNZL
31aleOz/ZXZm0CFQiyW+WKtRxb0vHQhk42i3jdurHZyFnK+q+hHgaV8N+oZdMj/g1FASbXb5rDNm
10mSgAZfbZXT6eaTYA+36Pnz92KZCiEFCZbsqBEcYQh49aHSkvfPnoF05l41jMLMzPGDgLgTNyrg
S2Wr4TF0pWMio7v78n3lBeqOj0wp9iKOCzdniqE2MyP4Ziv7bjVTvdJ1jyfqE/MwkzBPkxn14sfe
bHjHQkmNmIk4ZZY+KJx4X9enbrdTcYyonn2909CWusl7zg7b+IgMhqsf3UnMtWOCbUWz1eJpY0dA
x3TaMlZPAJrHZ4gexSEC/CYLQoc2FcZctw6vdprCLHnTKLmjq13DO2wIUf6SfRzEInVb7+glLZY0
Ikzdrc+j7Kj/20XlD2w00CV8Dhgi9ohzomCzPgAHmhs+EZ9SrJ9oOBXCHuRNY4P+d0DkxyxkLEw1
sjJQ0F3FpM25EEUpuSYcnQZ1x1mfc/7rISbkYdiU+vMgywD7Nxae4sQj3Z7Nb+x6Z0XD0gtC107p
+gC2djVhULKJYTDM/+hiobb2H2LhKKz5QnMNHGLGTadlFGunTWJJgzb8hCAK9kQoV5m5pOJPoNv9
VfDOI5IJyv6kpvIXelE4LkCID0YD2nXV93JHl9nIZBfhqH0Iqc7npS8kWnXrISrSfRGECKYPM7fH
utV4NFpNL2LWBDDmXeoGit9bK0gop52D9ZqaVVaLmJX2ZRhyjVyiRN2GVgZ6Flvn/4LW95UuK2+C
ZHfxvFupWzSINSYW4RvFAs9P2j4p2nqlief11VaPZp5p3h+yXf1iu4kmu2xlygrEN/PRRZnxei5q
xc/rpiAu5rqmYn5fX+WcQvmDtWvhYLzX2vrtw/8WPHjoXPB8KBSz/Sp9wWy+VXkGCkp+Up/EUJI8
Q8mWrWHXGHyil4hF1TkcyLEtEVE5UfBoFnEfMWO8v//A0XxfeUUc7TXL4WCQBgMq6WDr3FibNSub
ErbryTRtZX+bUz/dodAkQf/3K3Pbq+8/MpcEcq0qDBYSKYw6E3S3pzDMFH1eUhqHFdKF/evJTeoM
LCBztVe8oZf+rzdjnIvl2iWl3hN+hPkhe5JdP1G0AO6LX5X74Fd0iT2cX9z3F3g/JSsjmmA9rcWU
AL/2I9gYdOyjsaKCQe0QhcPG2yZYjFhR248xKq1KL7ayH9pNFTp2MBxuCk43N7p8IcMUs1uWsWfK
xSl2vKZICAAPF8STUQarwMtDWAbl+aqzxGK2cqN3aIbd2n8RBexvhHDw6cO4kZsgecVllAmj3zCq
sHHc9ptKmyIzzw4ud5Zkj4Xpt5PUoEA38/EeQfStZR/Eh+LCDvI5v3CA7LOp7dLnAOl9jh9/G3YO
jtL8SgOx1+pq2wBXl5bSl2IYeSq4IAbfOUZQK2mWQnd7m/y11DCs1mCEVVCAQzxTL6rCjNQ24S2N
MuVSmYYk05VYOTBWsKSUNn7bw8yOnytq4UvSFZS6RkopdzTF469EXGU3gMl9fNlpksoM52Z1VvsK
IbybtKy3PgpgBGBdwHqQmzR5HU56nuc24jb0fKB/lQ/eKUPlrBQHcqjrMbTf3Sxou9WmvPGWIpfG
rTVG0Qs+ighX55gGy6bNKAy7OVWiYPRoTzPjDhlFBmcUpg1DBEFB0EkUzfPYPv/Hde1sgZOX3g/b
fR6AaLS/RQ90q4WIFT/CPWUgilkCpMm3cQd9Ch4y8y+1fnmcDdxkS2uxuf3/BXq7lAoZdmmGVfNK
xjzcxMthsd5A4nrvPy5mfLL9XGp9x2oPzEVzdlmjSNMRm8QjaBtXMzXQhFOfKq/o7fHki0ncef/j
cYvDxVipxbWLLjn6jXPTvCy5HuqmUTmUYIf1Oc3c/kU/S048ZYU8kGjDoL51e85c39D3Djq+cQ1c
dOgbdkI5fU8juRbDlqetPDSoxUdqjaJ52hhUcplsk9yV4whcCeZmbVLlpZatW48b3f2bNt2cQynT
Zx+Xhsrx10bgh9YD0/bkFHYchesH8vCX6fuDTVDixsvGMj8oZOkBtMIOCf8t0Enzra3QoRidvNIG
KGP8S1bi5uWbAcc7IgT2n2WqZrwoBR0ndUJPkzDDeQKrRh3sEGwWSgJrX/T8aLP+EJ7caGqyaOS8
mNbmDEjsXqY3PVyAhDwoNFg4XJ+JmdtXvS8Y2Tk2fWJaX1knx+NZCJHv+S/ICjLNvxl1JyvS67zA
wEZS/qPHrfd23PnVe5hpUmbU7a+e/jbAaItDNBXHBieTTZmQ4ots09WR86mLZCagBvrdPqvjioX0
sXUx3zJQOPLIOwvbV0SJubEjyToi84Ne4Wg3IHJgypu2/XzWCC3PjiYoPY2pUME/0FihfWLzWI7g
EH45UvQgh2Hn8i3w/Ftqn2hSaLsnjnJqRyhI43jVkiwqeFOEC7LS4U56J8vLjru63FCIpmr9OiUI
G5JS8YEovn9u2WfceKPmc1kJlBtp9pft3AVplqLfxANLapT1BIM4h43O0GaWc3YZRRz7CN/vnihA
F0KLHMr+jeQH/BScjp9Qmv8X3q53hulfOiVRzACFOtGY0yslUDhjFZtAPkt0+Qcsl4y53a69lBXK
OIu5zfpvs8QCp4zW6YQ4BeKQOg+Gf4DzKvLFkqeZuuvFqf/a9z2v8L1NUFCH18X++C/c4gUb2qnt
kbjtaoiI9bu7PQNSSTLWI8w/aEzk/YD5qI1CUU3VQgnUxP9TwUqLWSCJzVOlA4AVjs4DQqcDkznm
EJ6ljl2hDt7530D6tRu3deFfm8czBdAKQE0JvfNIXRPjIfHD4tNv0e7gg8ftmkhLD3KbsRYqa4q4
rL0oxy5M47iM4wArEoFI0qSw/bFr9jS/BNOPXkAjwASancjHUrkDW000Dec5mS/2jVIxSrZUWb4i
LSP0JC5WxvUWwaWia0UD05r60evLZj8Sv7q5AlmJfkNeQMwFTzo8DieXr6gEfiSOD/yrHc1rtFt/
lbMrCUlq/qMU1Uv5Bq4ZjCIHQguoeySNF0J9HKY0GApVA5yD9dS+G4w5RIFMHYgFMSO+o4p76g3g
hdIu08DGsWB+6QTIjnWBEAIogR9TGsIP5kRl3GYuRoDllIvDI0V+M5cmIveu6iHgKQYuGmUt187w
q3VGs6ruOaS44A+kymImzx8BAp8FpZKZbEzTdqQzh4PqJEFUskM13hBvwfvOoXImB+NOl5hQzDcd
sdEzctq4b4BqWpfJdGhE95k0bPR4LvKEENOnWCs9vl+0VVFYRjKj8u73Win2WN2xkQ5HBPxubKis
vfqRJf7XdyGMi6aIvDfZP4poeL8jJQC/kComm+2XLgXGu/KAn3BBPd6jHaZYut7liwdi/EhucpAO
8bYS9FDP8ukx688Da/zhO82Jf34d5zFM6kC/XZjsoG8u1zSfboCIKSL+lSDRsO0aj5kXoI/Mupe2
WfUB877QxG+Re5LLMHGjuYc+dvY0u/Wkr66RkgXHMIMN2db7VnF50fNA/YlbXlVYxTR8W/Box40T
lJ05Anva/upKSXCiRzJy0mKB20+0Yg4lvsyP2kVFz6VFyt7W71vaJSkVsr8EFXx3/ynhPmDPmU3U
3TXmjAKtJh88wtidc4+QwSSEbd+l6JLvnCZGny6CJTIKZwzVJW8HeA/2U1FHhdPjoJRbos+Mjv1m
lEgMdw1EjW86wJMbq2R9O3+UWn0RhJsrFuyBWRpmSeti+x8tr2dsytYfc0wtiX75kwSH3HAbzgIO
jqkx7ZkgglXhLVIsbRWAlblnUwMrYp/fztJQbKg4ih3g5anqwYjm3XOMkJcqxaz77XfMxPkOwM+A
dyhMg2/znqfmNrJLc6LBS3SbCxXCxXX1km439IuNLoY05mYRMtlOohdwiKdI745aQ5Z42ll+bIcA
8neFdGytLN6ThD9J9De+gqqi8IaiOvd1oL3M9JexeF/EwylUfFOL/Z86p0jXdG7f75hoyJW0OviC
ahbpLIs9tzLkzbHTfAgvlz3l6/EyeaKkgKwhdjhRiAp1tPh+zFZjfaaJZDi1frahd7Tj0oQv9mhl
kcPMRSpNWhjVwXCRvup03N2szaokjcLPtrK4S7DkgTRFkYi8IZ46KgEE7Cow47+CIZhSj42NHj9Z
MS8xL8aVXFQTuSdTUK87OyfIhD49N4bpsHm0aJr2FxVnE8VRmuC3HGZbcGd/BpJjRvU/oferqhdh
h82yytlQhIkEBmeFNolDp4j6W4dyJ0FyAyqsh9I+LL8ILfAubakgTAvAvNw4dalx78UwEnAmMMbU
gK24huZaGgf63UJwIyiRl4nQnT0685TgzefzlbL8yWF3iXT3+FHqsz7Czb7jKHlnPEdYbFMGt/3r
7+ankxzmYibBYrEdfJqZ8I0BijMdwbfhSzfUh/5U7TZIXet1i2kRjKPKziDZzkx10rqaTG4VAloN
mH3bGcGErkJPsIRH5s0PB5sdOgXqJDxmqohQTRTfZVj0LJJjq5hoxjeCD9BUfs2GY8zU6BSrXQPO
JSb4y4Cs0Ql8LWTv0YGNDF4KmHP17LvtvwROXzuLhH2z9WgZIfwPFDWGCC88ZCmQ4+eUQkWeyXl6
uV5AuMKOtzQUVxs2oop1IMshjDNw+sCfype0yzLk3DPzK4EBqaOmvz9QV2fGAq4RslzoQDgk6KoN
bvVQ3C+1FxoD+8UMEfOtSPEIg9CqkuzIJwiD79fX7ZUCawQs23A3AoXNOR6+M/nDH0jiN0L1O26o
pSdi1u+qQR4rIC7Hk1Ge3JgZnCIM+qryJT3b1313dmB10F6AF6j583E2MWeKXLgMzw9/Vyd2Id7X
2v+Lfr7xC8iqPzlqS2BqukkscG1vWgT2vM5ELi1wgcOSp3FG3KRFFv1Ma1wyVW4hUq9YWCZ8QzUD
yNOYQIoHKN8Oz4T7cANkiGd49lBLDfqTuxe8zQTr+og3qMzSDLaoLc9lGvg5uELuCpRLYuqjy9jL
KZ5zFNlUvCExYL+GebE3zx19S5okKGmvmOUTzg2A7D/J56zbHZf3ZJO9UuSJ7EhlzMRFbP5vpQ1J
SeL24jptave0OVtB6bujPRrZUoL4MNarGHQ5PoSzJfMBT/BDNQpVb1Wnd2gMXNOhAnnbb23IoKeZ
l6OUK0HO/K/NPCchzeobuXzbpaA4YJHrKWvNoOZk1I5kes7KC1sz+Jbsp+gPrQ7868LgbdgbqjO8
fchz6QuWGMQWFW0DEZv162/8DK1gdX0OXA4RbAdPgH+qUHPO3HJR7bYwOB0cSpTEw06lvkEIRFLt
+Y+arBxdYRgDXMGw7XEHzQjj5d0wQ7uIO0lLm3nY4NH9+EuMYIVn3D1hc07fUA9GhQymjKcYGzuU
I5/FC7PByjCKzMv0/35Ph+v0okC9kirxMaNqOWTViaTW1PSB4inuPfkKp8r0/JFRfVkFnzn3T1qE
TdvdLmTmckfjKYmQVnNJ0KuIjlfCHM9aPJqBSWt7GOBHpuaEFkbgBGvdSNCsWIJ0Bvgz78zq7PRb
0znAn+Ysxi2tVef5TM22b3SMdaVSfMEEJ7nS2jIWb8OaicfN0qVJYN8oIoXYq+47gtTA0zUgnrw6
g9132ugsMzLGDFxvcy4leAFh3KWlmBphj3jb4RJfQSw1gzfa566PiaInsN9vf7kK7LbJ82Mk6W0Q
DjJwL8JbdpVtRWA9hZTAPBkQfldQkPGobJN0GMAoEtRsd7/Zw+/GF2l0OZ9MJaTWSF3/CosNnfql
h17EoDigA4vLTMXZXEBwKx4CNgsnTuyiMcOemNRMLIwT8MB05UKTAGd5LBMFQj6oH++qJBWWf71X
5EkphPnmaj5fRFyDlSWvf5mbKU7LXHBhYagEumUdiodtmtYYAV5y55fXSF3Sa+GcAbOoKPm95dzR
Nr2uB5jNCEVzQrGK0//RYNbwCI6zwgTxVymfoeaR5Hw5KhbbrBmMVbWmznf971K21sIKwr8Qk5ge
tQM9geQ26+XmuQPL6aSiBZzq97kAb9vC1ulTlVagqPwMwPn/7GSP+YmqmEhZ4k8xQzHCb5wQn446
ybArqaJ0EIbSjOb8HrblP8j882e4H4jPrPPrF4q+Gt9Ah11vt+3j166Mwrmdf/Uuq//ZLXrDEIV7
Jnxlgadkp7xo3kS6LX84QqSkVm7R2jdBCOyNB0hVsHVHaQC1W2+Mh0km4SnQRJMMpuHZpLt+i+9a
igWevQ3qVkjBg4OY758fbtBxErlKhbnOjA+X7DwbKZfgHi4VhYmsLO1uagxieGzqEsbQGftEeFlf
HfGgmBpmW6r0IhNbHQwqypf9QgoMuSXHGkAhBFIQraIA3DUi+K7Cuv+rQMLBGL5phmLcq82chZCo
XEHmFbJ96z4/LD4PSYtSr34Y1wpJuD1vHBzXUNEXVaNRH/CKqIEQk/uMMbgQFHHRdjAhQTEcinVZ
m67AFnHJLA2udbJZBrXI8lyVc8LFFa2ACyN7vD/VnGKp8X+Hz5tjKBo4Mjog8Ztwz2qjXcDv3fMy
Ftr8xtg3fya2gENuoSxoh5kMR+lBSWdcJXQOvNRapmwUfXnRD+EOPeXC0Ps++RRJDEzr9Ey8xfsh
dqgEY8rkzYoxiALIQ2S4MD91w71gB9ysK68AFbuOHtz3wpPIEEpkBZB202mLHzlKtzM/q3ejXrRb
nkII4p17KxVY7shFAauJtMwYFe4+KK7qgQhmkhVHoujZm3aevnNr4uqhX3aBnNAdTyMNpxcPw51L
58W/pchj9te64gIH6cLsQSgl5tYuAqQVpcuCpvHBDRVVZtZByOJWCdp6Wm2wu7bcy2RULFVe1MeR
FNcu6zfyj/6u7blckn5rNwijnjtfUekoUbGT2PHAIuFiRQKSzx3X538uvnGfEwSPW82FBXea5e+X
/+g7bPPB7NIR5o0elVLl2VHnYZG5ZHgQyaguETSQXDbQ2XhpfoNk4oYvS0gox43eKfttKkeEg/lW
JLm9AkNlIv5kkdIjgTrfKg9fT3inyymcGsrmkqSRNFgDIVqbQz9RAGi9mjsxZzeT/j7lkPQd4vmB
7wgDvyC3gugNx5kKUIjA0X0VzeeFX1xoyzmQMw9Xd45CEB0OxGjv3UpDj7IM8CmED9lQpwptV7LB
X98e9s0dUt3hefDnaVuzzKTSCBSr3OuwkWFt/QA/nt4I82CJr4e01nfr8pN3FlxAPJ65bH5+1EyI
taE0VLzzZ5tosujgsouinQj2c1H7DVCwFWyzNrLIfLhZg8x3/DzT9Rwepl2MbHbHdyRyWZtgTNtC
I2xLVFSw45hd8wQg+cCGqEitrIFzqwvy3UcHKq9GVm0qUXe6QKVpq97N4VLnrpYD0fMnuvLDbNKZ
bs2yUdXgnM5gK75F8d34XNZzXqTj9PeG2OUsfhe6mqZFsRpGxIqYnKGDaJH5/MWVDe6OICrW37Hn
bZDS83c2ELSwHxvrGHXuLc6UX5TO8m301H44e2feE5v0/SOjhnnek1k7TNej9+ABvxlyXT+XgFJb
Wy5MBxbUGVnco9zk1hhWp6H7S91rq53+npmo4W0hmHcBjToSYu7uQte4oJ8RZtDapalrJFcp0/0k
K/+yl1vL5cC7D1jDPmRyLdEb608Sw50FiOiBYD8H1l8im+Jg0oJVcFvg6G0z2gB4A51dGvPKSB2+
n1fREMBjXpSNDm+FCMlDm38tGKEDXRl6HySAruRvJqtaAfiaREp6CnY5i6Br+fegFpBOc1IE0yjY
HNUF4d34UWbJcIFgyn+iTsSRQI3zz+fs875iNAZSmIA95pTCDkffmMBddNctVlP3sVrf7OwibOo2
bSiAEomkFdqOxe7RJbIBmmw2wWLv7e6Qs8rvXo6M8M+/fe74bnZtqnRtvpK+VYQSURNwRMUu6pc9
29Tlowyb9slhnLcDd4yIpLw8w176hEsBzzxVMVLlRKdZi/N36Mf2b/NswlETqb2zgdTiDWwFKCM/
lK66VfjmxjBFIK8iA7MyhaU8m5E7MALD5R8vrzMhToIxzu1jMdR/yputDNNIG61tmuuDn7V6oC6Z
rXmwSsYBs3AdxioX97dSLUieiUEYacLz25B2w0PhT5ieHuuUg/ojH+7Ub9D718mYf8c8+nMn1vyU
cTHf2T+qZf3eieG7aFWgfQOvp72l6Dvmy/kCGc92yHYGOQgbS12yOxPlw9HWzxPH6E25VqW89wxu
BvEPcJ/GJIU9AkCpDnNLQe+Z+Q6blaXt1023hZjCPG+PCfjJU769r65gmgVY7HckN75jIqN887Jv
cYPtPWiyz90za1ea0JCyyQ6kxdUcNClzY/Y5Kckc63liiPIrE1aguuHSGDmY7n+BlglWzE5yIq95
dIyXVepntyHp47VPWQXolgAWPeQUmhfz5TEzVmLQXfwGhiBKS1/dPLXBmPf2f4SRK7BBLJQJpqhU
pRyfo7uXTzK6o8tOzsscFAr8D8q+PqFAH72iHzrdODRfSJii0AQU3MnaxUYGqbGvwRcvSEtnTKYG
cF5ZnVTjroxER8aaoRdPyY68SwxquesH8HeemAuWsBu9egbZphvQTSziHBVyw2MV2TOhcbH6XAb1
jUyn/EjpERjcJaocMno3aXLUV0ZMA8FqRPRtI/ySaZJ1hNORD16baOuiNHUh1XjcdJ1pWrviTlrH
6E+NADvBeRwoR9ZagfHoefv8q6eI4ukxFu7RSmFfas6wdjk2EkCwERAtNebtRplp856CZsmWCwj+
2bb4t6Eov8okvU9obETdLeTREO332iMKWeWjPsbpSII63L/BJB9DBjtQ7MeI0YdfFnxvCaoY5GOu
FiX2FG72NPv7GqmTA26SdRBJ7laB6Fgy6wm5Wlfchy3PKqsyyYTY3yvkZiNEiT34Fy4OEjQL1YB8
Jb8DUuSJTBXkp9FtK4LzwvDiGzBPK99t8AuXFerqJsNhEv7er8dbJen4Lcp7rdT2IEqcE2aXguaY
H5TRmXlOy4WfMIGt256wOnSY/w77wV74qmktZ9gbSigMTvNocDAqPYCbb9LmQFCYSwqAu2ksX1te
n42oqsrAl/on1APzXA+Xz9g1R6wxq+hL4eIAnzMlJmd1+oP3HmvlZim3IR99sLlxU+fYpMWMSN5h
l7NRkq7YSH25GHFg4NJ712PerVG4UAZ/uAjkhZwNssuosOY1sK1LkrLJTCYml18sWbkIufokwqIp
tbeuzfLKSrl5DGJdUfdKHfpTIjQqeXE8kqzL6P7q426ZD4tPKYDba1vuPV+pYRUfE+3HnII026IN
vInTRgQJGvukML5njEAet5SC1+viqI3+VJHju2bb3sNqRdW/PKyCkb2x4SSzfuSazSesE4yy7De/
yoFOzEvXV4uZFblbhV0AQM8/mMXcP/ReSY8IobTmSRk0xYzkF0rBN3DHmheGqSoJQTXohoxogm8H
7E74/3HKE6daJAIGOzBr08OoN4wWFIwHs4uU32ogJhJgozWwgkIjp3ok2RlxDj5hDTpe23JytK99
ssNIxs1Mnw/PCHVfc8j2MViGxFyX2JajosJZvADKWes02cgwmCbZa3dMP9HFDwflB4FF2vuYtdo7
AZzrzEFZkIlmlj1Oy4LHKrqc64SWOpU2yYamt3meTQj6DcTmKeNP4fbHruDWZPhgVZ3mgTXv5TMX
lJB4Qr+MYRC0+Xsn4FOtbvi2Wm/ErZA3m+NljdPwEUfXZIghsf9JhiKpKl8YkVxz8MoGNhK9ZIzu
Jp/L9t6m9A0CFzw7yifCi1QVjg0dUHvrJ2KWmXmDHdZoo9uPABIM54vi/1hICf5mxCtGDzLaLt2g
JjYQnImC5gwKL4ZG+U3cxxMhafuccBjBdzxVO5yV900DnKsSnLLpnY4GnpjAzZvGTcoPoV4U+r9g
7gAsViEI46Gyy0gZJCY4pTwgSApE+hsJElpJrUdpv6QkEjg7nxH7pIKhbPGRlltNpZu3U9grjzhl
fWBz5F4xJT72HRQ+tLomfT9XllqKVrD1rt/hMTf4olDW9zh7eDo8RmIMJkmOF/9U7Ot09hBXnwe7
U4G66bUIggvNzIIx+aFThy2hfYns9EPRdi4zKo3ZGZd9sIsWR2pIBwl9e2/xGJGOjajorXscnS9Q
67jqF7/QJD3G1iXJx1DY8lGRxPuAwrbO/CPZD01+YnE0NNLdD5s1Sc/3KEqswVuM47ai/+rF9rsY
hxaByaZzm46u4Mj8zS6k7RmLEM59id9BZRehTkh9ORBzThOVB1lz6ienKxb+0jDbWmQ7UHmBrBDr
4KWbxA+BAIx8xtWsysDhUrwUij9Y7s+OsML4R+w/7QnacKvm6BvW69fQ0mYAdSvLOUuMo1B4cgNy
rPkMbkfFvmyFK1sNh0JnSbeR0p/l33vbhOtwoHDNMUZOxiPo21fLKbx349NTj9fUdmRTm7SkCYF9
9B/dzILQJUYyrQr+A8iiycd9tV9wtGUtishUkRGZid87j7P0pMN/Ob2ez0tCXCOz56SSffUu23pa
p7LV5tEsbhPrhKTucJa8sfLfHByucfou4AzdNokd5CDvhCGMeBvxc70isa/Rl5RQzLuBCRU7rR3b
kBmka+U3NyFw08b0gpUGfFXXrJHy4FQ4ssIsEFXd3yj7o4Cv7ItXRyxCpSepdt6x18aZvQyqTSm5
v2ocnLAwH+IaJRC5/pyjDKAT2Pzk6gpnMJPE5nj04k13r5qkub+8Kisb8+aEFlpdoDS4cyM1bZ76
ZMfAx9Xc/KmuOWusOmxU9Qn8flVjuV/xwFE7xZkrVERD5EjUrDVbrQaiV9YBhfOHDc84ox+FijPH
x4439iAS3THuc2cJGziARTzpo2UYsWuHZVEvsNSXM44MMweVqQlg7qdfncJURFaFSfhavuGg57pP
MQ6c3C4T5TwMux2IRQZuzWhZXW7CCVZV+ZkGRxKmg4+VziV7aksW1TBWx0r17nzWDxt0jUwW3GCg
cFKQjtgFFc7Ywa842/nzU3N0Y8n5MuAulbBaMNHIkm1RzYfaKgPSTmjISGQVtoQuAsAI0NlSB8cW
epZNv6r2AW3Cfv30rl2CRGIEJhkuUaYgy10ZzKAE76q/enEHKQdhmTkHiTF81N31Oxsdd44riPtq
aThCOb2tk/Ycw5lMp9jay5i1ON0LatUiCG9WQzQ4/vPwKTtTfjVlH18p3yx99hQqvEwvd1JITTCb
KDjNQIbOsgtjqLR00ROVau7avWWHibM1aeepfKmEbjI9XDLs3fUK9OgXx1bpVN4xqZAkTNVhX12p
p2i6a4wjLnwQkdwq0h/IFFWVG5OyWImP/Xq8lIKtj8qQauW7w2Lkq24ojsqmEVP4Gt/tJYtQyjud
46BujpqUe/hvkdDALmYoI+DDqk9fVfhqlilEXIqRNl+UGgI/x51aAGRMVs61mwb0dX/M/FffDhiY
m4mCNsem5y8NydW3NExzYfOk1nxqn5rLdZmHrxGLtPCMbHe/Cny15Bic49tr9WCO+Xp2uLGjK7ag
hTHRDghr+1Oabjf8Gfp4FhimqF/sTcDCyvN4L8/hDRghEabwWQoww8objCI9Ye/ivKTuEzfsax0J
d5j+HUJq0/Q5sr+M5O/857llQkztiQAVmnPAK+9cnKmOTAIWmdOoej0BixB36vBsM6sail9Yy980
8UMLYdGFbBnZAWRKzW7z15Qpx7NbtCwZ3KoKrQCiRgHshe6oh0ISsV0hKCmEKuV/cyGtIfLZ05x4
Kld/3YVPVfWH0xpBMBTYHJNHIoBWeVM0qqKps+fcvinokGLhYU6feU/xXWjN3UXBrcwTlbLGWYNs
IVL5zQf+iIeLCnmssHKPrSBdu0m8DWTv4dj62KX18mOaL+MlEgTyrdjn/4FGa2t9uC2nMRSjE5f6
SAz8bVwgGJvNaksU674kFTzM2cgZt1gegdJzvZLNR5oGXYRbew2uWeS/9qwUSwY7Pbz2pO3SkJN1
ktHv6fkb+Y1T7VOQsdIFmGg7R6nkVj4v8WAxbIpUM312/tfcSdoeML21AzvYdRv5OqdnB6hMvK13
dsQIIWBc9tbGGhtSWgYzS8d3vU0wVLY5CCDF/jDEMtga2cZVy0D6dZfYW1PUGr41qWe1HpUIOa6U
nH1rUfuUAmGgGUnvMYq552MbWQ8ZqDaSKDG9rZI2ERPZ0QtrL2uAImSST57Za9HGhnCczFWJpUKp
ZSDYrNE+gkqqRA6VXEFaNNVzxqsSDRjSIdO7fvGHstV4W1iyd4F627S3FAWjKa9kdNSVekVSHlou
8IlT2hubo4YfONRCkHZJonur2rFqlkkOuS5RvFOvaJ74T0bw9z7D6JYgDdUBXs1f2ue1zaZo8Ikm
9fU8OBEG0Chlkc6fJPEVGzLvjjzVjVCHMvd6A++wN6REyxG0V+OB16oeHvmo40KsCbf/IShkuZrX
Xu5vs1TTtGMMnfih3XHOYTYwu8V3vobQYOk1R2TlMX4vlS0gMdyfupGOY1J8zU1+xJjRG1Cy/H5g
RJCal5d7uQ7DnQejIHR3/+2b40bo/bHXNQkUyqDb/fgHioxUQSw7dpY95aK12rajgpTlaSkvQ3fa
aGRop420wyIGe7PmgErmflM57V8J/1j/9Xxt6l1cIh+0owo2DuVKLNHzSF8aflEK1nDo7zjX5Bjb
9tCDpC1HEZDHPlACQZXIFI5R7WZ4AtZ56Unyd8SfGdFG1ihZWba3sqqGoZSiqfdd8YjdMQW1pJHh
F5aPMpvsETjXEdyDGdDJurMKzPGPjrvyt6/+aZIk4KITC2LNQJG3UJ2rLa3XFLjWH5MJchpD8vsT
iTstP+P6c8s6vZ8ulrO7EBpOnVDDNYtodtg+fWnbe94wYWRHvZI9b4Gf/qXITzYpi2Wk6WdmOWov
9tsNWaIaODRNS/jaicKB79KNN5cB9CWn3XKvhfrNb5LywcZvKAAETVuLiydKg8lfKe2jEj4HIjlu
lESKYsk2qMo7NvRfVlo3Ct/mt04iF7s424W1kLQQcAboXgnCXsPXtOwmdHxus9Djz9RSDiU8+FiZ
KFRQgikHLvdH0Ybad4mlf52NcYu8J588qPx/VCYMSPJRJ9hpfiNl955iSI5UctCHDcziHZP/N900
tyKoazkWkxy3N+7KSqlMrcghCKu9Ekz51cm8k7gC2sUf8oY79eWL9+YZroBgqUoScrIUpu9mea+4
lLjT9XAlQwJYvkg6LJNAFM9x7tcueFjVHKvgExAp2fNVM2cRUkdz5CwT4UtLHpyyianX/O01Nk5c
DsTCWB6hyTFVF2OdCVTQKl1FX/u3F1OfRD85mNLKwgFfaJa57dpYkwz1eiSFRSFC33iMJgc8kR6j
+zgHgh6ti57EGCtljH9Br9JbvxMvNRtgvtk3OaZyw7fK5NfbxZ1KrCzFV37aQkrfuJliczBe7jS+
Tz9m52LpRFkNzZLL8pdUHmykfFbU1xHoon1dPZMWSimA0ue/D8sPRe/S1w5tQqoYxQOVOO6nD3Jb
rGGNLu6A9e/nmWokVPRO5/jsfLn6CxhtWcL0EjQ8aOvc2D8Ba+S4NYY6N+BFBK/XOhvgdsySN2Bk
1AOg9UdY5qNM5OpZKhkjzVraDYcrYcEh/7pJI4Gr8L8dPG2vTnVhNyHkD0cj5DNGwU0VZENT/hjp
OircxQva80K013ngYJqFd4WTQ7313+usY+pCXxpu+vKC6QZENtra+he6XTC2m23tCXEV73AP6MXj
Nhlp+KbXfOjWBcKjKm6iTMA9SAKtfhHJrMK06p7h9FA4WpG4aXVlfuZf38B9TNeqbv0w5J/t0sRS
tCGgNFTUQCoxZZ9cNZ/sdtU19m5Gpl8SVUwqMWNurF5CQxaRXPFiYHxUMpmyH24+b/EpHSTnWqtN
0acHIH8bxj7wSvk1m+2MOq+YWGV2puFJI+LAtiZQTJ6jXfdZqiHfRmx68pv1MVExSeVDQykpVo2C
T3ZgeODNCq4atkyYQRHWqKwn+sWpDmDwu64myCEi5cfrFxq2O/1A/tT2u1SuiZCkHSw8v6HU159u
rCKp/D9VSJ50CsWKjgB0iyYtnGapxQHWr2Ry53qd/hMBEyKZWA6TveQ5DfevR/QNpC++XFAV19Vi
vSK/lUYtojQP1ahN2i+URQ303F+2j0BLMIQ89NuFctWexZ3PQ52W0BXKHXzU9CKx0OhToECr6Ctg
p7E3fOaXjAGmJhgsfTEd2nRUA/TTIQ2I3Zzi1AAMZAr94K9xomQjOk8EyfAGMrVbEMIS69DQdvoa
D5oby/e5fN8mSE6XsrQKoiASyuTm0e2gYCqUMVxEzzVf4ITmeyOvT3NHmPp4I4gRG7XGEnBhL3FM
OfZmBm5/dVCxrY/koRv2BizyAve9Pgg9Qp6vueEe7JIWbewbPM17z03EgGI49VdwZX2W8yOGojnp
ctbaP2Ln+lCF3Civpf1uWNZok3Njp77o6ONbnMlgUSXEcVTVyx6jh8J921BSbB98Z2jrIIrLLUVp
StY9P1qwptc3qvc5FDg04g7ZbMaspgiJH6RUE9Yc3XN0fsE/8d5/qS9AVdG5m6xJPd4zMZG8Re8V
1m3bERWazHfUvkCISZEJpTvcrSzEa60znISVctCIGcbz3dpnwKsjrt9LZMRddN1v4NyYLNRQsevv
VF5c1400U0RdU+9I7kgaicauUU3A355Bs5SOHHMnbXOAB23ExSCGP9wSgsxiEaYcNot95EDf7ccm
p2j7px4mpaCyxW4XvmkOnfcu/y5UpVVOGeSOr8F8ojPdbbAzUWVyKS94kjNpM8LTh5LgcTZ/9njV
Bz4T7L/CIg+fnruqTMylhEi32Hyxlepl8RE8ULxLDjIb2aKrV6KvN+7oXW5O87HjTE9qF8iz2LCV
UBiI9Ewf2Ar3291kbF6uSZlnqzZJrm2kGJjfuPWRqvoFk/LjlFrOaks9t8UI1YW+JMYQikNarnSZ
dqANQ/YE/SqJuKwJaSJhochJCJnVJPz78qGpu3Yz9tq94JDxkKPhBW2zwnR5c9fLqL+UvV+Aet1U
h1+lV3nB6IhokmTYOxqgOMgvnz79OtsAnbs3mYslL824jRSaRtk9q+VPtDlMzdpOjCqu8J8ESt4F
Fh8pvfyS/C54/YKAAXnWi0UeMyYIxK1vfp/5oeXhaIHmGdWzwYixAAw5rYMPZBgnRtrI+0mELQBx
hS4j8m6p1Q0JoZjAfuo0F1U2hzX7WqiaZY7lYHRto0B5TWGd9nJwAsEySUcYKb4NMY+9PPJhVZjO
pNf3edvY7dhaJQqiR+3qjKFv5KjQP+yIsR+sRRedCMi9TCTf/KbU4CKdjlBoRCuiXB6MjjGQB/3o
kQ0YGpRPg0MKsfIS8N0JqijhernOd3aD4byuFidfLsSI2sU9OqbuKRFDs9hCdWRc5Qzdzugn42Na
6rrHGbgCzl8QpPVq6o69sPJfPnVU7t3d0eXAcHsMjYcn+lCvf4RQMOVYrr+PCMDEMJ3YkFoB4D1v
2hM7WpAx6RGopOmN77noomU8ce7NvbEilMAlwP5AUVNVbDOdV/4dME4lM1O7bUGi9u1Dx7zI1EL8
XDJpPdpM/CHtsAxbs6dF9TZviMWHwyiozV+ev+2whDihtrxN4ug0pxjRWaZC0o94+sEcUSqBPoDy
/uhKzF1gsf4plGdEi7q/t8KstExcxqrTxk5uMZ32rdnuNjqqnlb2z4GSftAxyeWx0MCDXhYwnW0T
0PHkcbwpABTkqfzu26UanPYEe24BnSOno7BL5yiKAhb7yeJTzY0YuTQ4PVm/jZPdWwavqpr7/eiV
nS7Ht0+U6cZ++9LLSFx0z3ArAtFrVAgXGeHgsyYJcfOmkM9G2ZIJ6HeB9g0M0V8gVoIPr0rFYeZ0
82HDjSGCim7KHzX6GHUwQmRBbe7KSvjtR51Ka9nQHeoM/pHpaN/M0Epc1PSZta8O6LxDIY0KM+sK
KA7FD3h5gJcMKxREl2rNDoxntE8G5hmzuIP1JC7/8sTPFCQttSqJj45d7wgzXksWOar69jOM+2SV
yf++pFIp3MLGRj/q4GSnv7W/eDBkZasOD/fEJR4b3hWBSMybbRh+UOBgt9MXbQ2aCWp5x2m++mg7
OldgGvUAYumvcCBVdydqaP8GZcCNMfz8avt8Je95qlQibXZgp3A0rvslVvUVJboJu/lqb4b5UiMf
aMEiOEVxqyDGA7beaNitdSB+TzYSROXdvyULEtuMJE+heEdszEdbnSjv4sloeYjh5iSG7fCvwCZV
a63KcRVUguo9PuadzNq/Wg0BDKTX0Gs41tQVjiDbQIvx040Vf77i2Sr1O3d1Bf7jRKbqMtpv8HlY
KHoPkEZ9LYEzkkcixTqqCU+Jh/R/DizlLVuM0KyIFQLyOcsxL4kXlkhuSnYnb/QIOdct1Knzoju3
V/e6bbZ6sR/YtQ/iGg49ink7QdIPrG3n2v3yBp9Op6WGjYHekQTADJI3jz4x6g5ZagcRTJtYaR6z
RhOjBweEZxKy2w2lhZI0hDMl1YvwAIVPe2EVtHHypvClEy7tDy9J7q2U4q2f7mdztuI65dNaO0F8
eGlWYsgq50waxIG4/vR7TBGHk2Lq3GSMGV1YBwdhlEB1JqZ4YpQllpd5+Vxg9qvwWrx7xyoDfUAa
RQCzFqEbtUjq7HwuMtDMSbxsg10bW0f5A0Zz6tLyp0nAEiWffGbmiuibxdwHs1JXkb7hyEAQUDH1
Vxz/H1hdNsfwR1klc9zVQ3kAhizeIDJKK8UT0CWVf37AMMbXYhwRc4ABGWSgh0wCoeS7m46gW6Sj
+EzzSFJMgzWpFEqXGH/YxTXpz62uT/FKqoDKiaXSuEj1atQcQ5m4CInmtMCMrTzpqdEcFTytO6+v
HdsL8PzpyAxcyMdSJXHPHsiY2OThuBoimJ6GeKQLox0O8MM4tpvf1yJPVyEsles8jz1L1Oz61JeY
dD8Z9i8BDyveHwh+PT6qSgDBhtPwjrayDlrfRKckfEbiaD0LvCDNYsn0dxHrFwUS+7pJCRUEjiDL
g2PrwHNLVTmTH2cH7aiwPlNI45ItDMLEj8NUqr0n6JrJkH1aDgCPCcZn4IeKy46a2HnMnm/uOiqm
tZqim4AkyEDziRn4vOdf8eACRDUojYw23kYdcGgGczZY2szdR/ShXwG7YP7Xc/PHyxaF7XNrwiOu
gPU83GqlX178gjZYHbgUvyEZ2hFELEN9mf2m0TNyzUHjHXDePowZNM6WLsAKhEpFVZr3WKRP5sRd
8xIsSoPDycXGE+wNQMIkjtGkReUxM0HoniK2vzmZGnarG3G0DX2okB0kBvzbGiFOufvnNXFS2+rV
ciKi+xXAxRJIcnv3n1eeE6gXL5RHAcBMFM2nCQo5AMZ42oPYDme6IIWEsYHgVNAerE9I/a6ixa9U
TBfrMM/okYnNs2gpZtk8q4Rc1nz9FJcdiI7d0EK0uRlPPB5BnS0vQOLLFSaPN54+/JC/ZHvd09SW
CcTfHcQtOlijBYm9i6yiYsM7Ff82KnsGpgju7ugdq/1cMp42QM1chzreWnCC9qle9GiX6ZpUH5w+
tWYdrOYnsQmXuiknN75nqi6WkbOC5/yL9Gc+ba2TgbDpbbM2RZXzMOZZRHfqzVokHV5m68JPOxUB
3QWMnXD3Jla5at6568Jdf2ITxPp4Mkk/L0tql+K79qRCWVRXdzTQboTV+z7H9PJiQQBZS0ROUgAO
0J7d9ARo/uGNZQ8rQv/Ncunf3CRYhpiGYPHLdd1dDA/zqqXZIA8OyLZ4jUZ8GaUBKM4VlPrGuFvT
3ZKEU/wtkgWklsdAr2LqS3SWrO3Nu+1bVbDq7prvPJerza/KOXVNQzl0l9FM36Y7PJp7X3FvHzyZ
KpncoIytvxkNfK/POp/6J9oolHRsBVi5NV2b2Pf1fdyw5or9MsBMRPiOT6dWo0lWiNf1rnwHQ7iL
lQ6G9OVBINamA4irZDoqZjCTlWxn33PiG5QfPI3STY0mKpTlx7sabU4OsSF2pnYy9zUOcHzuEUNx
OGIMWInoCV8H8V2jwz8c4eTKI4mqxTtquZJUliT1KXUC2lKxJurEcQFexZiV5GF7ZqIsZPKWE+SF
yPm+X75KPYshq01W5YC17bzF7z0CejCahAMeaO2vj2efH+luWlj/MU0fGPCbUf7f/nqLJ5P/LjYW
do9FrEKR1rSiqd4+S1vdfw+/AkFCutOQ0a8VLrRIUBDxboDFGC1kSkwDloXg9Xk8L4bemgIXTC8W
EqDHWrGesTMWqwMqGUkdKmQs7MspMV1tGUCSHetZe1TIZvGqCL1nUIxp3JTthTOo7VVa03IbhlLk
q7DrDyqGPsQLyClAPWTld8qIH1zZpP+tsbXlnox3L9ZebuaORjN7s7uRFhyodz8npEoe756qpnfJ
7He1UK0BrlF38Eu3DzAqMIe3HYryzBXjvtewwOGujaBIRN6f2cZs13ZstPXJISeNBC8l1ku7reSb
SWMw8Onm2csWtkFHjvw7N3a8dBwSnehtbcgNiYcHmTmCgpMRce9s35Vjq+Ziw7zio0EQlEYGJzpC
X/UV4tBk2dCD67Oou1cmc8fUUGAHfZnZbhl5IsUuO7Z8Hv0z1+6y2NybKP/8AXS+2iqHAv2Sp2D+
jxHmAvFjnpyXZ9AW9f+3p5QUHirBOgHJlU1Crx4uAF3o35jLpPTCrI+YVfUCJ3H8JWEYH/0WXfRV
WpDsreqzUZVc2Jx9cptBz+il6YdEUrlPy9uZluc+wOpHduDMYEuWL7pQtPhBzKGkyJ+TchV5WxBE
UeQnv+LgIntZFU99KmmNP2pAm5uTmLKC0ik77xWJMdOj8NkEIJwlCFiD1OZGGjwRfEAdvY7D42zo
OwlIjqtqZtF5Nzk/5ZvG75HRse6cceK/vBG8hpbl4PWdTjSp+/NbEyU48dKdg0fqEjAPQTW/9yZC
KcRDFc2mM0g2Kv5ORHFnRazjEAE0sttiX6g0vpeQCXanypzh+9pGLTA81dnksINSRS7o2+jh4nsC
JMkkPsTFLo8IAznBdtN5/pU5BFLcaa42uXFeaQ0Cx+cw8I9wZOLRupyPx8rdqiZFeHvrDVASFtFw
vy0w56CSuZp9J80PsyRtGmLDqFBf3SjE/jPuhPuwXSh25dROevz79d9/VOCsZYXwJOahzE9STKyU
vzBVq+VRG2a6Xi4VoFAmEIIuaXwYqSOKIOtXljEkKFrEWz8q8eHmHQmMPJjFaQ6Js+qnIt/PAnPx
ekNNStoLrerTJeVjPKuF8pndea2NL/WVVW6w1aFU6zUhBuBXGh0Gvuv7mkNS4PWKIdphPwx1pvS+
/R4aKLCPXLQH0N9550Q8/d47w2MvkUUGClVvPKRVlHsakCbsejUYP77dHkFMzjT+JyTY848mrY0n
fJ7umvcO0RfUz8CnRnf0cEgouONHoTkn0vcYMlgt3bp4o5Xcy9TWYL7rN+/5TFw9f7jFEtaHHxCI
TsC/Ybz/lqi4GBm5WcF9gJ5tFuiqb+BqM5atVF+U333j6VWIenTtyvDhZM6eyekuEl69/bM6u2Ko
3dH19hIdp2xBiR78W3o5AEm9tKmebENF19lilRUV9ybyVJXJLkHM7lLTsSPM1utlbaXaEiAS0TdE
9LIsfJ0IxX7hRFEie+tb5jj6LD/HcQHB2Xuy3MyyFokTBE0sQUZcZ+HlFt9Ee0YHMgio6H2wp+q8
o5PNTCJOoYS7zWvpp/OM6MJOz24yjmnvYeXj9TH2Li8QWYcQBDscJ0zNpZVPG4ZOFFSZG6ZDW/PX
rWQlNed9fVTP8z+cN0/0iKpHn1Y2uRrk/UeV5uKWqn/9YNYPOv6kO4v5isXSt5Q4HplpjStI3rw+
EkNIWLyHfIBi8DHAl+TA6djmqjvFlZoxSPXUaQoug4znrmVjk2ws1xwOfvWKkKdXMrvJUhhBZtKe
JZI8NtIIsE/ZuqLF9SeQLivurr5uqtVI/UQ02A06O5ZOu+MqCfhaOHna/WtDM+xuFxohAs10ub96
cNDIKjs6wmOAMI+AY/a/Hm+ZUdBORc3jA8skZskPfvGU4IC0rLWiE8d8MQq+yXYKDBlgUxyai8iI
astVHeF4Wb4sgJNWxYAoI9Wdj9rKnyg0Ed0pCjrcv3XEju6g7n/ftsss7eBeQ8WBIFsa4fAuvPTq
XSiwtrP3yCXF7NoMHsNdGuoLYDwAdT6UlM1JolbtUGNTxz7uuPytyGBJlZlQMrZBDR3Ghfyd/3jk
1W3mUKbhUjWA+rEB3mDAzLGGUJnIrVT0KKMxw7L5ju4V1CuBeJPRfdVHP4qWn2VzTkYKY/xG8zM2
ubyRdlLkroWlDsNiW0Eb11RNiHcSMZ3tstrB5Y9mMZUoPipTN5l0onULDTSNwzlfE+zNQsW6VjwJ
SXnf1Mqy60bj1bFMsia6lkykVhCFH8a0cSj1yLxozc7zT/5k1iRRelwpUjrz54Cd54++2BmLE+XT
8pYTKXcLmDWU5C18/cTk7Iqt6+aHH+i0Z1bzciVucSfWOApiFF4bSGEvqNu2S+8v4xQMoqzfVcg5
Pd0GCYQW1qZh3bNyBE56kadiV8FzxZt5yqdLOH0B8lY+g9zDL9/2wXZr9zi8r29uoYnXOzshq6MS
tZXJTK69cbm9/pKHNusCsvVZeVZdPBmcTSRxfqfB+kg5M221Zn5o8e+w7N2iib6AxrHjxiZqNGmh
3IRntpXsuPyAXtco906ut4BVSBOgmg/hnR8AAvo8a/S3xDZ3DawDtULIEM7HITGXBt1Ew3a7Na7q
sMYVSGxrLfjzyhxu6AzeUmEqX4UCGWW5mSLVoNAKFtD/dDAcbPJwQQLpm3Ihl5wHTXpXJszUtw7E
yfBaIRVE6QZVJ2qJnqmkXgU82oTPx60HcmTC4TwLCmpKQxSefTY/OwLUF0Eai79gstmw4YRvyIFX
G8D8i3E4QiixpABKXT44++Fl3dnIqY/xRGgQaWITfIjph0lrSgAESPlHlXEEKP4ZLF+xXwTze1WS
iEWPbXm/9iuMMyg8IZosBkzYdkAGoRgg7Z8Ae+Gd7On1InGLVWBIpSYFnvMirK/ETJZHkMySbqs6
AeBgt+qCEL+PUCFPb/MVp27o15FOdBhNeThV5DLJJ5ELV3XRhtZEhpAPbh4+EI8y7v5jKxyJGusQ
qtjabqyQk186DC5z7YytQnoIwJ0ovTpPJqfGBajJYJe07fK60yLcANHiKXre7CvcjYyoW7jNHMSK
/dxmXDdjcN1xPEWQUWPjJiTVnzx3d1bfp8/N0XXgls2aG0CAxmgNIDQT7FARi2/LCbQjRaG6HIQY
U90ba84DoIRgKGAx5h62oZh/7HqAAfYIoKRfd9ZK4RO4okpFngoXFDA6cbhlodipJ12la1dKY0Z1
i147gkpMBt4yNG8Wsa2KkgnFbHc+UWEaURTjK6RqDwe4V3R7EA6/Y4Pgc+syHIqrsLfKNzy+jK8T
2ytPTDCBnp1hS7Af71PzmjTr8ZAKxojX8vjWlVvdhkqb09SiVjX387VsuJ/7nq1jDbGej+JqYiBs
eO98XQGKEAuuQA1LpUqlqQMgj9IfwYl679HHyNn6rdSkA8JcZqXBTfQLO2UVqpGLzhHDOjb6h4jM
E8XXxQLTYBx5hD/aopw8uOGbgREK9ppABnO0eRYfeeOp1M5kXUcdiEwE89Kyy0/JyRveCg/hJpal
R8jTTBKCTLA1uc16VXa9krYh7BOboSqvyDDejpZ4B+YcLsYDruGfMkdT3/kQnmy/p/nBZ12Olupr
25ga3nPwqM6db1yOw/vdMbjQqUOQ2xHbsDzHFf2e1Vujx+8H7t3yHMx+ZgyTruDiN6vAHt4SNrYq
yGyqNIpwwBQcQkNcKVBtcLWEPzNiSIu9cFsXfitETKnHZ60WVJeFCLZXAK9igXGZJ2vPNDP55kur
keB0Oaxpwy8NWjrLYckbW0thlHnolSVqHKFQ1NsZNmxJ03wAOwqIBaux7E0+RSXcmmYkIl+pXpug
xM+iIKWIph8qAOyQgXATfk9YJmn501eY/ZCxLUGr9ZUXHpdEcMMBCnZ/w1QTM2AfGblPLcc09NRB
tRrwn+BEw8kRD3BWKay/JNHoNwSC+jJlsj7rQPQ/TPtTF1/qNUKh2VMOM1rnOY4tGlBIjrAbm2O9
tK8idiLnsu6+TtzBG5Zfg5ySEnN5e+A+WCMIWz4H5mVl6vAz02BLRkk4wyDUy1789bAexL4FJQjN
KYXpNdCZDfOp6GbHu/UhqfvRPodWWNrFdb8HDvX1viOk5GWJQKNwy1vnAEk1uITXw+xuKWraQO9P
gBQNm9FhJugwSUzhPQzg0ImwypAe5uucpOQRURz+FM3M5INW2lwld2/Q3V/4PPssQor88MSwx6+2
o7PCQ5HRR704/3mCvlqWZ5TC5WmQ1VrTHHjI7M7pE8qDGDJJgu32YfJjb6CkNUyJ09eo4FUzJxWN
Go3AG7Vn8QsTYWbA/z9+lPTys0nHJ0SGhkt82Q9hX3BdWqKPunZaVEPOAzxv2jhCRRalhTlySF1A
7z+lVnJoSpFQDln9KeBuOVrhVOF732r7NlElkFQcR0aUqQta1eLe0i2BFbF2Z4p0lpHDGUPBxn4k
GIDb5zpNFLdc63IpHm/CU4rE3Xy7b81nLPauag0pAfJ3wx42An6eY4bAHvByWFXK85VUSnS03AqY
+0tdr8fWntlXJ7tS64Kj6hDmU+MyjGKzWT1eqBzladU5DNMLI1TONWvOW8J2tHaihX7HrfG0MzJG
BeT7pCpbf7We0ARRxhderarEVZsOyW3PirQ+3L5Or7uWVUAvofhoUMW044VO+WRkN+7YVbI+mxb7
ifNKmzxbrYToteJl6r+nPr1CaY2nsO4PJlH/drJ4JXmEoehwnpCvZfI1BeYgrx8BN+McycNDHNxY
Griof1/dg4xp3EijdstN65Hc9GAMJQFgekd9Fg3MdDe4ESxt3+WK0WSJ3XIaMMf5dUXom4H71Kvb
+s/JDmvoIzVHuEUaBCwGDRJOK2dP3K41rYswelghdplLAjg3+KrEuOlgdGB0f5v5kwtw5Lird3fw
P34Q+ZBCQSI9ghvqetmSbvPSCpHuDJacKCAklgP8uw/IR8DsSRDH2ajLauNWnNp2EzwV27W/F3xX
614F+sR/VVGDYUfjKXeOGurKLmsNL+p8FEO22Dirovvt7KVtVRhYGWypMuLe4UFLdJamN60DEHmF
NLdSsUQnVatWOiJwwehTcdslzO8L6VrZHy+XoEt9FCRsJxPCtfccK3xS0aFWikwlIvG/nm6VUcgC
Djy2IPeH7W5ozOxW7AQLLwukPLyGvtqcVby614x3rXd8sYK+v/uS+abzxO6s6QZkWBkg16LvflCf
hcEuY185hzXtO3eOXVMxPdFfrXuTh1+cbXTeVWU1WGovIY6d4STmW76BLf/Mfz7bGiCNiJ6UmV5E
WgWeQiM6qvTnrDUnIZ7LHLV6urWwSniS+1IgGZtlRvoCLxL0RIRPyC8cOSjHbX1PhmbLjqQy9ObI
1xUBXUpb3a96Je0kDhbABjVkjpCvjv7uGoBfAGaG7M5/frI8lCW9BNZONUoLSauLF0AvdcBksN9Z
I15McQoFk1N4GlpD7JbhL8FW182aoudYIyaOt1ERclvvkiw2Z2rcG8jUucHDOJODeB84KnMJiunT
B4QzxobSdaIoJmhA2wqqJgX2ZR6A74wd49IOEhmF/fNs4soJJEGeNfDkaqRTV2vOdvPSJ2gPMFdR
IqL1K8wPYmUtfumhGsnpHqIn48ySiRGsTUCemLMgoa7FJRsFlTgtURK8lqKRHyKksCn8SGIkUzfj
SWCYM5+tsZCq7XBWoJXesNNMBl1u6hIeMwTk6XZeSu8sZf/J0nloweNKTxVLOtQtUDPS/vaYl//M
BY0K5yimeHKK1Ve7SPMN6OlJPbNmQY47ySU3OovbZgiBNeVZIR5B1zgeuPhfg8HpoRihdgHovuVg
J/sE8LN8+Pf5ma1nsAWveV3iJVRi8ejy8j12uPCb2IfD0+EcWy1HPCHOsHRh5u2MyOMSrdralVxB
jiLciH+1Vz2E1CjvbnEz/GwVcrsohDZsxP5pGDHriPwQ2qwf6Awc2SWC1tCuUOKEYrRItNOVFsop
x3/BDh7yKF0CsyDPQC6uFoF7ThAQmz4lpvA9jxqCsTmn7kNiN1SEl0XStt/2ovFyatqueTlHlupj
gLrXpXtxz3o8XSTF4x2/R5tkfOqRHRnzHrUfaTbcodEGCjD+cOqlHqtnmlv/G4DVmoescnLYuJpE
xq/G4IRICeG+OMQYyaKgOzGP6xa9HBTarOE4hh5MBa5i7WgjBtLO+qqkBtBH5+oFL/gXGeDwwFF7
Q+0HLc7HidXfELuC4olYRJj9DGLKqcR8EV1tHsFTSLp0PiVh4AxKgj8Gu7EMmGzrDCE5AoWGglIf
o21Xy65gnborLudPrW5ymQHXelskiCXlB0KeEG5Bzo7EOCFOLK0WqCFi7XD9oEBeBc+KnRuE3MBT
YfqTANj0cJU6HyYVSkWvHNRMKBcVwBIXdtKXvPyGc50eraS33p4zZRrPGvW/c6IodXqZ5IqQ8jrI
9iT7pJfHvQp+BlvfUsLXj/TYn5nOqD9tNz8d7cgXtCd+F0ZuSTzRKOsM0AtRKjSxVk4u1ga1OsV5
rygySHRx1ZUZlMbAJQBL0ecBqXQhBuGKFZ7yewWHg3Vy7gycyOjJHtk9PLGtxcgq+hXEQYPXi+bh
GVM3lgQ8lhDiP7K2yVHOoL2RTccmZ+UALuOw1obBMNeVCHMKmk5K5Zg+ENPAqSR1uaB9/8NwfWsE
SWiqEN93jAyI91TLyPmIQfj8jVAzC7EujrKOTl6pznspf3fTdL8db2NID9eTGjtjufvjFSZ68D40
6V+/REj8931P806m45YCCyZ1XKWyrHxbFZF5kPJtBdPtORkTT+0SafIV8exrh+TTrbrSA4tsvlsi
cWSUP7aN6iE8E6pXmpauWISDbZ3YwDobW4YQg0lCrU1L5x9t+AQ9KbDRhy85zsJcxye4EKER9ITV
7wERMOGu2iGHIYB41iGRBsG6TTVwAjsX3LQuMxgOwzreBH46uN+26L1xMTnY8wTJubsPWZZ40kYC
OHDRDPkjBTi6v28e6Dz01MsZ98qL0iKReeCD+WSzsJPUEJANjoMClEfp9dDZ/3SiXiOUjxunzrsz
ZaL3QhiYcOmjLOSKNnl5nwlIzNR3+0xB9a3w5iOoMYmAViQXgHDcpVA+RmmH6U5a+LuUWnD09yeg
ANmnD9CMVD+vfdIBgZQ2TDKdZE8XhGBg/jEoohwReJdNfS/yAFe9LfKfy6Z2RxRxyLtkkN7EQV5B
QVJZa2lwlGgJwM46BQDOULBLhcBeZrHIZ1b9Ih+SMV6gvefGZIE/l5nHzBzTvfHKrcc8AUUEy35k
SJGsHe9ExLQ9MHXADMCYZSOjqClsMy/gIw0/yVjYVyMgIvIbyx2T2oNhYLv/0fyPKuwnM2ul83rb
OIlDZeeH5XWVCq3v5YJyavuja3qUZmkwS8km/W04RQodA3znwdeR3nIZSeW2/8ArVysatMu0eVB5
1kTmEKD3GJmiB8+bdc6taAqKgcdnmIAAI5LzLdQzyU7g/dOfIcO8SxMeiM0sVhLgNIliELcGnfom
YUP55zHuDApibXYfqSAGrzXhw63Hx/jlEUzFrohLgisgSqdbIAAifNe3krRceV3Zwj4lVtp1yt5t
LGBoOAjFu707iLzqmf6/uMBqhOWIolD4HYO6yV3FvTZpBDrQk68Lo5dYaxcDauqEzUCNLGPeWO7h
lHznoKtsTZ7xRBnFH3a8sISJYJmpbPnQ6pLDGLvroUjtr2z4jGYEtx6+Vs87WCBzsN6rvQRx5mOs
F+EzKYkxj0E1BoYsz97ftJwsVuUiDr/5o94igFulpoAyJZCs4yGw9EaAERLFgEWpWbBGiZ7KzSXG
uW92CD5sFajJDxZnnbr5hNHMK3jO5LL2dbWO6SJjNlEGHhRTtNT+/1eRkNM6an2CvAaQrDlxh0CA
jgxqb6Dxca5B9n2GOKLqgX/c7Ao9OyPzJQTu3Il9xnPef1jCSmXLs/Xc4PcJ7o6EYkMcFiT1pZfq
UaOB+/Y1hk4SJjB022uVgFLRbS5jb4yFXpYhVG+VKEeG0jlGzZ6pqLQGF3PNFfu08Q3ViBFPfD/V
EJaFYPT+gK/pEnJpPmijsk2GjfI5bPgkdQT5h7KC7KabV7DUWHwpZnhwaTJI3dWz5M3Wvf3DqU9/
kZSxuWhZc8iv5yDYpHsswR1B91610vTch+ZvGLa1bh/whGi84wMXUIYORnevhsiMy0yKw2M15oaj
2gdHa6s+RRJy7Bs1g1nZQxugUR7C2/wzWsK+ynC/AKDs1Kt7z12TMqEAZ6bhQflOa/fmglahYdhf
cI16FNR/9RxhoAUhUII2JJhoB7FK4YN8NE2Q9aUe8GUBADc0YHcUDdlbXS7F/2pVkS+ZZHHbSpT/
pp0iOFAkucLOqZ0MbdcGIcZ+w9a//x3un875YAHnPv8qfWkBQ6tJermfDP839e+kepWrXy1LyZsO
6Wl2kkp/b3kYostrSbj2wRqpzFuyeX5g4G9jiU1IhrOpRXRfyDPA/TXBj71RdwxCm3/wA7d5/FeW
KZCG8H/p06UveIfDY6uPB5f13mOGZsSVKN8HiIYyC1H0gkU8XcUBRJFsKe9clmdJLi+XP4jQm6dZ
FZP1CMHzff/ZjVkOikTXbAdiEQaBWhdgFg3y9OfgdHSWVO0gjwej/pKkuJImUaMbVxocxPQiZAPa
B8ovxYR3Wnrpo6icWpXlWHHMkWSGBKQrdpMsqS7Le5UVTeTGMWx+0xAnIi0neT+q61QzvRmszpci
w7MGSgp3EMz2HVpcArkO7i1lEXMIhAf0+IiB1FdbIrh9m8b2XW41p4v4x+04oWdhZKatUiheOZk6
Lr9zsWnFJyo3ZwO5zTLUQfyY1VV4sq2OngN+EufyUGPYtq7kXVuaQ+g/pezP18CV48bCTRbtcgdY
qiWGhz28V83EPqn3T0IGNtV9LPDAgrhTte0D9jvrQlZ0AJZf2aVoICpwnT4CIleV7xDFZuVZIjYm
Kl41cgBUvRfufK4d3O1eyxMvqlqiT4Uh4xdUQw98w+3XQWnjatTAxt9hQGFOqh8wvVvZth6Ck4R7
U4Ey5Ab4XDbkXnOCoJpsJOnHCA6SH+YOFKCtIRA7jXmcGs5z5jRP+ya6l8yOiHDywZMKaoAwlEoV
unNZFWJBlI+Uli53HI5x5NzJ/pr8UpJL4oNkafOkmVdwErIZIx2X2VyLVXxUMan+Pz3a7rMg22hv
7sK1m3H+v34B+CoY+gIdYYK1PujCaeY6Ab3uUSn4FMrXNqhmvIioFoxBExTGvvU9arkQ1n7NqRqC
Ku/1MtVyNNIjkvJAasgKc0cXCtPXYcdt1Ux9IqxgntxXyej8arwiE8sSaZV6Xe9cKxgsXd4lFAwO
H8yuKv4ajt8blNHDLh9YUFqRJpLZ+8PcwwI+sjZH0+AaR5//GEZ/H3aINUBZ7PGzNSkeqVZW5p7n
niy6Pz3232D27UJyHTWJmBfa960W/1jg5JTFATakpJys7acZv7FA8vWb2UuvgC14QdTya29kAglz
WUvckjvnHm7khdduUz5ZFDQpdX8rTue3yfzwVEsCAFFXFs2Ce6YHaRqJif0Oma9S/0bNA7wLkSvR
uuF/mQzEV/XItUUZQpEHcvb4On3fp2xW4+35r1xEcvDawEJm9bgCAR6o7wMQiUMjMRI6a28HZTEh
Du959mMHdb3mGz2MbkJlh3TrP1GZEVefR4gDW5Eg13Vi/eZL2YaXh8rlp4BjrQLKq0bWKtySodx6
fi5mIJiXgPduw892+u3FpCbseTlpOjk36bt9HFXrCmKh1mLLbDXv8eY8YkrbH8/Hp70MZOrPRrkG
GgOQRemrnzqpvR38wS2RFaKDOodtpxm/Zi4L+D94bnBj2bTmX6L/rT0tDdbUL4GQi7ZrOditltgp
SwaDP53hDSSEW1nFc2k3X49OnPTfJYqyGD9kcDWk/kv1NJiZKel/SgwHoiEE62xW1FMFD3wTMBfv
KtmSJPyoQOPt4J7QK0Bydt2n3hxLjaNrCzRBQ7W5F8y8e13QRBkmH3oe2DLi1OXxiG2pGMFF3LGw
bJrMrjQGrCeLgRFH0qZWcN2eD3cA0vM2kUobFgORp8RHDmsYgeh6l2aC3OVes/1ZoSTGZbzUoeZD
B3DkQcO+MDojvBSIzNJzUGaoQVrAXuK5mR7v89RqmWMsQgw+vVNOwkpDQVCA0MW9SBt7nmG++/ra
wVKeLDm3mNdYrdX2j8XxXMF6Dl5s6PeT+D90U8fvRzB4RN5eqBUzobg/aQ5DRZOtWxdbKsJ0lbp7
V2vu+Y5lo3BsWFeLdtzO2VKfzwTlE0ggH02j4v2p3QqIXf78bMh9aA0jNPgCt/Noxf77ybFVhJl/
FzFxp4ta4NAZSDxQGBXURp8szV1Aq80zxNRkVTq7xuXb0JeFxXZGUV89QjpKqaUKG3eAjUwN5AVw
FnqVpIPccKu8JD2IUuoSquJvnCCYVj26Ov5Xhn1qg4rUQvJKOqnyr52kXCZgqSZ/JNxrOiP1kZyf
D81vAJAGu8jKjp4sy9ql7DyyFNSOFo1j7x55oNe1eYkagt3V5XQfbq9Ost90R0d4wuTAsFMB7CcC
N62yRITJLI/jHPzuikzLF81zIIDgKf5XwBp4YLtIh0T625wACtaUoEWAVhk+COlyBBpUMIjJvgIs
8nzAXOd+/vceV3XZhH677tHL4KIrYTsEOV8dptimEHNnFDsH/RiOFUdF7jfydB0Mc/bHgzBH4bXw
NqfBJ6y9j5wDzuEn+ufDRxLB9reqoTYJZ569X1ktPn+Fdz9DM1Vuh+raYHKoSkEVlwIbXYB5LcOI
Qg8850LVrqmXWUcq/Anc7JIZPofdSVi91ZpKUScuW7maMG+UrxDq5xoaoEDopqSFtNcA5WM//mXV
xBHmXFJe/sK2F7S3ZgRatlmlhTnEHH3Zv7Hw3i7vAQQ4cYxNfMONhnR4XVNqPhckl0KtltWBD+ci
wrn3yFPhth5KmU5E14QA6yGbS14HCyaOqTP+glOXuol7gkhQJQIWgPKEFJbUM+9n2SyHni+uh/bU
Iuni7DJCiwS9yeTJTwahKXbZJDh/S7ciVCD7ZSKSqfHE4LinOCjLlQved1xEcULxb2P9uPV9SzLO
e569IBz9XODsh7wZySLymjDFNxcrVbIcBTtACz0P5TiRAXIIsOuvkUEtfobkoFjEO1SfwUoQQ4e/
MR2RAcRWAjOYBvJXLt7wDbHjEO6jVGliSQRNIz5rNJ9CdbfnOPYklUdqIHHXr3xepFslXxx2A9I6
/lOCWsxXfcxCrMKpS15zRofmpGtHim+R2dW2+6Co0N/xY1rpOAvjTueRBufkLvuvkS+g9f3gC7JG
yMGX0LhDNHVfQUQZg934oM7R33AtnE0Gcc+7omFBdQ29sfaTQe/XyKh/feL/4tKX7sjVjpV756xl
UaxnHIkpC4VxGJLupsdVwqLRblZ/5/rCu+dcUp1vcJO9MX3XABQRluVZEOYMqEw4OoP0nRf+Y0zT
KoJhQNfR2Wd+b1eIZkBwTxYbKZB4KrKqUYcMso1XBGMyX+NbF9XZS3xMYr3disEmWIbNHxC1badG
MknvQ0j7EvOjTiYUX3zJlpz3tTaN7RKD93uKX9yT4o4/FnqIQW6fHUWrgTfO98k9iTDc606ZNgYy
k5QROICSNwSlJgVpw0oGT9IGL2TKD9zgFtKbplNZC92ZRTK+21NIui31alGHUszx+Gt11h4IRRHf
epZj8SMLFG77lNQZcR+vcUrYF3izy55b5cY2vOR2wmioZ13hjkl8Wxtr2rLbQ1mm0sVdmSzurj34
QhL+fzy+3X412Cb6OE/QoEs3CpNCmjuKuVN1pH8mguIufKqz2tvOl4jQWrbljPeG57EqV3blo6PB
U3Yyz68DYm4FBL3n4BIo7plN1wwu3w2ybJgaMg5DEzHHpfLguVJYJdeQKkNd9OE4FPXUAeOPzJ9m
gYxpFPtif3/p/hTN9LL9jMQ8veibLdGOwSG7qLCmMBFaj2h8sgDMLB8McJtOQiCTWd2WmpnLpmks
kYycrxrTqPFYaeaqLayQj/p8Mv8dkvfD4I3Us2GIUOMN6TpYRb+NGkejcs+aoFaro4Cpr8WTDs69
eh0YtdWjJiPV2YhRbXmqjqHcxjpCwFD2EOsFuL0lgv8K8AwZxQteplsKYJQdfisZij6u+4fQIfSM
t4xd8YFD+8qC9MrwN+j+QWPTRYXk+6UBPGzzLhE83HUy6P4RlII8LGVv3sxoxJzjGdaZz6eKafUG
HS1481mmAZtg7H8G1uEZpnpSHo+JApH6TF+MLFtAV2f/oY41s4Bbwu46SVdyBBZeCo1HsacyuHxR
T2+qrAHqk0BoV5GNbRzdkX5fnrDhsaMb4ASpGwP1KCNoLh1ctjD7yRc6AjPomfdLuBB8j+pIBboJ
V7Pzihr9mfpV9YSqBeDlsZAV7RzxO/oOTWLdmHNCcOSERWAzj5/qErWm2LaPXxww+/mjHw27Pq9I
oBCC86tuwfmySAcwINol+gLjJmIZMlSS5GPQ6zmqXx+AHd9MtQ4w39Z5OKIJ3xdcCnS9G+Qnpok7
wTFx+BzI6nzwUgXiBW0zcD9X5wzfGKp9i169VvNrYJRJZMRSqPBrD62FbG8G5rjexeT4eR1RApLx
vOcOSVDgyvO08dr3mV0StynCihf9nmxptWeIuFqksXfiu99qhTLgRcCUeqi+9dVW12/6Se1h7WO9
U54ZUUhaIRw0goAYJYKalR5hVFnelPHmiUiNMSmgAR3mnR9jargymp7jAd7Bv612NbTUH8/u4zTl
PDLqaAXg09hPQq5GZqgSX8kfRiSZIPveJjURKd91wzKMT8PT08dFf8jOVNGf8iUFRQsh8/WKHguK
ncmN7W5V2U8RoIhKOOk5gsoDu9oKEXOgwF5PsFZjVVwIGsr7ICaHZmwCCB4Wy+irZ6KqQXd45T9d
Jn916L8pFJXkdJqBvp3E6JgPZPZajWy9u1oh81zc1ddF9Orajh7CwxRE9VpzS5zhbsqmgr7POhLs
4B17tUAxDPcH9YA1Vq2XbwBmehC1JH/x/CBp0U+itCvNXKC5AQ9HlXepHQ+nPcuz3/5j+qFwg2UG
Fuijj8CNTPyLPFpyl4uJQthQx25i8leti74bvKWmzZT1bsors3LjcbCIJWLvc+r4jBMJxOORQeNe
pi/8sewfeS25zQbxGcR1Ocjx3gMboa7IFmCvWljcPl+gqLcGCSLQPiHHf7CBfFoszx14Raj2UpDb
edD/jVWl2AT96kTCPIGFzGSDKlMeMvftTgefcQoe3D1ABY3CfqBfIFgANRwarvMG/HSkr7/YR63R
MQUcsB4dAGQztENLndPkqJoj7UJmnd/cX0xMYRPw+9E7XtLqoUu1RCM7OPcLqaBuM96qLwOGAqed
lZwPTSTXZAlcDLyWb1ebSn9u+FdH/6zsCaFOr3E3R8jNangB3pSxa6aTfXPWFmIBL5KEt5+HioWx
iNCvPTXc1ZyAF5/ceF23SDiwdCFhhg81QHpANNn1tnYNl2pHxyJT7xpF3FZbqDfR0wqKXeYxfKP2
+2AWGtUI+Hw/ND9UEIAzk3th7P3ttLZnMVd5vKeMKKFgyU3M/JjS3BW30kJkbIjeU67Y9/ZzK/mQ
EN9VfvZHv9/v95iZXGRF0JBzoVBK1VyHk7Ji5+rje5aqfA4m7nE8PTJeWgF5FDnLPF9yOJzkQOba
tZQqyAF6XD70h1X2AZghpx7eeIM1SkbSpvBwbhXQ1EP/maijIaWEMBA4Dt/ZhHA187E7XQAHoKVx
GYaMo1rTOWgXxSd/8JLP8bEdBHpJ77PxbW0eY4k/M/mhhQBiUUSexBviHN8w3lJSYY6kfSoz+R8i
bnIA+uT4UoIPkJfOk+QdBDBx6oyjt2M3Lk2i7uCEU0FIh7HDgUM3VXG/ZgGcuJEkAdyts5fjvRUm
Q9qiFGSSP+LowwTE5Ofi6T8VTzv8rfwfXtTXoMMnhD2d8OHp6GqGJssc4RXIlkUE0hCmbWVbWp+S
/RRs3nWAGYLmqs47zWLF7yPcP7gpcpZgscS0z1K0Cz1/Xaw6D26mPPfEA6DeKZtxD81tsrXNvVSO
a9VUWg/etkTQ6AQkTaI2I2z8tIZUn+bYAJgUvmCyO7XALPHU22acHetgiyx89niXG62f8Rto7hPp
uTFb6FqWwxMegp3alldnnONI0WXy6mwH0gkw+iIXXg3q1uVtVwzJL+QCrLtIF0vknhHO6uFb1AV/
I2xwjYoAkEDMYo4Y0ruR4nPXHwI1UWadkZjI6NpIxOficBgn7cYERhODTzHTDFAXUD2rOQSSl8xq
9FfBK9plKShSPTDWbiDlEkSsH3mUd1/l/cdeD0JISIvnQNfzeVs/k5RulRsCXv2XW1Q57x7iz6e0
icK/Lx9Ubw70yYYkzdP1jljzXl3FAHKnQzm96w7mNrVVlH48BUl37aT2eP6ojKLf39mTiVLC9RTJ
Y42Zjz6UpryAcobEiP5VlREoSZIEMxTMdzKVRvqaUXPjBozwRapLH5CWWLL+f0X9vL/FriuIfmnd
1qZKRK10hGuRoxB39w9lIyiEthU+mu0Br45GjbmfPPSZTiXHtJlMhomhpRCM9Ahz0FGAS8uV6TvZ
69WjNP797JjX/n+MK1dEjKXwn93zF9VJRhnngq/I/koWowbiNwBW0AuJh7Tz9gPnDk57RuQbUL17
2UuVqOfLwTL4ZeQGMYd4m//rRDu7y/QlAEfMnde7JhfHxfapYz5kdqQFLWM0mcfDZtYIhE+VIVDv
6dj/9WYa0bzQ8x3RTCNoT1MIzkhXX2EXd5TuSTzRawvvdT8uNJZWm3RCd5jC/jNirHrI7FbcGXIL
zQaohoHrIDM9LmIeNGt8/r/Iju4QKoy723m9zT50lM1hrM5Xo0X4vMO03d+yfYJ/9NNb6gzT+e4d
vXoSlbBBWZ2BFu577HzEbbWzZe3c6G2TjQQ/exLBG0bFlZNAX6eC55i6p8+2gHMtbEG8O/mX6se+
japlBVh1eJMnRVqGb5wz4SiqqlI4qlzMAznJvsr7kRON/V+7srVkaGPggettdw0tFR4DV9YRUJD/
uXoZiuIbMOiMCX4eRnR2s/g7fQSQU9uQVeKcBtUdB+QcUm+CJl3DXCR9yZWH62U5o0IxTFVajbw9
WLztRf2tRVOs8+7lq91zkkuT/9UhNV/sSlNhidvQr1IeFmAMyC/5dDqFdkB592HLF44ZDvYoXg4S
HQTdYK3REWg1KKZ4Cm/Pp04h9sbO3OWN3n3FWOrFqXkGHBhhbcTW2MnRfFNhzcPGGo6MIw9vrILA
4VK+k3PFQNx+O8woFPr0twW/83xmD1eL02bq3m9Q9p57SC6SsFkQMUeit9fjV2Ci/k2vN+SoK6VF
0R/MhTs/Xs7ctTyUU7e60bLbukqlQLHiMRtSa/h+cRdrWFSK/gveQhV4mEyeUX2c39cnE+Ny2cgP
uq+nJmimWOFFTIuhpugcCf2wW0vqly2zHGZ++1O+4sFIDfQ3tBjtcpMl0utwwPk3Tqz7yyjcmr8d
GlvVcV0L7a9t+g35tJ30O8eB731+QxLHT88oVGv9Lrk4H+K6hRkFdMQ6f78NlM9ub5jC5UxxzEWE
ajIYYkzjyxz+2ep9aNgZftWlRFJuLc8NwNPoNVruhxcB+QegIGSoxKhGZYdWcTsTDjYQYN1B+jW1
qXvJqq5lNMSzaP1tw9kTgwKmmSjCRJk7nCCKAq050O0jLmt5dAcZWNGTjf/6l/VcUpspSsI2kczE
BrolP1IO9+yVamOF7gVMTVpTYCwwUTVaUjwDQlDqI1t7myDL4zjYdcT9voZsjHOuvCgAVNji6XfN
efgK7zh+WG1PSh7tTh4aP0RiEWwVKg2lEJSFL7vC9WfMCug90nGmEpk5V8hefHgHqByK7WC6J7Ss
f84Hd6yqvQzjl/R5yIoo415EJAZTFIM4xXIU82wMzgA48/Gba8Z4tjWKVHPbHl68hWaEMBHfs414
hIy9CLkSmQd1p1RR+CcYH+MLhLShHMxGY2gpxSmQdZGkL2XO5/bHIY135OQm0xN5yi9IP6b2akX5
J/rgYHNM50oxVafltPbvZlvUP8oLrsKpHNG6dbh+1G/SfyjsLy4AV45PNQXaleY2DINqsWTyWXZS
V/xH6RJ2A5nXylKzJHKniXdyCRQFa6ib/AboaxbPYFUh2ZUlRx6ciUL8kIKKPx4VsP/zsyWp/knH
MDne471P6MdXU6tacgodAkK3JDykcnffypLC1GOBlDsqTD3b1uKFas3r7ov+rdBzjc9g8gTH9N9r
6OCIXQ8y7QO3H7sk7ZF8k9CxjYmTK9EokCrXfT2eKPKsgov/QSTSCdEf2qOjgtNhw38hTNqXErw6
6naYCfkwN6rdF56q5oQsWIKbU5sVqZA1fQIw+gBXWp6NnTNLt9VVB4vLlmkuNK3k9Nj+P+uymYu3
hHh0Grvi9xQEfxuTI/c67mZw72rTQkVNG4B3qHIE4kpLQxwpwqB84CuDUa4UOHxlBHEGsvQ96H51
fyWIzc4iMkyOyTaUz+eVMFaO1TgktjTtZqc6PD0f7zhxmEfpN0yYGZSPYshKeHSlMjXTqJTR6i64
m/ELCW0GbWUkoR0vVkEUfDPXYMZWxHWh20gN1GjtNaK2rbIL9RSdaiPpQn0npp+VUrnq+mERniKm
XGcaZCZQ8R6AfzalMe9KgvZifycYt9WWX0sjdX1QLXTIkRW1w86U//5i0g6R+oUvw2/2ihxZu5eW
vrpwSiG/Eud1T9iKj/TEJGHBnkNdcG2V6+L83ySpZD6CwrwNSmiXX7ycNOdu5bV5qP8x2s2+4dfx
UpxpYMg4b8Np1jXIVPxaZouAoKFWZ4h8mKB8GmsjXpHNXXplOe1nkOL9jI2j0BLF68zXeDyPA26a
DX42qO+xoBxE15OYRTgqodYJJsYVIcu9f85D7MM2YmHXTvxBwHVNCw9Tir/z8RAXrhQ9lreQ3TFm
7tbdabjl7Q/tnmthImm4cSumA7qqptbBY5CahMDgYmKQrPS3iL0QKYkR9kGpX218888gvhSNybPy
5FVuMK3P5Pwc1/z34LriP+iC3LCqrhFEj2oTeUQGfK59PVITrZodhoCUs605AAReDjE6+FDzWqgD
Xy3id8B05afs2gOlqsRPBFYd5c/tMqPfq7Q323wnivVttJWAWpXL7XReo2oExWPbSSqHaFxS7RBL
yTDOSJh5SGjcJ9k1/Qhu8rgAfMbFqwHWdgY9eFL2rsKq0xeN3iGUJiCRaHZh5/emEvPhGE5u7+MQ
TEKNaNymHckjRXpxaSmjthOPICFiNOKIe9NUjXJnX3IXmdvI3L/dtsFt0VGvqubj5NhL5DlebgUl
9cbH7tcxThkgjBtnj3SI8Jf7OSt2eDFuzDDY/+vQNvjsUf730ciZ4iQU2D74r7ZC7qvUpVEP4R2h
7u5TkFsmk+Bf5QhxeCXwUgQgzYeXpeUXdKr088Zq1HcHE9zunmxbrmC4KFoqCc/MWa+/+YSE49zX
dxUPhDIzc2L0gSM2EyguAY+0bufr55VW1x3RsoHuyVPPeXLU82HZX5fE2LZPNsYqc/Q739bq64Um
pY32Ydr3AgMJsAaNOl5+5Vmf29BYSgWeSMP4Z4b1aobiWklC2GGNxl7Cod+eaqpllNG+EKenP/mO
FxZCAkL+hIpg1adyah0PgVBYkJEPugNTLEXNiLUDpamSrFd4+qHanliF3qOgX6z/Ep3XOt0TSlsa
TEIJxEJd192TAzTm+6PNpeo76w29dCAjRCr3o6+CQpiRi8RhwT/f3KAOL7vRDljKjReg34UYyxHD
9RxCBMtU/zksX8y6Iqebmf0vt1QQbM0Hnuh8PAuS3N9R0z7c+KHj5G1TU3eUx1vurCX35MbJr6HM
+UlwUhzV74W404fYi6gx5L9W/84iyba8xKEShCdThQgZh4UmCqm1UGkUT1x4dphIYP1rRSGYCb0q
HpTPUV4nIAvP4G24k4o1oUJWxsqX3CXUobDT/n5TAo50in+HuUsVhdYN/Ze5Vef14Vpd1qNPnGRp
vywGXRsEioC0ZmAVe6PHYP0qR1Kwazkg/ucvh+oZ8YdRGoOvtRmJxDCaX/1FEjtKqHAX+DWo1h6a
fKE+5XYhS3n/X4rS6q8lgAJnBkSz27kxE9/Xa/e1G3txsJSma4m1IOhTRF+undPQIYtVAqi2jU9P
XQrhqC6eFsf4D5eEmJKJextLg6TkxLJ6GwEpPNkFS/lZOkRMZqGEgQhK/HgP9GfqekCmx4shYTT8
9Rk60KYZbi7V5yDmhVGnfTM4vLehMS7UPZOMnSZe8RCtLTBiqbv8i1b8ElAEtnfPalGYgU1dQzis
Rm5NnuWz9MFJWGVoftRbIlwcHdFMCKvI2vjOcJ/cfbwAKI4A8laN9JMR3LQENqgtzFRMfIU5ZFQW
8DZJQdJVSY0g+Gyb69RrUuiI9ObhcYX0RHwuAEYbAWVZp+RVmglN/4eWQhAkEOoXJaz74sB9y0Ly
nsB/EoN3dPZCWZBebI/6DjCpyzuHCB7O9LOAC1RU56f1spFuawdrC/L3LHROXBDQGfcAvnra1aK6
tuViLE0erxaMxqghbpA7Eb/8QMHp7HoQ4SkU1aCfGEO2z6L1ATqQbsc3Pvimzi3pa+4MMbYG+PUX
BIm1XwqdR/HRhEw3xSF/3G/hIb7ke94Q32nrW0s4NfTVk2K7EcGrI5wHluu16K18YAF7V8jxyxY1
PzOkzOiUj6c+rRLLZpRppZrBjMDa4q9A9fJdWveqWwLos0Kwh5jUoyE0c4tIO611N+msl/dsoB5P
h3kgl9r9oV6MYLENvQ/fhNBt/ADv5R7CNbRzue8jhyxT9Y6tkphbu1i248hJjG4UVXKiXOBQ6WSQ
xZ+lEkMQaE2qCHC9A+UMbNcAB0Kg79qKDZRAMrQmNBRaX+Jjt2YzePBiV8yvsW4wg8V8Mic8OzFt
3hjIqrE8VvbJASMuzwaZxi9LCfa8PTK6FmlDmfnt6V9CCavDjaD/OVD3YbVI29wABndtwV10eJEQ
KiLWqNkrajtiaxJNTK8Pd6cUZY1/kcuW3EIEglWghDsElyvW7Nqr4Apt98d0PWK7m+jDfAegF+mz
73YuY5VhmgMnKv+oLNagqsLozpirkjHLJcG4piMECXnQGAau4ou5rog7Guxq/Tt3RNhCSHJEB9HL
yPgR6hkLBrxODQpgwYd7P8kUz6u4QJppqYohAXPWDMe71JK6vXAvoX395Z/h8LPJR9+PEKQqPRek
0obNgYzi9qmnCSuJlXxNTABjFrI2IVIJPzWkQI1mtDg8uNScmR6Vav1zDgElwcImmFhqQa8z3jBY
fAVOt1vcPox/mio12d127Ggh9E90TWFp6Ls22DStq1e2q4lkUHidAn+4Eg8032zYHJ9NBvV7FRsq
H0CyyvU/QLHJRNpZFnbhK6RQf7M3oeebPBwMV4iHv5P519N2SlcxztkE2DeC/CMFPVC20j27Ipra
xIQUIJNgXDbDq7QiYRUcqH6Z8QWXJbJ4a6ByrEM1dEc4G38gOxz1TboFeudmPwU6o5FfcL9h2c7H
BqQ6HkdPHvElMVB4RH2eD9LHH6D7Rw9l1King2f6TbvLHQ89Spf/9cvrRqXs9T2KS+bSr9IBrh1h
zxYGxxEL4s6uz/HCQHOsfjZnBPcp0fg/XmvbHR7CBixIqdloFwshEUzmprORtqRkHIqisqN/E2nR
yb53zzWebJf/SMOLs5smJsfOajhLQYWM0ssfqzFc9mB+XRfHr65X9h4Mx+pIxW0zvsFj8ZHuBe01
XewobYSIi3L0carC8KFFlGQUnjLHGwj5eAFhIMtS6gKTlFrxpPG9gyfWgQ2Mkk/CDS1EV8cgUn7w
BhtyGb+v2tPqcwirCWGDYxiiCUN3G6tongYbukP9bw6WJRoS/he2lDjqK6nOMuuIWtB63fFsQQ1c
B4CW5z/B3a49cyqVMLm8RpZNiAgLL5w2MAfPCHQeBmaHq3u273dh2jsBi7j+MhCfQmHkb7oDjj2O
ZGsObjHQ2u0Yz0+2laEq1jXwsRfqTg+b7Kfk7beXE3cu7uOHLT3Fv273S62XQmU22AHjN4i108bD
1Yc7zKKYn6h/fLX99F5GAhhX667Ry7ixPf1fNooHpiSThIxdfuRAashr/i53vNWpJm3a4+PxrTeO
1N1yVsDcMUq2YGeod5adUjn/ID2uyNJpzcxzBeUFF84uJtuymfo4QM9gkYqILnhYKpbS9f9SVMXV
Cev4831Ij94/9aOQXeYXj0te5yHm98/32wCxu1I8Mas0zPA+uXKckpNTVJDAPBmCu/aeawGI6LFE
6NQdb4ERtt3GOs47rV3ejij8JiWXVrNP6biR5ldEFspCyANXrinbI4uoOtuX82UXq5wEPd0V/wQS
BYo7fS0De0fvYCRD89XZr5e8KrGQ5smaWvJ91h1/zkObqmHOT3+Dn+wkhTER9vL/BY8WkpOyrUcG
qNuPjxJcWXuDzJAU2CatW7boz7vjRiZ1a4DX/lUN0K56T/OKjzruKEZEVBhCWTauc02PINVEo8pL
eCeVKSSfsZGOOz9bJ7Bl5xfbGo6q9Jebqa2sS5k48dNyBKfv1sb7pKozOEKk71D/7y9U2drsNUmk
5+BVwPiO5tusgfuZ/RQ7z3kyK+r5WwG6d8AJy8dN4SiY7Zsa1chnMtvjo3WxzKx4GDN6laQrqNEY
knjBkLpas6Yk/9EWhJRk0F7MBmIMiswD5X5ApyvgLJ72hRWRN1KdxHC8Utzrr65PPfrw2ie1d6Hf
KvbdpKcGRMyMP10TT5HfWM8uXOwFC1mPW4Y4sYl++94V1RUT9s5nyDkIJOJ6ztm9QOY2MJwJzacl
BLiY+RsUELmm7XbT+0uaityTi/AV8Xp1raYWfmATN8sCS5WP1CvofwczHtCSyp2eZHf3XNoORlBu
F3uOFf0HB9lfbMdDPqMnG+RzwMxMsNG8jx6mTa7Dz0ycrxJo9ld3pxq/kOdppHn0uhETbl+Xz/b/
R+lVJctUok2uPRJV44FtVbuL1W4Is2U1AAL41U6rcYUI4CChP0L6jHicb/YKDgKvs700DoGrz8O0
FRvvlXJTkEMJP3Dnv9ppzpWLpMgHhwDTGvnBGAtAaYQYfeIaBd1LdCMvcHqbgq33BoVVscacWdtn
Hf731FNLiO6Uo5lo4hh6U5ie0P/LDI669JKSkX+fFNujAlWxhQSeLvZH1gW6Mm8ntUD/9M8PaG7Q
gvd9XnPGuC7wTx8pCzelvJ6xxzlW/4y1F6Uw3WMVGX8vrPikn3QuLLr2sjshrktnC+eJ2mQjs8Zv
pIlp0s2VrON3OpMdF0juzu7fhtBZoo/ABwQa8+l3rqEInWaovic0VoHOpvlAVr5V3uKsjdkqbtMj
33MYoWr7d6jiqDkZvPlsP550WoCKtvTZKTQer+cDnV1lSIcGesXVnpQ5m3fBg/KycnuauzN1OOjg
Mjag2z9dosEWH3Gcrnamin3OBlHy5JpqpjD/sWtCD6xAx1Vfb6uHol5V8aIqtCR2LB4i2ceWJfeP
Ke+mtFVCwEo5+WqcjRuYSpHQk19rKIZX8+7E82U4zJ1H7QIIM128+7z9zaUVSZIvmtzP0kRpq5Th
zPZRZ8zcclrG8YHjEhW5GRwxZHduO9TbbE50gCohrq/5zdWhfCi/frSPnr6kne1YcWu54tMEakjZ
UVG482qM8WctouB6pVFGrz2sn/VwjqZ9Wty0UbjnjyyTrjtznNnFYFxLdnbPbCKiUFOYuEnQq1kA
Ix0h5KLGUXD1zZVzn95pTij9WvBUs3riHgsaqFFGm32dBRMKAycmGN9eJ7nadVTxaeacXEabns0A
rD0qmJyW2cricdns3oENRdiI+3EECXYTF6Diag543RPLIk6XXjol2deE1E1CiZ/Mp4CzpakzLvcC
ezjJiUF1t7VF7eh9myl2HpR+b0itz59UJusE2QzXZJRuTUlo3KsoyE6hDw7tiOmynMWKDAHnuLKz
xONvBDJPGBtqTfR3S7j6mmggMrld/YiKzstfkoj/c1RIKFi9uRhNKqOholiMbK/VNgNhMY5qSF/S
zBMuQwgtf8rz1+tun8MWEpAzWudys/dWby41O+7YsyPAxID6QaNtZkXZJUiC3dK4wYp9LGHLi7Sv
anev7sP/dortSIPqwpvFG0SOn7zeJbXG2hwfzjgiGLceaVYH9f39dmFpjqal0V3todwv6vIZJaZl
kfDNfQKfLOGyks9XPeI6HvfENVDs7XpiVrEHm9iUzMsZd52BXG2Xp5MZlchET4hj0ddzm35HDREM
6DZvgMf8myWPcbxbwHgpj3j96HiFpVoTd7lNKlKtIgUZKspfxLr43J8qSQ559fg9dyI/x9G7LxLz
fWdkyvikXHWlzVuRNvKBSK6LiULwJc31WTY4hncZvUaEuqP76zToVsrSLDZO1R1iI0YFUA2OMyjH
02qxhEj4VE598GGta9mDVZJ4QVqSl+h98fcTH/MWheUmYvxOU4xlyyY/X24xqiSCu8x3zbK9OVfK
SjmGh/CpQAOa7VDTD1z0zI7TOsS0T/JYrGf/UUjzQ9T1CvI7YPTVvJYog94kTfUrDMCWksOd2IGH
MNux510dqSTv2bUr1JU8YmL/KpsOpLiUuHvlyiMsOYzVOnOUTvEg8Lr3XqgfNnhKqrZP5fkmSzZ1
fYKRWFb7Mnux66HzNh9PR5jOH5TVXIMem7tAlSVqdEG8uJgfNpt8/gE/X16/KiqwepTtrGMOr+a+
7hDqzpH/VvZewm1SlqycitwtW+BA/PhRDYF4XSljCmFpbmmYrJv+yHTyNWIq2Z2soye7sxTguNAQ
kfnHqccRywkHMEhFJdb5QXBVagBTKG2xt9dfTtkIL9Z9s63YmgAPNEf9di6oDl/XTMv5jJjhTmu5
sp2uxwmHE0AgvrMWTCwJzjEDtDGWw5nzSXvFHYX0jVI4AAPhbEmyyiIs1fMbTwTM7Xf78qUMzMUY
TvcbUzVLBblMKIhMck+vUt1E75YfvqD+6iO1lMzOaRCzvjGUoSVN5BB2spK6GUgXb3VCh0goUdj9
fU+P5f2+8evyMnRZB7xQ3UZkxpyRut4Pj7D02Ll+Cg5Rc1wvPSkmHRJ4m7QVPZt1OeU6rYc4gDZO
kca0hnXAnV99F8uRzLP+ch4VtFXIFAJ5OM5i9bhpNfo8W+Fa7mZm/ppnUI7ZcqAD4+m4YHX9aSGN
ncHcPSLqsnRtyKtPbF/qT07fjr0KHMLFedUTA3U817wKIE0Gdx/RtWLt/R+wM3DjwPflotsNsyqJ
NueZFpPvbPskOria8IvAhOoOwqqZ1qcbEJmYI2wzOjjrHnKRTVwEZTDxAxd8Z3jXr7ZvIWAuWBJc
E17HaEqhLmGnMdrEQoMAr1NGp/VKf8jXlLEP8j0umVqxuf/fCIKaYFgUpCYWkNmpIJzdAg22YBTP
wM9+PCJ6xPlkXfUSmIgONu8z7Ha/yE9MkAXsfoyVdIfMSC1RAWEIa5d604UhDKuOkz+ZSq/hpySp
Mj53BAvho6Wwpiy50w14mIsmu/mbhBv0qKx3UPTUyRne0bSmgFZwx6e3tyCxW0rYpZsXi32Y4Cbl
1i78mMLG4CmBXEIPfzqy4MwF0cagdyzLHhuqz6IL+F3nPSQJjfgf+/ArqgyhXxep37WyTAXlvj2y
u9xBUCfK3HTKdwg7xvYKa6g/IRe5JjNlKr4aB2o3ruuxKwwARBJsL0G5u/y1kFZfjERdJCPbdRP+
muDDInwrgyCjBFIF03GkE5pkKFEBrnWurYGJXZul6iDpL8Um77DxolPswYyWJdC2a02wKnGrY21J
/LAYvZF9hgOZ5frcNNz4bNdZwkC4saKkw8P+1EZihHR7XMOG8fPVam4Yr7zMXuAa/hzHXld7fGxE
P+T4t6o1JjyVJNVhjHtVV30OlfTwRhW9cKgk33nFyy8X/6fAk4bby/cK9OA+Fjg9l9opOCC9nex9
+AOzD3xwBaY44R6UgE+8uTBQbRU4DSZwS/D4SqBZIM6vsp6pe0krWXDvbM8I946Kxzt91QsrJ8Ib
0K6Dcmgj2vhYZlCkI3IN9vTudmVHft5UlFilz2gWJC912qq+y4QU7X/D+kFJcwsHb6q1ZGADM8pt
UbBBjZhRoMBzb7qUNxNqnFgkW198vOmuC4lmrtpS/m2PzNQLn8MNIKIXFIXbVCQW5C380TRsKZ3D
W2TBugtlvkp1EzkPh7itWKrC7I5VA8rPJngiW5I4pJj7nQmkmKGFcRCOttHWm2yavLiioPIogZfi
QtRYw/n/xlf7GpLk8wpxL+ntpWBFn7g/t/AF65nu6VfyxMmucgLU1XQpn7ZqnniHWmQxTSPUXr44
6mL0sa41Nhx7M/Ag3PlDnyj+zOuvIDeKWptp1xiTjdYqEvQeyQF29fwFZynyMWBP1tQO7Q74b8IX
dEWk46tOkjw0/wxnBqCOHEHIz85Zf9wGz5L2fFZFAZVbK2M6djLfpWKO4NmNVO4asF5z6lXPd+rm
caS9c2nPjIIk71T5fhVLZdkoqMxPuhWtD6yA3aYmdgSBhH3kQWpHVLZH4OPRYWsjzE35FtATf4py
6YgYF7Ot5sqEc6OGz/vUE3jzKZ5DMVk35dk3hvlH29LvKV+tC6QuEcdn5T3xI0UFYBVJggY0G71o
762Xy9CmRSxP7W0q3bw3o3xvC5BXdTX1+RT0fvnxzgUfhLUSQdwK9ljF4XfuQzsTCRiYyAqvA0pS
vNuWt7SEw1HpB3/9+A+UHY0bW5/kjxYviHiJMCBvss5UNpO/Q/kFNx9aD0GAiiYRv7jueFTqRZuA
s81UpsRZWr7t+Ou1Fe2T/w91DN4/1Sunqhzhh8t++THUBR7xqypzPJ1UI+hT/fB6xLyzRb7dak0O
8FqPqZpc/lPw0zfa4wsO+Zp7mgLA85DqK3Q+N996xwwa0h4GbCcpMZ8cpGp73BKsT9yf0ktgDwzM
JkfK2t2+DhCvG/57J9lkmnXf/PJDs8g5FinMOzaJ+IadlOZhmeaYwcnoGkBVoLpAoAQ+loJAeTxL
owJbEkb1YqOnx9s1dZ2w65SlnxNYqoemtFcwTnKApk65Ljfz1cZuIR022jNKci6z2WZmSddW731P
PLd2fdsd5y1ywYztYdLhFsrhMFn3vFSA1VIhTdNqDuUyIXws/x3Y8bPMtJpoZdx2LUFXqENDvS8N
5hjPHygsqBlx1nJczr1RljhhlDGhs2b1JJLI85+tdWrjelDqJduMyQf//0ap+Qs4Y+ZfMmVIzzoH
aRcP13wXalyCtXOogQlAr6ZWfof5C1pBI0eUtDwaNY2BgJ/d4Oawg2ofB6FSyubjcNH8UQqqNKdA
eqw2W8jKtncRZJaLS4BR3Lh8CZD3rfkeX8P4pJj6rIJ2UTS+i9Dbn1k1IEN9ZUJJUq27vekCHN3e
a8hnsN040+jrWigmdZPzdoZvCM5gaiwn/AkJ41fAtyNL51Au4VG94GWE6eCNDbzs7e0Bv0exVcBq
6aoc6S6/IUxDQ1VCa3RumdqWCs4FoxzlP/rFBUz0p3zIIW7XyHKcAtE5iYLaqxvuUhl55fryTGKS
+Q3XJ1egDm0Vs18PzEUeB02F4AQ5HyEFtibaMbVlhKrQXIoXfmrPmQxd1Zm6gD7Z//crvLq1KAuR
fIKOg+g4rgueE1ihawuDB07RreDd9C9+RvgVrzc+JC5BhXFQrrpolnBULaUiwIW4Ztqb/9G/LQ0o
CC41OSdYIiCWxBGT5iy2mGLIrCP2Vrio/sVjDDlcWkGEkArjUQe8jpuhcZeZC0IramMn/sKBg95F
MFVXdM3YL/tY5doFoVex2s1xTolRWs7cIDHkKr8tE816ONpd+g2Z/gFYqMeZNLziO7yIUaIL+MHE
8Io+7CFkMTegzSp6yo/UO4KdsSbtZon9NW8XiqDnhaw/hC9OPB7w8oYGKC/8ta6sQgcu0ckgxbcg
GAHBK8x6LGpUhXUlbX1S/7HZzMqzxyimiqkzJMBHLplVo2SKXoH9ZNhJ52SyZZ9IfwK8CoCb7IlF
1jdAjjr38wC+qUcRTM3mvVHwmR9AEiRE/kZe45+GmdEnGAKTvNXZef9KMp6ULsPkEMihh0inr0I9
IkoVput9H4v18koA8pTjQRVkXLe/njATxxWzc0NeUTPXLs2m8qMRNpZR0nK1+fUOnjqbfLd1k4N6
Hh2kBS6h9aei2H6YuSTjz+v4f68CjghTwTAn4/awGwkLwh/VCSrrhbkLPwmYC9yvppTkJ55D+lnd
02jYTtt9OycC3i04s8HRv30Sdk2q/fXZYar248hNAn/4JZGxaNO6jQ/tyYpQ3Uqk0MvovBW2v+7v
RLaCR3o5oKe9K0hQmEwaYT91khMyl0yYOO4ysIOdaX5F+0/bNzcWVIEhHdbVshLLJ55Ek0GbNY96
8Egygz5LYKs+L9JrFbGtl1lVn+p1M+7OE0aAXfQzLhg8a52yu5jbZj56FcCsI8PFrn/MhGsEgwsU
8bUYB/x1XjZNgf6413FQ/57KuNlXn/J0J66p+HWUWa1uApurSgOlr9PkvlAbSEYOu9Q4L0AgrSVy
xmSEnQxa74SHpq6aYpA+0xcnz7BPYNGLTcgBFXnwysp7EIskgfHA1zyAcEDMGMtZlxuWhwJKKTIy
H/sqUNcFZBlHo6QwTyx1wbnxqnsNn5Sgqee7iTiif7Aca8DgfoHM0PO6IqNebfx7GxhAvJ3oPuDv
4Be4DcOZl60WUZtgSbi7NTZ12vmSPgwK9AyG0gxE0nT2BqZcUsyl9YVl7BCXYD2h/T2mrRZkAxH9
TLflyqfkRGtUXFVDITFAA3lGqs+91f+evErUHa1N95sDyqF5AC/SGk8MYDMgD8UPJAy9gF2065sX
Bzb2d/5eNy5jhZUxmlcEvpUsQno+aLMdu/Pu+8XQQK4r39kA9VSEP7SOL7FBaF+L6D12cVZw5KBg
XRX0E8LBh0f6h/ialufF33xzLyRYj9/1SJ7rnyymIXJmo/I+k8SVhJdZ6Co0Dep5faXgbuf5r6Rt
RclU4ErGROyjmKsoBc6OoVjfenHYL1COpLWVQvj8RkC9NcxaW05pn3lZgYBBbtpifAi6pry0CnkE
Y+xaHGPgRxFfTCCXFW4D8akf+CG5R1vZWNccHC/dJqP1Qb2RxyRCeGBi2HRFEdpHttkZ/WFtyiJM
WG0JzYIIMDErrwuCIXE/mFB+OgAUIO7atTSGhYlLXlsXNB4P556Dq1rA4SAHRKw+/Iu5hjI+cuKg
FKmS0vo4+tIy+R17ny62P39onpTrouB1up1lQ2QU19s2ZMr9fLcnSPiR8ApNLKGRHjJVnxqij70E
Nr3iZSPzI/XZp3RFOot6cadF8JW59BxAVQqN2h2+qa9TlXuuowVItraYWP8Dgg88GIEXKKjAJAhj
mHq120jmKFqOTyIRYjYUGuqKJrhFJ9/ohpZ7X2FmBszbDOOvJ+npriuoqJzsAMk8KF3jpajOqLCR
ljjJJwGqV+Yac+hVAYQNNH7s5MxdzojjvusUi3i1z3CsQh8sm2jKg1UQd8pKJXpKM+VlblORwUUR
gYtxcI1CJdVasUsMhzJZj/nxCB2XId3mrOITox0YJbMT4DW1Lmo9VouhmMetlJahZ5XLDxEIGZF+
rGaiiE6YWm6vcwHwlDmskHpOaL/1cyCZtitPrtNy8uxitTouduXdOxkQYG21+4DLUs8Hk9nB6qcG
gOK8etRFy3rzqdCUg9wnHaTkhoDpBhVyqiw7jwBh0yk4Z1NAYvUOBuQ3ZnqIINC6U4Ahgm0HK4Mm
bK+SAxmKoFy774dCNoScMk2oah92qaHEg0fLXq0dWEqt64gMi5OH6SdUIz1+UElmVog6vCR2mFpD
oIFyhhsF3WnVKlL3OYlIPCBOjacDld7Ero3zLGrFkX8eDY48elKb25wpU7jHoNVvFtRsfMo+/ghi
COvaLfKYKNS5+0hvlD7skfvXMjcrhIrXiIoTDRLf9tn0gdo5z9U6buCJIv8zqxH/0jtFadTUsWIt
63yeBa3saYVGrXeav3PcNgEhL9F7lHDWrVqfhKfyo/4uiEQ7Ofxsh5oYd//3ixuNc12z0ub0W18F
ruBdu28wU1ajXRYW4wYDlt0rRAszJ83nyXjBiPcNecl3PhI3xKu/5imYaWJlEI6ZxA01QmToGXU9
P7AQlZAoz3dNKB8MtEKpW8lMv+MwDNpSzJkxPslUoLPUp46Wo38clVNCmp3m2TuEEBIm/3pkCoyM
0YS6cwcVIctN/3m8dd47EEIzea8w7oHW7FC+v375XGeXm6ZIEAJr1l5C/+YrWCKepRVQez98Vq9V
XKgrS0Ot0myuhxhuO2xxtCbWnyIMl9CdCX+EnYH0mSEXdiUTYLB2kqsx5rYT69BfZx9aX6zLLsj6
JwZOxmDw49oAlJEguZpGDhaOp8Dm6qjiOVlqHIldQqiZxMYt+qCtEvSHhYZ4ESCsvTTsZyUYil5f
NBQfdRnIBl7J3eYrF1MW6r3eH5kZKM4/6y67VYHuH6hBv28A8VMmyLlgDa7bdw1BnV0Wbzjz7Fvx
XkGs9nSK0UaQ1ZqYj25V7KRuxExQhqqxPfAeQ0pTSJ9qPf90HCH4FHb5NhBrEsIh+bMMoYpOXKac
8nA5dHVk3lB4/BEWWHmocpavFvvTUyIkkqmhmprIAmy42FsDZe/Ym0JMr2vGQVEhpJXUk8XC/WlT
A0eg2JAUieBkA0EXxXBwdZtHBEa1KI8Sts3ilsaHTKWJ4ECsktrq+lyCaD/sgTFQKZuO4QV0EIpq
951a097QE8RGaolbvL1EPV7cjMh8kElz5Ci346j9soSUAPbwGc3eplkZFMMj/jBkX73OPP4UX0F8
eUoC4ydwkIESlzPS84rpyRoWNA/BYAgcJDOO07K6fvJhdycBm1ze1qfrySwQVuDNJoGZdWpUfGVQ
QkFFMqpAGfwnXLW+Ha0ETZyEIrmD6tFRCb3Czdoh+yQXrGTq1hp3khYhhdN46y/PCc4kkHM6EjZI
ayMyGxdi1Wzq4B9brpSfNRpa48AbiKZWZw+y1EqbBmlLgsfv2xfJlLj//txUm/jaTL848rla3kT4
KstFsphkMbDlSpTkNNOaA7GHYnru0St0v+PMBbaSPGkZhD5kiSzV5GjMCqP/gQUx8VRKbqZDBVkF
XniXzsa10Un2WhKvPyMXksxMUEWWcIjrb/xqbh1q8ayhne/ZozeUPa6Av+X9oa2N9iUjQOL84/1E
p+UZKXfRFsOtlpyr0u9ftM1wvUnrJ94XwnKis1zJbTQdiEhGi65jhaEy2NL96AfWyAQ6f72SphT/
ZKL35ajyrbqU3YyVtoUM72EwstyTY0hzKbAUk7wN3bN/SZVw9CHvhSOASJAID8joWf8wl93nNGmQ
gZTVqWYnfFolrbhn2p+dp+UdmEBeKlsjfMkBTYt4wuspi1p4d+X0xm2eiyU9/wibmBN1q8XT8rZ5
w752Q4cd9LAsbEM/rHtbu1Q/6pmb7dWv1MBuXCn7gFGrWKu1ORsl3PpWNuWWZzbjQ3w/MAsyIlSu
KxmAodsjE2p26XqtF65ptMow0EEz2Nle2B5UYNpaJ72VLAoI1HyKDP8qqt66PxOCgTsDas3S9GP5
fokJVWrTc0UMq3R9FwV510dhXqhsMnrFKr8iOuIaYNtfJNQs1D+UesbTViOdtFUW8KySEelzyT7a
3Zf8szFL17Gy5LUJg5vkgEplEmwbbTz5e9Bx86vC/9ck8iChmN/WoiuiEjMqdCsXG4ekZahDAE5R
OBxwB7MNMr6FYuD/hoZ76KzaB88Oe1WHpYLTJNYxJ9ol31e0w7kyb1l6YDVNKJoKHAzyQu3JGCKf
rR4CpvUjttY1bPg0G650NQpCHWwjLVm7Q0phVBSE9zYSWe5/m4lI8vt8hbTO1eKzw7JcMjwbNpRZ
R9BkNXMc+WSAhivt2aonJEQUFXfAyezXKan7EK9LvpD0xblLf2jnJhJTI5feXWUHbN5nKvBz5vO2
p26zTSgXftvH6//nHvIO0Es7wAvh2to6FoFT8HTICzP8U6KGrXoeyWpOb3xhEFvH9pA6fgG0hmVd
IRrTyKK+esqTvvzIx3S5tUVC+VickUMqCGDN08eqJxthNHRVmd6cnsXh1va5Bc/EFXh5K1L5wZrs
Z4c3cICvQ3+mU650rnRNVhRa9afTRGAKQtNGFdOsLBVQN3K4pE1wh6fntN9mSBDpy1Sl8TN23MDx
ALmkDF+1Nx26jpp5vQQgZpgdM46gkUQmU9o9jjcz30Ujqb41lnB6/np4bR8S3zrDkhgyr0wSVO0k
JPQLGj7mi3hy25P2bn1QFXqQpdIOcPzSGKJwyAMfepwzKxh3Q3z0TTigek4A+mao4EDQdfzRYn+P
4C4SdEqhF55/nwMYQ/IOtfFN6BolMRI89fDrK4eu6gzKJlvUDN6qScYIe72+cTdcdae1ePGg7JrL
TMOnmWi6UFNBTWySXPoIFLVOTVRuAZJx4kQT4VS0rrmXPbRFNQaALmtgU/7pMATl/uNysxmRWfXm
ifPeSW1lrAHKW2FLeiIWuYb8rgTT5DeUXVpQmfRbm7qOdd3XbLFUEYXTyowshiNmFt58lRNEPlhf
tONo48I9HCfPtEt2cKvrx0ZBT7txK50o+CLooyjIqrOgsGKLVh1r8ho0FIX6c7VKQuEXtCVbxgOi
HoJf5OIwzyxi0rGzDbDvd4T+WCb2O431lH0+3kdhBoSFejbX5/hLCKNlJTcoWI9Fd4bagkLJtYMS
N+Z3x1e5mgwGKz9s1Xx+e09b9JPWOM5SXTWOM5VBTRiFVwigqSPG4ON6D6dUk5tPh+tRSDrjlSUL
F8h5GKdhXwbN+p/fOoegzvhqapznF8/H5AddrLVoas8xaG4RZUz7pg49c4a6V/uboqPEbP3TFsSF
8/4n74hFVHUEr1Avj1Vc6qNnxxDOXUhALOSVkHvdNrFBOpJfRPCDjF5Vbhhdepz3f/YqrZk2JFVQ
LEkLdzV9o95gg6z+d+Yv3V/Nmdl8iuQBYMAhAPMD0QFJ3uSR4AIHxL1Pi7EPbYgt3WVGDSiYzgos
O8oOb7jAHhafNVV86Y6yHVGzqogJUlaqpIycMyGavH3cWU6wMQkP/RLO3ag95WwzhbYRtiXOouli
wkew1N0aq/oEPCt3RS4EvEg8AOzzCCw4k2w+5h634qyiQxtky9X/G523zlQXDidkf6pUiWZn1mOZ
nNtLZPNsoyOqC/+6JpWTuP9DzuqFB+vSaP6GPXyv82LIJ24Vvs5UavPjEznOqGofNWRVJtgu54t0
MWsJUsEsXA4SfIpdJrtd7B9gQFuoNua/zorFKVyZXwxAyFcmbk+1Te6LZcXe04GjfN4c9EsagaXM
ObF9xHXEImvFc8h1uAf3EkolpGLcVmt2eJJKdh6hh5zZV2W253Hi5z/jeMayo7lmxs00ZuFHRWIB
fM1VXG6Ho6p3DZrI+xLTyyVoIIFL2n+urHnYisLthxJoZ+hnT7IeSrN+SJlUn3sY8p9qbxBIi6Hq
q1cUmQZ05TaiEEAPRV82TECU8gmNLisSQdELYQs0HiniMxYpLRGNebnfrjd48nL8T1R0iK5VpkfA
di/dgSyoJlNU6/F5IzJykcbLcTL9xbGg2cRdnAQ4YMu9XH4IaB7RsZVGNGcnOsKHmjFDSG/1UjWq
yslQnhf+UrmO8sIUIfsOKE0M5qlATxD9J5Wz3yZwBpjlYte07rhv3CPXbBW+dNae8GjvZRohW8A8
vXv+d37kRHnxvdOS+ir409OBA2c334b9IzzEePsSx4Kg2DsBumLFaVVrCcRVj2BOZCImCbNtFmQG
34zSMSgIW80InEn9MDmtktWo/s7HV8sNNHd6ITAgpEdAbGezKV+kMGlgIF0KHE472ugq2ptR48y4
hjLQElz7I2Usyt0Y2cV0kDGQAxITf0VdgdwdMh+7ZVP2JF+HjfweX7GtgmAWaswx721Tb3HJFkQX
DNE32mDuyzIgv3rRCEdTi0Lul6xr+wJmD3g0Sm43nJ8LhRd0E41H5QppHGLKsce6uITAphhnV8FG
jeOzegA7y/p2xXTgngzcFzjlq/vr+FCgaVoehyvYMzO/yfRM6gJ8Ta0H4nuOouCYlBYaoZSe5pA6
2R3IIcglbSzwna3yiNfph6/Q1A6yj4v358j0nZlrss3Db46tEqAUl2wXoG5EIrQA4sb4/9ROAe+2
NA8eSZxKQU9LegPdF1EpG48DMu2PQ3Eb+ekgVI9G9cYPky8KRVlHnKwhRR32a2emSMac4JWEVS7p
Jco7uyvEe3aQn342ZJM4T5ZnUktjLM7vY1+M1r7vLg91ReEi+h1uAIMkdXnw3hPrvm24JTlvRFQe
pWMKbKlS8nYqzvrTFv+MxYRnZkOG4Thg9bNF1XCB/1pbD3sjUYlJlt01W4hTplh8y8p5xEFiaO+Q
9W4FVZnvTyjieAKa6qeTrgOK4txo6CO+SC8jpGcTUxhXKA+115wU5fKBVLlCYQKD+UGhR9kFlqFW
6tKnDfex8ybUDu0s8iVjS9dko3qlwbM9Qo3AWIyUsP3Xk7yG+y8osWor796ScZ89nB+sm+ApdOG2
2sy8MrsGi6UjCa787Io3hJIX67HWj3RErkuqlOcFpl5cUxGGz/AfMITgpNbT0oI+n5wSHfOPCJ52
SEJ/af0VEPmMrDq07cmVbOCXMpBB1gjsP8Z2lFYXA4jPCSwjUOl/WU0SJRWw7snKlxwBRnk3KShE
/ytwRMX9u8e2AuIDYnpf3rzV3EDEy/kMcgYM5wGhpna6uXOpSzZOY8jcw/i5c1fO3TCvvLlPWnQH
eLQH5pynV7j0SLEfglbD78ehPU/s0FF3BO2KuXvAIgE6Ez++QFWNJYRmTZe+c1NIrzw9PC3J1jC3
+9Y9xGoBdlTzYWkOAStoRV+dJzSb3/PAj5Cs4vqDS72DfLMlJeme0QQgN5s8Ze7YdFW/3GPQDrO4
wtyrNYFbI0FMO2re95ikKK/9UHryZJu3YGlrh2SZ4//ZmKXrzIfrIrAeOPVSivziSbMptQSSAuay
iMXNZ62RcAwPpy31lHhRpcTmATow/ZlIjARveHdNLodVVTh4C3e7nQRW7wdsrkcyuPy764o5ml5h
6omJpP0R0UpGybSERUbLA8AyzOAjIpu2RR2evAOG+D0ZJMFHUNwgna1ShWITxjjCg667/xJUjP2H
eq1dRUG+rQPc7y3ObDLLpUmv5IEVhXd9WxIrLndkPEk+DsBQbm2rvOU03DxwH9+DlSwmtZPgryu9
iQnqDuem8OnjTr8MIAszMJGwU9sVjV7QKHhlSYh8vMQsRnj1rWrEpuVyc9S2oWWfydgYA3qYuyyG
Szo+Wmi4K4gUnUSzMAcl0DF2r6Uo8XWwfKkV9caCUa0aQEqar3DH4fnP+lq5T2PqF78XoKqUintu
sVO70pjAR3W3RoZHEfwf2suXRElMC4M84+RiqWXUGBtboZ7C5gqPxM7eRtK60ZuoHJsPfLjaDLmK
6+fvdc9Rq5Pj0QzFp7W63ZqKFbxgFiBNCtBjgN8tZRB0tMUhSBiNCZEj3lC8W+ZYGedqkrsx1on4
1sm0SXWay/nfHIRo+U7SFi1o6nnD3f5VEbx0FlEyJmMioAXuxDTIar3B8n5KOx2JS/aSYernB0+w
npu56W7lG97okHtzyrZO8Thc0ZaUDsIuowWMvjfHsiSw9/57Hm/LAs60yLf2nSBxC9rI8LkP5fKi
7f2X4+E68RINU3nrECDDDGC756yd3Dj+52DeQ6w3ZYbEAlJUwYCe597EbpvTsrMyDtitJB+lDV0h
OXJIX7UX6R2otX/pC+M6EseGoDMEIJ5wiIaC7JXXjTrfzYeyFidbfdJBHLMsrpCwaAZB8sk7fCfP
/HWhpAQx2kfo2AI/7Kttzw1Dk9Lt1fRGk0vOH+FawaMIQnq1oL5cl57ldIR9TzqEWTPW2v6EiNU1
frrxQzHbUsnFBgjWWNDpDHzwmwBmVvyIdhZD0rL/7rztnJXw0XMcdTBUf5/18146JUBvX+l3nTda
5lt7swqrO638HCOmOPedNBEwSXaTvEKoDHKzDVZvmvjRoIfGnMzGS4eu3Vewd//pmNO5WWf/KK5y
ZsSWMAIes8HVCPPBgMNwZDWDZmkZfXSsuOuybEB5xQaujQlSlJn02Q8+bHExknO0NNW7tqUNWrHC
+JHwfEpJxAzYf3Q4DdSjukxH6VfkbZlvIKRtos4My29Ct13ajk1vSSvb7s+PLi15bqqm4Icmm29+
ObB9zJsi+FV0f5cLSa+k4jRmtTQ8XCpp8HWqgmUYs/nhvkcyw0xb4BR1/eknApKA4X+tN69KNWAa
9NQyKzBcXn9xGYSvbT0+ISs/wCV/YACOXo0fT9Uhtul1tZpcxUjeDYiomrIFwhzjn/EB6523ILPK
cROnSVEFnmJSq0EUbVr3FDtRoz7J3aFrobXc4t6N/kqi96GcjmK7ZWQy0EI+XW2jecOz+nvE5JwO
Q8M7A3CNEy8XyUjWZ04j/pXiYwPhycqSPQ3gUk4q9nTLqlyv94yOnVfh0c4a54j+oeyP2gYWBqyH
fPXiyEccH8KtHn8Hp1jS0Gcx8AB2UBPSTcOvnQFQ2sVvOefSg3kwAUAr1oqJOZRmBZfP1wMbYR36
YKFmBYr62zlGIUY/Muf4j1lyt0Z5rsIc6lxQNvIF2lAFNRXOt2JAkvrLqVpV3+XKRrgmdHkS1luC
hNod4/XkElJWh8cMKlQPE/YFUwlSThD7srIeYneJxymkucTQedZxXHuLTfkDA32CHwwzkXh+nRD1
CGWxSYtMf7X4iCEcrZHa7td79PQLvRSc/ccWsJRY5CCvUUTAU+//ji9OXzcJBw/vmZCjAd2a6pEO
OF2phbzg3SNef+MGPoysFE5ZqzkSqZ3xxyBrfNyoP3pF4ISvhhjUcrxk4qADXcmxTk+HUp0Zi/2V
h3lptzazHhLxT0g047wvfAhG5o0tOdum9zskFgnQvM3lQ7x/w3HGiXGCsBAGPm5W8Zgp8BGE/W9k
3tUCD1hf/0sFzGTJ6sowf/XY9SE+SdgN2BU6aDFDWSibGzxKChJd/15C3OsnKVExAi6s+KW4XF+I
QqPMKaD9vUGPykYzE79VOxlIg9XWj46YxrJ3vuV8FMtlrG45joZ1ZcYdTgXsLJzKT6o1Zjt3tQbz
b5XZ95CbqQ4ipamed5k1FsENlmnLBgcY61E0u/oGnelKBvk3zgCrkr2DmaEtv0YQF/upeG+ythJ9
Tmle5ylXOoGXJ349XDnPn0xrAn8MivI/loUCjmt6uuC5t9L6yQmR4BThl9j6I++5G8SIwD480mgu
9LRJRsfqUHUKNKlazk0Qar2m8FuCfhwAgkQ3/6Zwzu0dvoJ9oKr3XBFvgw2kN9/E49z0WzSJ8JVb
W+hCKhlUWkE5kJb1NOD1sQDh+qAN0s0TVNYf7GrOiMqU7rHzEa2hihU2ax5/sqaI3Jth20cBvDiW
GAsyUX0wqb5n/qPx/JBtK4SpEkx6pG+Z7HO4VwukBbxyomM3f+xXmL2u2ObaUinFnexpVxk4C7xz
kapj61Tu7zTuLg8sAz7jK2iJApAracONnYFNotxVBniAD8qBgI+u8i5p5iooEHE/8E6J0wD1oxwp
KE5MM/2a6/Op42XU6CnJoxYjHipqnT4HtRWQzf8j1CXDnFSpWGgsE3jswXdKqNJ+Uc5RR7NqjTVb
gDT6zFbhuX8Em6hE3gIkh3YDEvK8cvPLn8Vi3egMJtne3NFzwV0oq/xezz+/dUUvvYjDOGoUeDLW
qd7Aj8vCNjGxeaizHAsmWDWO82h/Ag+KqkKT13ntPTlf0k1BBbPiavUJS38hQO3AygUfq3hXt+Vy
XaRj3t+xwzm9KbA2oo7hxjEQP4Kj8ADMyTt4aDf3YeClCZI/DHHkFWXj8smRFq+T5ksuCYtKLhoA
DI89DrezwKYlNL0f4pjuSrnCN0HuLMYmCDPpzUe9Ga9SMa26AEnUM37AhjLAPKPBRrb3kBnCPRdd
dQzqAVDu9XBlEw+2I+B1sRiwPhV2tCLf4yyF3UF4MsEpP5994n4UhrU5nc4Bty62Cnzbi8ghoQRO
t0DSmaJxkcVClKUIrOTB4EBylNWKTkrtqrscE7t7MWhX1LS908c9C/M/8Kh+4cCIhqfupk/9uzb1
f1HhJMAvT7N9SwnjxzgCYoPKcNmuTlOLlBid+MtL+mk/kYWipVup80yjljcaa6nxndGVbjOIz+Te
nA8gDWlFzMjWA8IcYFwJ3GF7CmpjPG+e2tgnz3g1bIZgco0ROf8JQzvztIXGJR/ux9a+74rqaRVs
qOq3L0SAUt+4kehZiQa2j/JCQ1j/gD88ccIV9FDcCizm/PzakYccys+N0w5yVKNO4DVGTGarWX0e
Iseyip8vPBINrqMc18gtRmZJHKDkVwbGqBMlbKaNc2JBLJ8rDTIT1Xn+Bh2HdiK9QbRZknH9NhSK
yEHq7RY2G0dNpWmc4LdIVJOWpC7HnNgrjnJgMxy8WRV3hlKlTLCQ7BwwY47ai/iV711q5wzymq1V
/u/Yo9kAzWDSNwB1BILHvH8AiyiRQGWUAWuEaAcya4J1PoiLH2/fSsqtgPsDFw/PaworWwZ/GBJ+
jjQBJ3lL6xtQ9q4RLALYNAJrqH4lUMxixdpF2a5r0aSBK9hiTzrjIBFedqgnlvmSijCipSLpYmC2
vjon1TeTcUWcuxDoD6qNgxcxjWw2wRgNoP1RH29W97mPK5Y6TV4xPL4H8ITAX1cFezOQh3qEKEzW
vb93oBDD7SVHExdqIUTJDiTuWCp+vfwV5Gv4H7QkxVZzv/bdiKkoIkuQFvnp45KF4F/5eQcgaKZV
/2HFGj18i9dj3/VMr4xnYuTj0mOiimQMeMFp42eUsZuoUmvlTfgH5rIxmB7Neh89braYe3pYwtMk
KX7rsxIIjysKxZYBKo//FdW13iPmm16ESsjv2kolxlZtMZcbo+flvpVFkkOVzcrlk4PinBUDQSyJ
wZksGk8ePbCx+UtFdP1ks67mi3yXMTzeWCOw9Ftl+vJKEV8+yolqJHzJWZSq4wsBm0BwQ3F8Z3yt
cStB8tdXWNwzb76tlzlz9vgDp0P6RFYq7z6gaZie70GVS0UEka+bMxh4P7km4OLDpVZWPtnK/qR3
F9cJDKoa/HwGB3YfmLZ+cTOM5dmxu9CNVCDiqzp3ZjKYO2WQFKlgUfh9JWT8etdh6E0ShKUlnJBN
b9PDn4ebozXE5j/XSGTu2xi+WE4WpfBwdflHiknbMqI7Co5bIqX78TTxrupGVhu7I4wQsOm8kf7f
i11nESbjoP5LcOiOVNHTJnUMPczvw8aULHdRgPHAmrGmhwysig3s9usM8KhbZm47c9RhmCJBA+hE
jAyOlt/fNiYGo8VQKFecz6TyP7f0BlSEhyB+WnqHI2Yp0hKLTlDGixXdZdJkLZqUNO7wOGO9f9Jy
WVjsxWu5JNPLGcrQ1bMHVe/v8B5Wex2d4fNLPereL/s3XEaxg1NgQxIoMckvxi+R5aLopzWV7SIS
yEbDaqm1qo8+iYsFSbqaiMz0Rb+JK+CKMJiguwhOadDUu84eQEj8g0BdOtvpIciO+vRn2n/jpwDz
/npBxlIQvuuntRqA8QI0oX6nBbmKGOjsvLZ1OuOS+UdjRtgBzMHGNBXjVKS3nJlXBh1JdQm1H+8e
TLhvf7QwsI3eWcArAL9zxZouLNAq/+/4fXCx5q3C+sULFahvdcvGiYi9b8ylpTHDDHM6qy9OjVKc
YpugpM+OJNWgqt+qHCSoU4MQa5YXloc2d8CiZpiOls9aXzLq0F8aVN469WeNNxTALooIbdOxwAgm
V/dKhbXSXW1W9G3rLd7NpIw9YPYrL8gUuPCNw6I4hrvOwJfH4LA0Ap1b4DJiAQBCvHEcJcNH+cCF
A5yy0t8OkC5QZgR7ChQSuthKl/9MFvq2Nk5ZHZfaIx8femOEyqMkjOT1CbyiwbH1hl2XPquBqrxL
TWwY4QZw0ITSp+F4sWUMr24ktlECvs6hupDWbqMtN80S8gs99QslMqMY+dPuHn840kxzXst4169J
z74ykRlxoeer1H0hrR9HEzh+xYVKjvXNJsaCBOtOulPpk0xjwN7uNopDQPGlnJZzysvwCnzpt8+o
+s8pHKe4s81mHehduNLOLLtM4d6kG5dYFtVbhe93CN/siqxXCMomk6flRRUATpa6cf+j1K/W78yp
Nf0sP0YFGTk0LdZ0M9M+wn7QBtq23Pv0fS9kvXhRl/9I6rIZWnJDPFMuF3LR1mpy1/tXmeOBATpa
CX4agUvgHphy0xueryDz6JpHaUw89Hi/Shn3ABuKXJDJlivT+el2ayMq6GPhKbMKRiUfW+XSOWJt
rUQd192aqQQFqM8s18hp+iDh6g2ybOLX2g3KogU9i6G9iw6MhHG6aY4S/CohnMVishZl0tsWF6qQ
k0pL+IojIwFSkmazYxLcoVjSVisOTDJlfsZS2pDkNN2L74j45PCbF/LcXrDCd5LEJqbY0/Avu2X3
EB3kQ7pGVsO9VBkj9M5Q3ry0SYCVNbR2/79uJRfK5fU0aRDHNdGxb2H8aoLkb1w68lje7Hx+AvNf
dZAQ2Ef7BeQmzxgURmESEUEi+vawhCqgpUyyxBcQ9Ij6z2iEyZozYbsYvN2/1rsNgDgw8X99JXlb
aptlPvit6um2ELw1QPN+PhY/pgsNMMiZzbxT/aCou+YeeymveL13n3DQb930nh8u2H/KDnPJH5KB
73RUXxUSkxHXgzKL4c+IwiKj2elJhfcReKq/PgEK6wrtojT9R6EE1Ny+afdzn7O/UpMPLLrITFBA
IMYswQsK4n4ABqHMCYVRRefM7X4ewbrgpbAHor9L5s6BAgo2BfzB64KaRhweR6yiDJNWLRM+wZTJ
aLxEZZ+wyoEac1eJObvFrbf7VwVDpbhXeSrSeOtePefTc4A7vnB7lnlSdRKM6maL6fqH2jXkDnGf
pq99Zzq8gmfXYfEQzl8akYnEOXkfqZInJzzGTOiioEYNR9AWjvk4QzagABQq5smbr8TrnHPeP6wb
/F0v/gwL+KjhQKcqtFMz6zftCiE6CYGYqhbeI1bv3wtmTWjVwqN0eq4SEvrl8DwjgaVE/fRNzVyp
0OT/cMOJ8fhIDpWV0FvE/JqV0i71Ek0yJ9HMc0XwcTcAaP2tX2366ZeYq5yR4Mtjb9G9xkZwmQc3
27gYXvYmyp1k0WAHQ3lWfZyfqywJF/BE3LTzkfsORn7Aq4Kk37iBv+MiSX3oYshc6Q0NjcuHgY+6
99d0jLLmpUWI4XVroxgMgLMcpn9BNQEfb04OvG2lRrARQdEsqgW7OzQ1g9/eLmEuXSyIddmSCVqZ
Ny85VWm21BVxQbBMS4F217XF0uaJuZ6Y1Mc/AjL100epw8h7fxdWVIOEuIXdmXO3jWIiUr0PQzX5
y67daewnfc3QDnM8+wgaqIqZUoBOjxbCo03jaJTVfCv0tS4y69ErEh/u1ZtWcQXUH0mOCdRwuM5s
55Oi+ZRF6Ktqqb3N1a5uzsTie9VuFVeMI/L8ntVfJ/uLyrtjIknekDhg/Fb6MTblj9y5A/+tEPaE
xtjGWSo+sgdZW6Ehv2cEd44e93XyYyx+x9fS6fOm1w2ZofnRPjD+BnJa5uscabNRdGLC+1c6GUEw
QSoEPd1Ki4L6ZUUlsHcM7M4daWmR93/kQj9y3sktFBxE9oHnQgYl+/AN3an0cIpB2UNTXaXFnNbg
G0IHlaNzkr1hyalYXniSkTAkYu+JdVnE3zVMbuiV7BtSHjPkKY9hTw+c92xNI35VwbaMA1Vw+b7K
zrx4V+kJcqimkJk3r7Q0gtpZX2RUKdOpr7U1ORQtdMi1n0NNIk/n4o1RYQwDHKYmIYn13f9QDj9u
VME5ShRImMFT5/xXgfVR6oTOSE9p6j/rhLAD+kUNMkflCHeu2Cb+RvcNIY9afJzFHFzMlqvxjb/4
Lx6lFHrR4yMUEtkzcZEJnxvTmel2ao4CjcRco5xuatLHkA9/BR2+HR2ttvM6nD94JPRUDs7cLGHR
SfACC3oKvs0JlHpr+MUrRFtw62fr1FLayl9kkTkqIftXZ/U1fJASvT9aVJd0K4nANesj2/KfUMtg
jb6p6gS8GYrJC0mLBX9ZFsMSDreSVThULbH+sr5VJ116V9PXZtdoDSPkBVFUHVrynpSNOFQNRqy/
rxs+cIUW8ltyNG7Iad1G3IpsXfYwkun1CT63xbWOKkHfvkjx+hsfrY/1shE2Jfbv2deKKoY2KVnx
BTDT5WxlPO6pg9D/sNkTv0E0x4DFBiaaJRuCvEmX728yPEoR0EYO54ihLK3cdiv+kMi143XWyZo1
BMLVBLH3w0kParQXV+3LnrUaoKq+ZI7LEwWg/aGQ4zvPw2aPzVx5Hfxq1go90KU+nj/OQtHWmEz0
ZpgQ6vVa2ldbXMoQULepaEIMCyJ6U2U9yzBaHJfdrpwjyWqsqJFN++IqphlDBwasbXupANxUiU4W
khFhu3/XI7Ui8v/3jWTN1K/aQQT3qDMcW/KbvTDqxfP+46ErCSHSEh/qM1sHHGTkYvVSk6e+CeHf
j4XkoaAmbvOsyoCbr6I8lHBoFoq9h67exGbjUWXc2gWh6q9kXE7mhljZ0FQW4TcxkCFfRDZKi1Uq
Hf3MgHU0iYX72JSDts0lj7WIY/18bjG9lyHIWW5XNJ87BaT5HHAUfN65ZZwjdWjNvphpB688nVMp
M45gtMSDOVVUlanZuX29aROEq6Xl5y93EqE8c7f8R/cMvzY/XxAuEZcl+m4ns0u9ewRqlf517EKK
2styMKusLbAbLVcyBxCOJlcbCHr9X00tWqGURDW5VjgNE/9Ptk2jtf9aNpFU/rYmnK4AA0h/H+s7
8+N7hM303hsiYpuM7/fW7eRzoRM7RfmaH0elLjMEULSkZ8CKzyY1hEMj7SLrGum6UiWOLqxz/vhL
arQ5OGkO9C0ysQON5WXuT25tEz6UuWUpk/FqDprEyhRlT10ANZ4ZqXkvXiy50VJLbBqQ+6lHcdZQ
9AdgmnbLla1bXGHYQj+nFWHgTqg8g03RVkaO9PMD48kNH2K4bFQc51ZUCw5Xc6K+pViqpaNZ9oNJ
3FR69IoVYVL/lX8D3+qgfF7+tpfPxlPc57H6fGIBCsTzy9dCj2Wg2myN8CKUyYD9YN8J9uihnkCN
qKXVgkCTEb/UnHSEfBfwo8LkPeHl6b4U+L1Yq/vmX7fFb7FvAv6EV9/l79xKcCizYE3v/geCIfh1
EcmR5LvQ6nkgxJtbNUfL87WEWPsKmcmHWIrknBGEZBfc2rfIYvjo7KCI9ttY62QgAxa+2Z4PP9ZC
b4a5I5TniBx2cRKMJU9kW257obZmIxvuOrnNJowDM9W8M1MT79ugofprT/stL8mkdC53oE2IUNuX
YD33Dxf9Sz6rBMYC/OlWMGZMcZ1U4HeflyBTjyLcRkuo3hwcyAzHtRq/4RokoCt2KU90x9ng91QN
goGKqExa58xF00R0+SLtrNDV67Iuy/eeE42QT1+z72iovl0d9/WCi+Ooa45yl9sml4BOwVB4pnTa
UWV9ud/Ge2n2Tk/uRm/arY3F55vdT89lR1SnIpGniices45in0b2+mEIlfXrfLFgJK6TbG7FSBvJ
jNMuBrkq/6QSKzQ+TbUuQ2UOnAqgt/LxOooRp3eezGfNJ4IIVIN8N5CbGDPKD63AfaL/E/znJ5V/
dJ4x6l9CVEPkgtET9D5sIMzz5PzZT0N/my2MvXo4/XS5CrAn/lCnibh1E7C4xKHofUecVY1V09vV
x+ICF/cZNyGLJfM7G+kaHJI9G28JMTCHmv4MtSWip5TAhp9qNMiF9Vyl+E4GGuShzMpRGeEArDBa
57c34X4O7ifgo1IjhYyH00GosOm3NC/a/TXF2fyDijGMGnmEg7ax1hT3i6Vr0BsgBagSJHa4I9J/
3z8Ne+l55UKbq6cfziBWAFxugGYpSja1p+ggLlwKlNqIhdVS2SyvfX8UoiADEj5aKLW/OtpfBLhy
1Y58ok0zeVtfClQWVZidc4GZfVZuSZIGZMthaOatYI23rp2J16Rv6wGufpAvuBx2/Z0iKVktP5LV
IxlPgXu+6o8kt6FoXi4voZhdQW9IKWZwr30nkoXvHxrNSc/b05oXi3Z+g9mBRBnbrkzKJzMw5fF1
kSgfg/BziZWF/q7qb6Ao2QtgZ+KSSc74OEdbF8rECKt33vKboibTdMz1WrfnmIJ+QMnnuC84wB8O
00E0SmwRLRtj6iSPDmMH+F/faKuXwQVo9fD/32LfSRP1Q4JNuQKkrXZdBOxQuI3fRgqMeZ+vXAgd
xh41Wgrt0sYxqxYRIqs9PbSz68R9Phd221IaQ5mEbcJuoktwrMV8eX8tYC7j87IKqUXq1og49WJO
uvVQ8z8C39ukfYxovTkts5mnABfnelFKimG1e/aGVh1nFi93ITQlLFZMeisSMrjxwAJMcnIwDso7
Id4kDLKImbvRCKMLxsf1+1oM8reeN/oz4KGfTH500KgTR45Bw9vUKPy86N9VDL5bg+/fa/HE3u4F
kSPJrVPZyE7ubfbIUBtCsWSy9jmPtKqdZB1X80/b6KiJEjsrEBuD9SCkYcnkANSy+82E74ICtO9R
HRqJ5qrQvdGVckiBISRlyiHKdB5V9g621FCIgJB+4sCmk/B+ofU/mHtaCAVIh8PeicOO/yqzpz15
2sBNr1olclr0dHmQ/LAtXIm9kLDpZda1C6KmwPkZN1UAeXfOoJ6R0hzScq3Wv60VvcO2N3DZkC1r
rhTTdjnVsCqsDAEmCwczdGcAVYmzqruzeFv5SI6nPQl7wPftQx1yKoS0RehrHbv05WJuTzo9lHzG
1hj2BReknIw2EXxX/c7LLlf54wfCsBWf7E2NknIjN4k577M8lWnDuHf0MU1Bs/1hLCgDMhhTtrAy
rWDSGblWuGdZQbniucgsH0hUIHM22u2tf1plt6iOntUdS58X5srGuMShQ0RuQvL8WXuPJN3QcL3b
1PI/pJ75asag3YzsafbQdB8pGdsO6V+MG7YRiv2S5EFCfi9NHpKzA4rZMUvg8qhOld5EtM7mnETt
35y9WN5ECztt8/O3H8nbJKTnyCq7Tmqf1nUs117eePn/TtjF5cSbl5x0GgswD8B65wa5/I3tkor0
OInoRTBkHfmBL+ZM90dtuWXMfXOsWgfKhY/y/8n09JJH5UGrYZNZoxwYohY+Dnwn74SrT2P1ptsQ
VpHuCB8rhkynPSA77gAthEW5xzaqamrt+cCj+bWgE9UowlXXZeGRmQAMrpPaorRXQmqmEb6gMebk
gTrhrNeQ+zfUMkSjklNpb+s4UHrm66TdW7goqDoniIzJRtKNdtG2S8/MWAHfPORcIqsA90wSxZVo
vDrFqzqNNGQaGsN84WtFDQzvwSgawIMU4QX4+4BylMljhg3isDTGcFSF3Mee3jxrqmUXwlA1pbvT
taXyeMwtnoIutRRnzt8lmRTACUffPpjSg4i/XJP0rsFpNQ2IZY526Q0cDxzoZS8XhUhSF0v0wASe
IPwFYfhJCHsYNaszB6Qw031WwX1f74fX0lNBf/HLL2YO622SdHZ4zGcJlT4u8Zp7KbPJluDeY00L
R0hacm9YEQS3kGInfbk/psEgU53Zkea44cY0Oh2kUnmZKwYfzHplwSqpFdpknSQtjMtGjq1VU1Xa
95gjfZaf33jtRhccd5qPJ2MdQ4+0PfNLLS447jme0ZyTPxsOxzFMPEMj2ijbdGs0Ims0MbYecjMg
2n1bVtSFkdqTxzsp3qyTehdI6urcJ+RWU5sioH7Ccf/fsg3VsNqyD2Ad7brVhJCT7oA2k4oruSSD
svcQXnaDAFA05ZsPxhOpUKLINXSqAJpFKbhXfz3ML+5fwpGAdzeQHnFXH4uIzSvaZureyCHjjcql
jiOi0Yec229Mt7wxZ9spXRSHF623XlHLGEygknGfixRSC/2Hc51CXnnV4uT9sLU0/8+PCuX3mPRr
MG7OWIRXJKa2mV1jfbcfPDRE+PKWg4Jz/X0rxf7VsmJyw2brZAongPnOcUelsSNhsBgA7JdTbc5e
g+gqGY/UmI/v8DL7Ohr8PweC8DEFBmV0conYK+XbtDIEDUsPkVPw9iBTeeacBwqIjOuN4TZXB+rp
9sARBBkEIrBJ0xB2UABYbqk3tq1zXa0lAmvdWkEmxQrXSHp9fP20BdsTrR1C9LSdy5XqIgq9PsXZ
r1b8qLUklWMLnfScsIkdjkXmhZYnyAt2N4Pde0cx6KlNLE4F7xGGEGvZ01OmqUHjPhj/K4TgxsDs
hVa70JwvAUjUkSsqJWpLTEn0VopeioHCSg/ECpp2hdNFTOlpqyhGRPmCMoKMPwi+mfmAD8hNr9YO
KmC4oBe/ckIMBGvBd9r5p1sGon1xkkwJtXjR30hf4yzSYH97LGtziF2yjToaKzildEYTskfYG3N3
08QpHCcHjF7r4KFFoXk8f4hBRKpow5GqGYXHuUTEiuqEtROzo7xwhBQ/L3asIo/U1UYt1OfhD12g
Mt3NMLAaPp/0k8YkrFsMm2Ymb//isVwFaAxYSK4IInTcpXl8fFFTyB3OucmKh7NQJDrjKDlpEE4l
EHGWFl68UVi3NMCmaIvtPJ+TiOH0Oz6J5wPU6D7Yc+yp5FcKQT4ZN3yW7KmYheWVULNU0I+BkBs6
w1LXMwS50dlADP+lHfgFA+lVkEGZLbsosx3J5xMqYDaHfZMVAfEuI/Ma6N0VcgDER8PEYZ3MOhTn
PyLa7j2lWN4hNRuEVDpwdO7ywj8BjcxMQF4qh7kmENXsSA5/ChlHvtU2ZFA4ARNMa8M2mWBTiMez
/Lp85UWrvqujHd9YtniWW+rLlbwz6l9V6kSk/SZvi//KNYoXGFRXdcn90acc8mOdSxGw2Zc04/Vs
xOXNnNbIVDF/OoZed3SkcfMhehAkua/82MGBdhKDSqJQ0ZkWyqCASeDCa7hpmFjZUXFqutL9DNjp
q8lyJaXk7MPdLU90ZTSaXEHfC/C7bz8bBJwm2Od8+75E1QPWG2BRqVcLp/W+a1gCLlf7D8qdMpUN
PJrFv+OeDdc+qDfIlmGXV1fQ0niroOfDqjJ5Va+C2EYdqH0hy2Ng9HxjGqD3dnvEu/H7WQrsRcr4
oxsIeHRgqNSmNGR99zpmvxFypvJPRCjJtrWy4WZJwMMDoxOhUi/jXJnX79QoBsAn0pLJo70YgLEF
Q+QRJYge/dGTeoyCnJRjcaGNHv4XSQss3bHoHHnXTThfoDuhXmaSfKKgS43iHkXvS3FNoN9vPhoY
bFwcjnU/nTulHfdeDWNNqx3SGMQfBArwvOixO0sHmBmaIJ5wXTQrixUmYW5crlUaBzf3zAGASuWn
JlMbbC1+u2WIKj/iUBOt94G97Uv5j32fowsoexTpebmV4rNGzusM2Mf0nsg9imp20OXcKl/LVrcU
NufAMFbeWnfGLlKIPmk/hHiXDNJe7Nshajhzq6BOkFX37atx/9RdKO0gjkBKqvTHYDfWi4d8NqPN
xxGbiwlhM2jmgAE72dT1Vm6k56rJn0CNzKF6grHDS/kigCZMwjWdWGgclCbWShbtuuK5Dpd6DYtD
U0KI9lu3s5OmI6zVvVLslHcK27In4Tik72d7/USCcOGPbd8AXzAwAl7z43NNhCQxzni9JWeyl1dt
yba32w6agvvfFI0onWG79Z9yiRVpPrTY/dJB1jYvagYWAmW664BY3/7MyzGJdGsLa612WsPO7J5o
KsB6VFqVeFLxV6wg/sDs0M/6hWp7BalSTZ8QvVZIpR+JNvr3XUAfW7eZqKoCELYt2VjTRy4W3qfQ
Qpcm+GOhORssP4xybxTBnuT7qKFT0yT/i3apT1BC8m7qtyb6MplqEiwJKozvlk2GBZqZgs8atNqT
J4a7gHWzr4scgTnqdrAS8dOCcosVTU1iU3ZVJqThVU5F+eODrHInB4+Hy/u1kNcaamDw4VNpNirW
6v1ceEQCLrk0y0E34mhkYKFiFaSnoE2f4mqc9UpN28mAy+WVW4Y6SMmCuHEZaMdO+Ofp9ExG7XJN
tyKualohO540QRMnUr2TLv19rlNbx/U5ws9jwew45qlIbeSd/3xcMUcagoj0AFOFhNtp2EID6lqg
bbAXCrEi/05PJR0F3WEAwMf9rdFpS/r8IMKfl4hIo/6n8qLt06iwATRat5ZMSMINyl2g0elIobKc
pvAJE01QDVSxAYh2AaK5N7MjKZHXr79zi3Ajo4OFWUiHkJxkUAWXLJNas1iBf2bCYUii/Ax9LqJA
JUSD+NY7K4hHXXslvM/3soo5eHz3+BLvfKskIBwmYXxcqm5Y4KFmU9SGpNR9fmdoedelpktVjsdY
mSGyeMDvWhVnvWi+BpjadTZvfKo7/RV/geVa++0nN0M425QeYql0SlPA1YebW55umwVNacREjMMk
EQiTZakW1ubd+YoAHqi6g5vof2CuhAFExJ1K5KJBtRfK947DJY8cEdvJQKZpeN/MWMNzEnWPP9H7
yfoYpl+/L3UhX/LPLm9eL2pMjAJREOZIdrvVfvQYW+Q5GAN1iUOSPisisTGTM9cDgoGUjQzuuSak
1srWI3XrqboUl9+UWOZHdVyCwTFaYOuLxj5NuQ7YZaxTwSWlPyKqH5GYHBIJTf4nplW/YFPmcKPm
jvOUKMODmtvUNytAlwZtOtp4uC03YjdA0s31JBRgYkyvciq1CqJyR0c7XTtwP6YvRM2vngYX0Esn
hhNLLGotUD6UtzGYzEc5arR4Rzmqp7E0hYCnLBGp32dxHmWDo+iBHrzsOQhKwgaqucp7lavdYbKM
sN4gS1cWLpVtFMfgWbLCv/Ocw7+b9t6+W+ILU7JO1OoflA7+UZVpkKLmv0nP0FQ2UuORNmiTyOY3
AGiM1/h8uRUDaB3wF7uqTfqpUl1elcC985WOiV0R3Rey7navbJqHgykObjSlrimmalmIz5K8fKIj
hOmxkiZzzjW9QzUYLdtKBlqFKQa55oy1CYA76DsrKek3KTurm0XTka/8X2je/Rw5oghPChOzj9mg
PU1L0regMBeKkfZry/oV+tw9YOz6sxRcBstLEzh+Z1LAtIAAEF7xSdITtxPh0ZD27Jk4wSZFYUB2
dYaGbN3Y+X3/dE9eJhicF+7nXBj2A7fi3vLvJt47UnL4JR1u2bkQlL2m8MKRiYfBVQ44OJ43DqkZ
uBY494Ry3HMttqzw11VioPZQqk/eABEGDAWHXUven+xxtOmOvJvgSZ6zJuYpt4/4Yv+7ClaFCDj0
ogRjrCQ3y63NbDGks0hOaerIAoP75lbjo1MppYyL4lwBktkwziHfhKBbBy9HTa8pErWhBVho35mR
M54jEmsuQn4RPNkrVMAXIv+v7sqS1peOlM2vRVwMu1rw2RVIb/EUZxwl5XonqpTYvP/HndQKNRy8
KYlJP/14qr8Yacc0ruWO4+nqDXBpk033suKIEfMcw3uaK1gRFaM4LhL6Cbru9ND1CfvCC15dG/P5
ygEHPXD3XetiBvoogjnPz4tMr+/X0EPBbvf8wn9mArDEYijp4uAijGWKhk92eJ4R6YSLl6EDnjSY
+aEJ3iPilJ3SJLGgteX99WNhUKM6HCLwXTYHCEVNv+9Yu2ygXYG2FwhW4UyL8fIBbn8dWjXpaaAZ
RSofrUQ+VuvozWys8ywV01oAs8dbmneCPbaScxYzlUSGBcz87R0dE/PxZzCLNS18n/DIRxX3C+oK
pHoa0VQwirKCC74n5ghff891TAZH0GhTHWhe+w5MOXbc67w6d+o4cURfRDnl0XCtDvZJBJBe4xMI
4xMs2APOb5m3vj+R5Yy4MtyMTHzQgR1gUeBX5j9A7dCL3O+U+z7ku772JpWMv2Szw/+15RYRdtm/
rkEA4sbagbFznDQWPXI0d1Wd2ETLdNGsVVhseV1UcLgkLztpuOdvFvHmuuoOHPEPbrY7A2ZP8F3I
j04P7Jd5htNQB8cvYNJHF6ZRpHGL0UGADyxGtu9p9NkY4UA46rN08n4V0zrtxCcPx7hXjllnsK1x
1SSqRfQlCYkwdHefioOkJEbrFw9RxsSeM1+9xShamfoeFzSr5k2QazACiXmqYlZDcAGdV/cE5xNx
HI6v6eiEEcbJrTIfr4NlqYTa+ugQGaIOrY/GP+eH74483HdpZVMckU4PEiHoJDz6sIIBcRo31d9v
JEBfioPgFy4qkcmFvhB2ofDY+fiHq1GclUaMHKLVrCmiOkIel7G1wygdpr8yXpe0Vo1GKsUITgL8
hPKgwTo4XYg9Nh//QjKpS+2MYj4TGbRs3NWSP3GzTyEqX84+3i1x8ade8rPR4NOw1ZkV/cKZBMej
yDIq2K6riv+oAGWMsB2hPVQLZrUAm5Mke/iZLkCzhVaGiXy2S6TmRW2VSSYNoaE654eTWjAFSjrK
PCjRk/IA5XsxWxGIBYD6b1evh6ZCsqTOEw3MVoD1iaNbKXyqMXKRIzcH30z44NL0q3InB+YgPiOW
Y35lKXpUq6W02NNpcCLLk+Ng9VJfAwvQ9W/LhFc8byktB1z5iXsemrmsiEOiGzIrPSIMyRbxxVSw
/21xQeJfHHPQTNoBRiH65AggZE/E5ZDByyskQEgs/mPqU8n3DWS7lvuTmOy0ozhkbXR0BiUKjz/+
7q7Jucz4Mpni5884cu7ZhZTzfP3O5w2KqiHpprOp1SfLW3O2wYTLoAfUfBWRkBXEjLfrTVav9v+A
s9ie28shSxuMr4Vca0qzMeqrEZV9Ekzc4xwsaKPv4mfbfxCQ6eTZyUbikNAss8cQmT3rwjOCAxot
pV2ej+BR2oE8X21iDLC426Q+503+i21Ve/TfZMOqSHh/VFeQewiinjy/MNeRUYpo4QXFxsavEOJT
EZG1Iu9YWewlNWr8s4cE47QiDMKi5/X9oYH9ndd1INXVhmfpTTfkPdhqArCUKl3NJB29DMH1VJcJ
XPxF2TwMTsM3rg3o1pBl71/Sj6S2Guwly1YB+7r8Vb80VrHg7Yrk+3u78MYn+10US4eCNrhLFwJz
ia1nXifjOchh+gjPlzJH2yKAbMGR4cWrIH7xvY9/riI7ovnLG0MZy/y/wuqnl7ccSKuzn4+bX1KN
pLTt40igQx5ArJ+7cY1JTwS0lSVbC1mAaVHaIzsKtGH17DQwPNsq5ln3DYUAveQoNZu1yO/tTe+7
fDy+esTB+JUegWCd4aewbp1hdvbn+ID1fgUSwB2HlH2yUCx/wu05DpBK7MwV9dXODittz+cebzN9
4OAZ9n1wF/GLSsqSEhU9DyJwe/c5ZtJBO8plPGb7OLwZlABevTAQUH2lUQogzgj4rW1c+1HB1olI
UxlncX5dl9mMxt39BAO1LQfC/rU6yb1lTXoQNWC8x8aD4gZ6XsL2HxI9F+M+MhI1UHwUkM4OuiKG
nUAWFMXNZi6onbWUVZTYTHN41CdqqwnapNk0E0hjRWXsfRjJZ6NEUqgItvYxYAW+QZIKr7ZuG93I
NFyaNqk3iJzJY5WPsx0weO2qZi6PiYZeVGLAwTlDlzTA1mOqlIqa40QfJe+M5ry65aDxUHjlRfgd
mQ6DoCWXufr4LLILoaEtvGcn4YAn4UR6cHTwWwhVqfHcaR5ZAqiZ1ZX8ooo8/JzbzKNS+KvMINlA
pjYOzu7Nv+C2HTVJYViZ4+jooa0aE2jVAxFdlwnjJTw2rm0BukF/y6SABnJ6AAswAnSjKDfPfO7B
7pOStfV3Gz7vKcyqDCs8ZPoAy7kPL2mBtEcGTlBo6bUSNsyrrYeHF0tj4AIz+Uoj2s+5PWWeyDKN
x6G0qBj0UnQtPo5qZbiLfK1B2m/d5n0nVX61K4u7Zka9qLUJO8Z46fyqmYGkpA00MlI2nrO5Q50/
bDO5YaPZVoYk5j8QC9oVEZ/vtBAnz2ReRi80XHyTTn85CiPB29XAeIsASc6K22JA/Bkc7L10xKOJ
w1njJGghubkrU7EMv7zIVQrR5rnNLGMGEWtMLZSfnquFS0oUIQd6RsMb9bspUA8FTmZ+D1iL50Sb
0/vo4Z8bHjv6MKOa49PdOfT4hr3EbizuxLKf0pV98XnZLqN4WjTIxhmpHVA6uPeBZ8NQYESvhcZo
ld2KITQ1JjcgUHpT0zqeIdo3IuqdoytgWz2GhNrco1Jc9AfLhac+LnM/hLpnevsTjJa7zYOJp9tG
YUdkJN9Zm1nD43VNmQ1Cj+asobw0gfh8xrhg+61FpfUX0/yPpGx5AkQOOG1T9Vc6/HGz3+TsSV4M
aKiWJnmOz37cAJ+/VeGtFTknO7grSf3Ve8tCHbWCtThE2bZsYvybVqUxw1qg6DuTDprINwUoCDzO
RwjGMGzBmxwsnCfzurhU3r+Jyj0sdM9MZ5LHN0FFy1Q28ExsW2rlHj1G42vhDXBnWc6Wj40QJCgX
tG0E7+ZbctHz1jvvrWF3FPzr4VhtNWHsLx/N4PEh74k6gqGAaFGOy0TXLE3iTw1vmw0+14fvoUdH
KpczUp+t+32w9w45sd626FkimAFK7xR81qnwkl5Yv/5BVwaBk+/sK12NCTWI7zCPlNJ8PBV/v/Wl
4O3mLoVjklGLK87c/ceTBghAyk3xOlIRICo7vms7OaLzhw8LQdnxjnQ9gsSrEyVjSgdS2vUpGWpR
RYtKMKch7nDSx29SC2kPLIf0Sguw/eNOoy/XjjGp/4RVPJP6OtWEGCOpqa3Rj9m4i+/OmSaRVnsA
6CY0pQhvH7sRlmkl9bPWFXOSIRveU+J1xgGmstzxLbMP5X8mRAKMvOuptwwy7G3FW/ANBCzIgKK7
VnaQ85lMGR53/1w1xU5+8E87vnzgXuDO+5N+I0YVAc0O4p8xXXNC6d8chhyYB2bZtxKBBVQNTrqm
UML+8CLH3jkbHaC2f6kXd27wCyGuEi3F0EynrXaGMgFFuoZu1Zn265jUFik8+U5W59tjc+xE3Qd1
JAK1VKJIKlc4upDfkNQvf9l741o/VlS3ib94rzh4DxkIKYXGch8Hlbbg+SycRxysP1vfyswCkF0Z
lbqdIhJxJCnE39AuIO4p1kBy8SDCS4SZ1YmMfYIPVICYBas2nQNeeUsxCvulI/kWGYjMsxqcyDdB
Mec0AsoaVh1xlukRE2RVuNZD3JmV2CX1sAPcZpbc3hsRYcwmgCw1R93DBNhUihCIsM39Di5l/nrG
Q2s2CSGIpS9H4DBhMz1zPe4R2V89gbovUgqIw9SRmDGO9GDADOnyBdJfIGcL88x1Jp23s2GEd7KI
QomPmWNyAC9PfZRFkSgtYwRUDybMg1l6L1FkmNoddbmX3RY3T28GNmBCVmEWd/iXN9xoCLZwUrbL
4NyjxcwuU9SZD2WqdZ3rBgbqPZXtD63qEjnAUA4PLifd1iNcbD9Lz0PVPQ+s3Omb+kHUzy47x6w1
i+kSdqVITeIc1JevFcF8SmuM83DeLdNrPholMdwRvTo9Btq0+oKKwkB1HXx6pOSbXM+MhbbzzsyC
QhALUrhMi95JTlH5LijvWV8QF4UcFx4B/gY1shXO79TRo4aIPrJXms85A8qJp4OPQ7fGPSAevo0i
NzHH87QUgfEiNFMq5SctWP/d7E6v1CA6tMxk2ys+0G1gX2zFDUZmO6Ad0KBbJPXRe+tQxgcxR2HN
HLp6Z4gFOYbubol/K7ys3ruwy2q+I1c45rzLJ+BMXv8joMkUyz9FcJRt6uJ9r42BOihTsSCP5eHR
pVERz72f8D9omHSox8O0qJOoUw6ilTttEQPupeAWUtB71VGAVMvEm4wWuMR9/opAP8GG6o7H37/w
cABtDdpOAEUraKwdALFD/VOK+vV4VFFxBGEYoOB3Df+fWhXuXeMF9ClseQJBLC/uqVL/gpsSApAT
opjLJV6RHrXQJfHRTXjuei4aplVoJtg28KJw7jp9kcAINETPWH39AgLtxvNViNenq65GTnoCxABN
5IxKMyMBuhJGXvHA9mD5ZswmxcRY7TJ2Aiih2nCCObEmR9PraMDC28MsNYyn5pX3gz20iEble2pk
/ZQnmL49NQ1Md1BZM0mfdaEcPmX5uLvqhM+hV3TqPw1ejVf74EMxs5ddphtw1jt8ss4cyDA+wnNP
2p/JmAwwlaw9gdStFylMXRW4OkUAkA3RnpEUYqpsOhgCQt55RvULgBlZ8iOqBga3TW9yBGh8tW5n
QNoHYxGCL8alRPs36j/CNYNQC0KsOCnkzx23DFH8sga6iUhYnktn1cdg3iIzVz2hgj2eyVfTaprX
eROjtDSeKn4TgsRsAVih79aUEWJeNmFPeJn+jwVrfwlSQZDXAy0Rut7Gq7eTxSscJ7l83nyyWyrF
ZlhTm9cqAQxN8/GmOsfK4FVdK8LYYEySIB8kSObMcfHrUCrDtQSKokGn2LS1xCkfCSY3ffNAXdW8
RxcxoWGzUqyDivPfBhXT75uUrVpB1s9bfDNl2guPmTkrqG753TNMh6hCyYQdOGutVWqA+I6pZSdJ
bjeRWEO68o4ZYmaMHSOYJqZvKTCWDu76DR3fUN/zNYHi28yAL7jNmq/JKDScyA04eT0nCUAVoMwX
emitzBxt+8Q2G8m3EgwI5pBJqxFaAIiCfmx0TwQbuoEYwJi6WWA0sSYkUqcKLuSaZtigwGfbNGIh
kSopxZPGPBxE3ca5FAizHKSJiOb53rGRTe6JtC5/M70R3f7jdHC+qBnkmEZ+I7w7HclT0sn008cI
k3oTqqeoLy0TQ1pbyZMLPdFbyiu6XfPbUaCI0CvF8paaeYcLHaPuTBZk1ioi/4+NUcY+twPEKDns
gqVke75QLJawLJ6yZYZ96kiRUp7TUydsa24BOmXHi8vkbzbe8iP5QaOlMteECsHRzbekn2+gFWYJ
jSgmMfSxLIUjbbV1NHgtAq/W/nkfstS5CJWG8CwHokzS9ICoo1k6ZUpsiW/WfxrH+X+ZkldqKPzk
jEVU7hVs/CcAXc0tFa7Xx/ZK1fVqiojYam36/RQvTIMupKIkj5IlPw0Qbezt4x1sGD78Q4e+MtVQ
UY7CCBeZH/inbgPq+CHZ2r2jwZfiRG6BmF5tJwNWjVph6mqdMs0t8AgJbe+r5O0PWY10IufWg9SB
n+UeKhtdfDfgM+4FDCCwJGyZeGeRXDUkvi1M9glnJrrYufPrmbNw8dRc/uwBvO8ihDBBoZO7Tu7Y
dEfCJbWm9krDpKEm+KVSWaKWqi3PmPzlE+I+/TWrP4SjCMCg4f5g1W3Ic8RePCr04LVAeGkAx04O
AbtIODbUkfcPOKo9tAIIRDabJSRrzHXbMd5arbgGJEp7qzOnBG4m3SYdECpg4jtuBWd3HrtY82fA
aHd2/FHhl/PwrxDLw4ARUJENzPSqYD2OMaQW+uTJiNFosYo5SEkY6BO5fpapROfzW6ubwDDesBIK
jERzvEpXR35ZOmZcAftzxhZBNE0N7owQOmK68mJPaVtDKs2LMh+H9mgdvpYWlrC4WVrn2lhWMEfj
lX3MDdpYOlVV1UY6pAggduLTgGa0ZHje6v1WBxrZohN8X9CcyLFOdjWbT8ioE3vyPfODIt7jqOfg
5PvSZS0fsONM2Isbu7N/t4T1V7GkPVcfuHW3UwY6dXmmCTUiw2dR664zsP3IcRNkOCFqbb0lokMd
69aQsCtoKjXVQdh69Rw6eMCRpTNwfRgwyRIUur/2JpBE+vr2r+8eZFitUHgGyYtSpM/j33ZEdUUg
UieKbqgspZmkvKhvbiZr6VWfb4F35sJo66x2ZDqu1Wows8YHXSpkV4ZIbzRNN8Af7wR3B/V/jGbr
on+zl3sWSvYBZnkLYAhFUMbZ4oC/ycRHqGfvJSUwWdYWUzompUNyeAmCO5RYWWtDDiJbCEXa4xdp
9EoHVxz86BX+ea+yBjpD+5OW88prr+GAfYFH13uEAjCOe2lcqM4Ab//dXbvojdhvInuOaxf/aaoS
e0XhSHHiJgrGi/UwSBVye0n3neSPuHsG79YqElN4dfV9VmOQMXYTnLaeWOZc3/4ROBSLIAoS9kKf
HbEc4SyktwfoeXFFYTjLU/vg7l7ODwmlofVebb3IcP1g7IQ+3O489MbwoqOJrkc7UIhWvOkOIlU4
LDKTVzkLkwgwCXmmHOmyByWz4NfSDfp55uyOxDqEmkduXg0VuGWIGFBpJkeY1niY//wlPcyiBetD
tajxt92nXmrh2MKZXG7gMnVHCFLNTib4w09zz9AtiwH0hRkTTrGOfPH4EulAT1sD85YWpDHenfSv
KAuIIFqLLFUrI/h+uTKFycw2B/P7G0TqrbfP3n8PuncRWsvm6xPkhrRV3lFNe6pDmvubWR82bLkN
JOiHiFmJ0dUFUlRz36eSlTuJ02eqwN22DN3UAEtIblv4Zd7EJKxQ9Tv1mh0A0dcN6ZaCCLEvj2+r
8lKNQdcrOtMBavPV6eSHTfwZeTTvCjwEGvn83bCK+BX+8nCx5OYEi0H/6mxbXNiAjMhFkUO1qpYD
DbVJdU9kxLR1HgDFT5W5Y/wWccQP49nQU2gsP6P8b23xQi7/kWrHXFubq9ypZ0z5lVW89gWLd08B
zqy5KfQpolnUqq/qmhWkt7tQNB/TuDYAFGRJgBNpWbDNmO60HikErFyEsej2hge3ytoVp9nOi6WL
r4XfWueX63sqYmnV6YlBRJzYJNT+p5BVb9D+f1Bdvy7ZVOPeKMeb026UtP5tHZ8XY1Mas3LoGtDP
/9tq/vOEMRQQhI56DeDwmrUKWeb1geIQ6db/3JuCiBrmr6bY83biQdCmPoVoRF0E2DY7svM3lMH8
k/o9AjEb+LBKGYZQvILiJa9ex/QdZP75rdotMt/ssrLxf7gDz9zFKF4FKnslQBXYZhYyFXxprPQG
zvjdWyJ/4D6ylH01qKnEAlwFoi6C2HzbjAf0Cb4VtIEPnGgymEg2hVFivSiyDHobBpWFX6KyEqx9
0WZrUA2ODvbz753+gaN3bhaftOGIdkE89h1aW7Kfv2txkZQCLn9m98q3cPhzRkjrwScygZRbPIcK
E6tBaMcfKb2bouerZ9bojZKh9EMIv5NZu88avY13r/btf+CgmoHIhtkkOhGgsQ3gMlWXOSKdwkH3
P5nNaq1mnj1mJrUr3oS2Uf4nm2msRlDO1Gc3BgAD6WnExXSONekYo8S0jTawfQzgkYI53mMBYZXW
mn0zQp1A9bCiFj+o49lF6kBQS3FnmWpsJniygQtXZH9drYytIqmF7nazYvccnoxDKcXRay3HEBg/
kNHg+aDGBDHA7fqDq4a0qm4PuRmYVuwbKLXD5J3Puj232CFQz1/La/bJo2MYvFAjj6NbtWXE/mpP
i6XnkSMTrvAAGQ8DJh8uqfHXVDH18Pd5ikg5MTdkZ0Q22wqWVemEAsuVkwBxd3XLbxAIKGRxOH4/
DsK1xvipm9lMwHK8Q0Hg2GkSboeLjYKu7FAbTFxVjT50aHxgUE0E0ofL5I1OtFjJnjzVkW+HEuDZ
g3L7E1DB3mMX21PvO6/3V8ALPLrJKRhZvY26vruVgy+Dyo5HDszB/Op2ZzrV8tfYSBSyw2i/F7zN
qSLb42PlSZ+2OIqByfAM3q2PtnSbss9rw6P46shzy2rzU/4e28HnyUynzAHoajptdnV8DWeHTywR
+/1+pNz4RrJOj+Uf8u84uBWe6O4wju9IoUoy5bKd/p+OPt26yejL5VEUUWpV7/noS6pYRr2VtWzi
ubuqkTYYLM9nHeJA6obbiCfsTRfEMaABHzsi79QTtYaU7mx+x6mz2159CuQNqcufD6HB/Qp0wT+J
wcWBXpJvgQbt9aLlGtJSMGEOylH76goYbI4AvApUOgjFsrnLzIRPUqvGWfCBVRotQrStHUQXxNF+
d51e0foBa9xwyqMaCWUev1q+k57rtz9QEaSxzoiQo3LTl9wqn1AueFZAuZ7jOa5C+PJ/Xcu8iUdK
Vw4yivvq/5NSCEi1U1gupOMnIUxjyoCUNyyrbiRnOoN1mJ1F8qsaH4VLHi37dc1yRW4hJTLs1QMX
nNKHTlOQDVQJA03lDBLv42L8q15t2pGKRwXIoT6wjhGx07BCAwSALgpxR7KRjx+JMVLLZGz5qj5l
O0o8hOpj9OPUlLna8+mwUzQqv67wFreyl5nj9Amv2J/qmNVidqpEyuruJP38NSI3CH73OmhXkYUf
xE1oyMXhcg0PoUKBeyr/kA75c45cpYI/U+NDQV1hm1aMV1Dx+s2ioItY3VaeOyQu/bjKa/ujygC5
iBn9uqiVgI7ZsnBOVaYpcn0eazYydO7bPEckoJOc/TG89nHP+l4BbcFmCGDE1pH6N+WR8figFYyw
BcaFZrwt+w6WywmnhsHO8X9ISUs7ra826sXxrZ/oFPwBW7/8IcHgV+IQSOJVqRv+dctThVfKFMDx
wCw14pquzov3Xwrcb5XTH1fj06hbCkJEnL3MGh7Nq6g9AlsPFKLbeUxJE5twndtkNBXu1zBi+er4
gDMAKmuIIduDavwYZ7KkDenGDuwabIWbQB+O+q/6GTYrN+i6Dz2B6Slkz5dcmqZ4ib8WujrphvFA
4M1iTNQtYyLvST1ZZ64nsV+1yskxOWiWvDLoNF8pYMs1389bZYzH2jON6Il7SFupZrc/5J8NJ8W5
FnWajTDr7Sy33grip+YZ+Dwdg2WMP9DPyoBibIExTYTeVm0642P7L84FK2WVfnf2K9DA5GsjjXYk
rcfNHt7RRFB/Urxv673zyaz4WFP60RBIQmdCeGA9iIGLU8sygysZ9mDhZkGhR8692jfExmub2LIq
nqNZL0Pk6HbQxhIAwlO5HJ6RqGl3fsqgAd3f0AveNxe3IJubosyc6mJGCbqiLZUndBh2xdd/w0Fg
4ulPUSZuknl3a9TshpWdsjLQ0wQZrm4cTHpetB6hpCG88CEJrfA3u6R0U/AxxWtYZLYpx/jjjX49
G/yE0LmuUT5RzCV31kA35z+QbTUySiZ9RgrFn3pwdUhNaK5hvHivsPp1XmZeuYsbIbWiMvZ66u9Z
qEeDfPVC4ZFna12+3tkFHwugGY+3U61so9MESNcFUmD0L8WHI+/wiPCd6271B3nryd0LF/9WbFEQ
Q7POyz7Jdiqeb+OIb90+1ejoKOEtTLSw0Oms1sH3s5rtuIMXIic0n8co7LIWs2xivnVexLb2s+DS
d5jV0/Q1x8mSIHua7+Q19r4+79mJqM603C0NR2B+VfECh5FbuXnf1IY5VTawOK/qjliHPaRJf2Oe
kvmSauRV83yTz8PRr0GFMy6Wm6VnrXxxAEyLECVjuy71IzD1xx+2ebORfftaRtm/FODNlUcDFXy+
3JjggBdTMHTBP8B+9YgYJn7rdNe1siWf7D0OuXWJfyChr0YpQL9oZIs1d4QhfDmt4a3IlNWZJRby
yadXOgTyy+N9iN81OcNiBRHNfz8SobXgqXj0bDm4aytlRdJryaUGjj/JQHFs7GcrQNf0BHcQotRm
UK4mgRTcFSfzjOayS4GaDVB9E8TxgAwm5bx6L09dEsqkGGJBu6iPcNPGs9FuK7XXeSZZlJl/K6tB
knLjtHmLQMB6gfSOQb8QNznMrfy4/ghQyQUj7wi5N4DUw1OQY5NW7Py8eoWHg3ryf5L4e0Q2qZNZ
88nmjWJulllylRvcVsvvn7DKCArsBfJ4Luz/bqmg23/5ZkPGEMi+rbesWoECqJK+ZCwci5A0hBZ9
H9LStPYCOto4mavNTxROHRVmwaVaLeR3ChIfjzZV3Kd4BYj81CZsg38WrsLvTltv2Tik9OP/tot2
BRJrnLx0o5p5EgJY337XOpcUqJVWzuaUGs0PkG6IVeHtLIi4AzVhA6QsV6NuwxPH8u5GEPixu8vR
cFnhvfSYgt8SIGacTTIbN4TJRfHoEIZiVfgiFEC3SWWSIcBkmAo2hh9nYLc1qyljBTkrmuFnKzl5
8XMGlExMYTMBCYR0TcWYXor3YCXE1xafDUnS95KklFNbsfVZM5whbdUK5jwnLtKk+p0Dv0hEAEAy
ZUbHF5ru4uWZx1BkZgf5rD//Ur1hAXkEjwFTNld94Ud+ldA/+HLz2hAV32qxlOuNsJPgn1q4ls7W
U1/WgHA8f8Y0bcm4Gx6GttMfwcGIAaPqZsOSuEzp03dzp7UC/sek6Q4iVtYmiqcY5gZspJWc4uCQ
cZnLFFMBRhZO2fOACcEZiFCpKonKQX31oUbQJukbzI8dOqcV+i9BjWhp9xcOfRvAU/tjfRv7WEcb
piVKZQcIoi/gc049mPH01lpM6XRURnfOeCQhfsr/BeQb4iJUvqGnzySHHjyxdEMtri4tn5GNZEiX
pFdfF6GdSnL5v3sNNe5LOYycoPN/Szqeeebg+pldkkAKmODXSMiJiAFJ892YQqODozIWXXGqNsTw
6UhUvukD/1xG/MhcOeKEBO0BHHhxhSIdyucmn/VVVpRvYlyaHgHZiZe5Kq8lQd+T/pykhzL/qGbS
70Iz2AK0Jzo1VLAtmZbHr7YvyrDwQCKvcFj+G+3M9r02fKoMukI+3SuSoL82UMIByJvKDkEi+ULE
7QfKs/b6FfgbHNKx7qm03ips28IR8BR47+1LvLnEDHA6olw7f/hRPhMsBb/J3/dlfokBnVnJ1Y6r
frsk5IYgdi8QNq6qWQYbVHeh56Kxrqm4GaiBiz6yP4oz7i6qkPX+AQLaOTwUpbby3fxUOHW8U3oe
JjQqyo9S/toHd1nY3Hk2fgpiaxMP0myvUe13UzBgOpYJ+3VO8Rox0x2O87SmycClXXlVZdzc/H9N
mDQT61lhYkk6zpdNgWfRUZhEt8qSwnQR5zrFkTLeZD79ANbegUNFS/y9jr9eVhtISysrofXlrAnY
gIQOpXphyLWDrwV6NMaHH8TZ8IBKtLW1RtJiDbcjx3tV3VzQ88iTEiIxBcEjDIjHblnS5XOfMtjw
4ENxKCzEiBiJUVtod5mmC+EcZtAzfnTQHvVsBt/6W+RvL5P12yYonfS3s8c3CGAL1CBWx7EOGbwj
JHgWXzx2dOTc+5054xZ4pt82QsrZreBJ4k3jrxRiftMg5QT6L0y16TU0yltgPqhSU2nvraM3cfBY
mHLpT5PvArsXfyvavT/D6cKrwtg6/ioRu8siYb3tYu5yyJRFOlGadQy7QvVbAOQW842D1dVCIiPl
k1s7kS7nHJLQZjaPv93aezgNe6yiaZXKw+pulDrzx56mQDRz5Z4fyTO2toJ5rqSFREjIKMK4lYiX
YkAPKGLh6WoS4kF9UWhWsmNzSCSerr7dqyrjuMkBNODLbsNB547BgZPYJ47tNPRkARslrff573Pm
QvsHhScg5bdHrHCps3CiHjFT63gtj10WKy6JflntFBnPKtI9zoZQmjxRgFkBmznWh7j2FfE0cMxC
EtC0F45W0FXm/wATzlATP22NGoMWMEJJeWcpjYe8GH93MVsPqrP9rYMpkOMv6POhi3n5W8LfFGx6
DOi3JNFH2+Qz6pSYJaT7HQMHdu3vC+i8NLu7sfQ2NXrcgo2iRhhR4Dz2VKbGVhQOwC5Sm3gEAyRQ
uWkrcbdniG/V5bFkMPGt1ZQMYr/XdCb4r8sIFrNc9SRFJE5+cpnMKy9iT+XdItPXbmI84Q6SsMSW
iL8aql+mG5lZgjzY5eFGTYJvwzyWSRODQaghm+MJSa90mwA6NrD8yZfyg9os9rZTWthB2kqa85aR
TjrTwTzIiSC6gutj80CQgcWoJoDTAsFcHBfAWa/4omjcUDly3EDgr0xQWnc/jtYAy4lRG4ZQbnkc
WyQB16WzV4T1ykw8UEoNFHmk0f1+aPPPFi8EP4cBD2Zm3R2Bxcw6tIBT7OA7JFTwx4DjiOpH2CWX
a/4KwchHYtfT+Ik00wJonyrF4mTgsfPt12wvMUBtdu+YP3Nk8bc/vAc0zyQewr1Q/u6wTaQydzry
02T7it3FOYw7NW+F2UODMDM5Cqk1UhAu2b9VIdVAI26M/0WrweIvLTZ+U4JYCuqU4W4iSaAbSbu3
aGAqandrBuhPa5W/zIV3ckndMuQuppEdu+0ez3W9xpcnGCTTodOrpFOg5tJ3uCUZpVigL1/3smv4
7YAggHorOYrO5wWV3JuT120eNoil5VKdMhPa0UcL36G0vcxN9QDLorEPzsdOLMHqZyPmhXsabnlU
qLU/NBZvmFg+2NwREmkhfC5tzUWY5EVOa6lp667xjJtuKVO9n1l0NlEoCPweJCt6jUlsOKuuoNJg
9kbCek+SKD8jP68AmQfNKJgsOcx/gZSOfLfDowtPkz+15lZ4pCmbvqwNjJSbr3ngThOP/0bxBS37
AI4ZU8FYoOAJFIMqErBYxrC/BU4kKJ04lz/GHeQdNAZs47287fap037GbJcgHHM0/+oASjLOOWiU
2eXOQNV0tc4q9/LFKcf5kDta3Xztyi5AsabakfluNoSXGbPNk3DAuRMIQhqV14Ou305SXmsoF5jw
06dlbDKNBg44ebGeFM0n/54vP9OtWv8IEVbRydRrT86i/7gQ574S/UmwVTkJDzgpCvbUFrT1SfKs
uv8jar6rW6uQ4+HAnLrbL25Y5mVrOX+qLIJ18NQYZdElR7njl7dElX24TH2mpMNcqRZKEIwDlIDB
i211q/fEqfkiNhbL/vJw8MwbmjpcoA+9R7kw/3KXEqvNwYM8tpmnwR5YLUiVbPziwWHscwIeYv9H
uBP/iCb+wBt7WS+ziFki812EuckmkR7w5GYwnO/HyUOYIlAiTHOZAI2itv4mxzmiJvpovlFNkKcm
Uh9/Zeh81Y5PDQT/n/jSyEPgreTF+M/nAHskTcrCXPwDE8B6NBMH9VkDvuDG/7NTgNOTewWZH1PV
8vPCnWfRgnXxKMEOp4EQSJ3n7VZWlxHmdNMhYfkuOmHZMlal0qTe5IgeQ5Wyv7C9w7sFr85QpEed
bUv32n2zawHgZOExbnr1hyNDAPFbw6sfNOuM4Q6ypjbMZX6eIRJIA684MI2bzrVyR9ML20FXSHDn
xznMNlKToWqbbhVk7SeU/MZwc3WfBUsrNMGONwQ8f553RioX9Df6uwFvjxAIki9FlG2mdUMzCWdz
k2XwUFSWc3aeB2DXASaE0/9gMFvUhH+9PQUYnGJPcJA4JKK0IcjTxwjgQYTwcYN2r+Y4rC4dXcrW
XHexgynJUtJwx074GVmSXjJeAUsuOiOh9YwuOaOxQ/8Q/PauGDs/H6my5GqgdZUNbWpsxdi985SJ
o5fGIs2kO71BEnpMAMhHJpBzm1dsHBeZDkvtGNRs9mPuIRYQyv+be7AwiSiLqQNsVVqDPQMsbGR+
A69LL7xPERLi9W12EpMReZgXC9UonaBSKCUSrGxAsJn+8zyzDC5XQIDnEf5ByxltFK7zLxmS9bUF
az8r6lvr4Btrt/spVaNe7R4uXfevVnV4CuOYSnqYC5KzgwqlkujZsnCDEl4JEXsnN2DfZgkql0hG
AcmdWA1FyR51ZiXhuKSTHg0uB/ssrHr09OaoV2FeKzqiGUol88ksg5kxZA1MCavqWXLwSfyFRL0b
OORFAcsLY8pwLsXH9ON0m+VHU9uRt/6bm9pBT6/crtbEkYiE+5uNqV80vtQIz4aj88qzZHi0dl3q
U9yQjqWGGLxjZbHrCNMkqU3w2k0WC3xgW0T+6EYShrRwnUTlY960ROzIa3tJGsvct1dCrlkNtg0/
7N9VIqvbu6SX/HYYr+aktDRVG5lnOHYSjk8YGZPShiMIf1kdmbsIWVVg949P+6BsTq04WL5g9M9O
Deb61XXK796G7Dl8nJfCyvm1mLdGYBiv6uLSD/9UDXorEdcozm8CwcUui3I37NTB4+1FfTkvZf3X
78vk0G9b2LMWkHBm04F/b4BW3x2Zi/kO4mmOkqAkngr3RUE9eSKEl8GiFyZfWudT+/1a1prWLrQp
VakOFG8sa7MpbgBajrlvS0SLNca0G9e9DVay69YQu1gGGQXbGjQ4xx+MBmsN6Jc1/Clpj4/CiGlT
DZWxf0enS1R1klZvqAI6+YRWAe19Z4oza9LVKIHAsM1ldLY2wK94YG4SJHs54wDsQBCXNKC1B6uV
g+/u4bEncXPrAyix/Lt+sG58tfpkze32/nlomAc+gWenPTzsuc5arUqyUm9QbzAD/2nCpP0jf8jH
R5UfKQLoBL4HHsxs887qK6+WQu3kwRewmkJBz2fLLiDX8VYFiOjL878Yv8N6R1Jd2AAErD83CA/c
ZmOrdAFohs/9pSiBL76zin2BbDBq0yF+D1XYGL7Fe9M4JfaRBpEfFlRXn2Zphz8GTtQ/yGRYSKXE
UUJUF4CdFos9RBZt+sbezGuJVnB7e1jwpyOs6DHnnJHsqt0kaNwAo2lLCLksLSHnB3bLAd7UwhtD
5RTtW5cWnJ7bEzPXYr0Sijs/oY1eDbXroAf2Tbnw1JG+Kzl+oh/3w/Y9ZnxOPVvRQEOtNWD/6ZyQ
iwguvR3pF4r/FivKY+Tl/M3fLl5Gg6J7R3GPCJS/SpvZ5Zs8+MCo1qf8TonM09mDonutdI3y6gOn
+tTpSAeP7E/gSkDiG/brhDX3IVCM4JUibUfUbX4+3WOvC2j+ppze49UZEVuYmrdLp5UB/beMYsxW
dvZvy6O5zJ7udF93d2O6YJfPzpWuZjgn2S7pmnMHEw0W6yT3hk2LQtrY1oPbbwjndX6oXxDia5Mx
9VwvIgF+enBIKRSRZ+4I26kt7cQ4qknk69sU8d76o1bTge0m2I6ApXfa2mt6w+fBtzW93VPMmVgb
1kyGrrmecJx5QRpI8JJaCpMBSSFnQ5Tn4mF/prc7XmPX4V6tyvzpCa96aKBhixBCNGOTBJrZgZTU
XPpvo/9rJ/2BV1kAPtF9RNs9ec2DPFuWqESpxa1pP66DkVpvMdY+f6k/Raagkv0bkmNxbkGxh+76
d//nnnAXeyGGfYOvSlgm10vVJseNexqnV4RwTLc+cc3MJOIopmLTyE+/0SXyTrkBGbfBkigCH1kB
oDROVwTOfU1BKUG1M/IVoaLKJ4eH/TgqFCjnQBqXI2wMUwZdifsvFS5t4ai5k81q7zwD55m72IN2
reemCcUa6k5QVeNHneqj7UALiOanneCYe3IwrMw7754HvFA+9QQxLgguqnzskTI2ssIzIqqPAOS9
Nvqt5Gwmpn1flYHdxjE+13A228Fb8eXrxLp0i4i0weKrxL+B9IPtkeyyAp6tDN41n+EfSwjlIGDv
s13JUwFQ/mNVdBqrvS9gDJCfz8GqEHFABvFOYZop+6ygQcluNgjf7MWB9QqBckALCrylk8iOdBLm
hP7JU8qO4uBucqpQirYD3DYOOh9zr0Rvl7BmN5r62+zs4B3MLMr6bu0tEqXjNFYFrZneTkO7uIaB
L0lmg2nEe2VPH2ITqgEfaD6oDXv5TeGZIhl6NlXaBkfC0rnvjMYFG/p0adUKonzV+IU4J1AhyHFz
gA6XznfbDZ10FtN3gxwpoAI+wvgsBnGPo9FrOoqwuSmIwxN9nkl3G9Lafs0QapZlGrzAGge7td6k
xjNRHfvjRRH9xxpoxe8d1A2WQW3mF0rnoQcTnpfJaTZWsGfGorAiHfAKv+zptouZhnoO1mL2oIr4
uKqjBWP89Hz+Dqo++7ck2dz6jNzNH7PL/3XBmwK+rq8HcGolb1O6IkuJokDjOoQ8myeeEyJBlkBO
qI9FgSsuz8kuDmKAdX78+n+kcZnsyadQQdR0U2GvjRQtZYtBC4WwhyYhcRap/x9raZ+2c75dtp0Z
4NSFKzLpH6tfznpFJWVqNfCFfYO1O2gph4brl2gf+yDDtwoQ9sTLGUxZRn9zgjIQBoOmWc62P3qg
Q7sq4Ld2r0iioVWDqjhF0PiyajU2Amx2ONCXoG8wA5z8QcvRgKuGwLdl6+IC94wYC3/wkWQIC8AH
f4a9pCd1SXTlWIym2DjJ/h8fv4uzp3fos86Cq4OU/a9mAVeVgYFlAp11F1n1mOyQkKgfim7avcQZ
MZr3AjwXwjsRk1UUTPtWlsC4CSN5kExnVXjZAEkE7dWG07qMY8fWWcONi1XjjSU2Ge3uAx62WxwO
pTwt+jfaZS/j4OeJFF8dxC/PmTFGOCOhlYrFK/1jPT24F/hfpxGXjnGNtEZMIe8K4lIJXrkg85/m
yTeNPUrEUM8bKdiJJQ5sN5zxgFbU5HRxPbHM256mkhgOEsrqGvYLS8e57hStBEtwE3n9/B0j348w
rkYvG/ecPOMBPLhbAuLiVHmO5gP0GoBTY7tfAHFqcdigfnP1t65Ky0qjPeQTsNGYntALHm5bjCg+
ctipjYJTqsz12v+eehNr+5flcKPmRUTTup6GIzYYsyVdga8XWdw5kaJSub846AdSrkENR4kK6W5D
KBsEfgIIVO8HrzcOPZKyLOULKiqjKv2LDvFKPh5p4/f1O5fv8M9jD8MrgbDScBGyuTIz0mHUX3CD
YRlGJX9IFRvjymGmuIwxG2oPryUCdBdcRdFOZU9qTFh6mwwTjhGkpmb+vz5SpZyP9CQm9A1C70XH
fn/+g8T9ITlA4EXCHgK25ZtWmBCLvgAIMPfgDYsiRRI+LB6X3kQtVgGNvzY3M8xLTrr/gdvYNFfN
uCkdjwsGLUTIUPlj2RyN2v/AI78QZa9eQkl7gLnJPOUyFCl5z+SYgBGyLRDV6q+7Sajw+Wot0oMU
IX37YmUmx/1k39dBL6N9mStHzvKYAJ5pDQWThAw2hETx0Y2uNtSmAF88jURtcGNtZQTuc9tKmC98
b4tFWNfzQLtpQGnVcVpduza4APvWHTfE97gXITGlaWk/5rkAR/L5raSxWPvcL2EVn+HH6bMjOFES
IVI9KZY0XJ52AwIjG9Lm/wkN8SkNQ2ubP9sw6nfaYLGIGzM3Dfb3uPQ1lWNKG8fRKWRgZs2F5fW5
nQo584zb/tDdb5AqCQSYVA6IYYTBojaLxxGPjU1HPD1XMDWEshK4NWiSMA4t2ijwpVWptuyw4QeP
ZIYiD1USUabF1cN1BlqfccBBA9bW5IooJ3lEpKrBCgvOA1VegVi8micAtZWUFfOjGG4gqxqYqHgq
DY0UwTFCF3AdXAoB9V4XRXFdgZiH1HV9TGllupa2IU4QoiVv7Iwkvqt7AbfCPTZ8lGmCb9Ahezxt
47plnW4mw//stsE8kkKZSynPgQR3Gm6hAOfG+2PVX3qwt/uwIm1naBhR4c6dxf4kxC3R5Z5AA4M+
jmAqdyOsRGgSFXGlsKz2XMMkYJptDB7rU8EcRVAs0ehCgLnYoHpu4aFWoe1lHd0JGUC+mLQ3YLFl
y8EQJyPO3a+KzrLrwLORST32Mb8hifCBMmmkr5BeyC/aedUKRfVGvz40ejT20lg97PsxYPJVmcPd
mQz/rmKorw+ks6WzSVD8hz4PH1SxLXsiF55mqB/hdxYGdzEbfYymdGiQn8N3WmTI7sTpHYdgjz6i
CAwBW8ytGazW4EyyAyXf7K5cfOb7XmOooUjVFEUPtpQpLtNu+AEn7zsP6W5OHYTlhkFQf4/NRXTD
nmy7LetJvkLdURoLLW0H2zjX8m2TgK+3IOh2Wjm7r0pDL0t788cCGCY03F+fXPZiYGrJHaKCecB5
AZoT9H+//Sh364btkgbgV7fM1BgX69o1X/sl8jfdXFHEVZ3bH8XFtlKpHW4l7CRVF73iyOZ5xNI0
LA5vsaZroZp9zBwwiu7fpIkDVk3ay+/JDtUr0gdxAwbRu8q8uH0qatu+sn69FJodpyl+MhpBxR1Z
uyav6hi2jT0Z4U72nS4AW59x+4fISL4B4E6rxoEbxznyVmSRG+/EfCjR9cTt2eQ676BMfJHuV9vV
rJjkngFULVYPbucs4DTO7u9d810qycQUVmHdByaEYlCmiGM+ZF33ilQ6RJR/BkrR57wJJHiWvAMl
aTP/ubdI22SWqMHeQ8PvdHXJ2abMwKTXjNXvCNAqWHUXVd0RYTqWiGSI36MIY3g7/ncPe/x+9XYx
9FmwgHWsx0RTIokf6KoO0jwb4MRJppof0qgt0PPNcTjFRuU5PPJB6ffZ1LbeihIm1d6U6RlM8jWg
lPW9WQtl/mvrwCEmfB1NVzokltYm1/+wqS+J8Ootu19D7oGR9bUbsn5HW8yTJoAhVN7sNT+ywNls
BND5S1wairNpZu0bDjIvKZlPT4H1j6D8MJvTgGC7F8YfSMGU1RPqm/6cUfwp7i6LRqO7IY9GmyK8
ck//Ap3bzmOG9jeNbRSsJ74yWahvRfGAWQH17b+v6c1qXLNBfluPVcYJ2mMr2CkRYnQ7TRJrhwma
WfrKxvfD9FDxta5PmOkLdArw/H83Y2rPyZ0pxu9MquASaonUCisayEv8QhbpILcyihDkdGuqtcTZ
bR0Hlv0M/KPJ7FJ4Dk3F8UWcWIYKxXkkrpPNlc4E71X39tIXGHHHLv3ZpjmloOY5Dg65BvSdbNWs
q4NHyTlKZwJWwo3UzZZoXJBke7VYlMf5SIY1QHbQ3KzeyzgY87TMEdN6NeXhB4TyqO6nCc6qswJm
He2p3Qgno6fA2/VxlGvaSMd8Yrp2O9xDzgH4P7v5hgGcubuKhoVUG7I/KVickdeVc9y2kKBFneqf
2AP/f9H9lWzFCYIZ8HdJnHhtvWhQ+Z3DjAom1TO638S7JBfZVuc1xrCP4k02FSDl1MggaRusQcS/
TvKVZrONvesFjz0vtFFscIkTamdJWzcKAfuF2fhFRnp3xkANsx+IVGxjqeULYjwRN4qOJ0+kwD/0
MSoTyRnpLv99hK9BN3S9YRd6yUN2FqXEZYuuCjuTX3NH4zc09KBg/efLeOsIkJulyjrHtVlRZxla
n8uE41bT+zKcdVrM40fvY7AmXAvBP2NTaUeLWUnB0V3xsCsLBmY2ihwr3mWW/7BFTZ35btDhGNpH
jwZtx820DLKCKSJsEXoq+dQrCGMuzg1tbYfaKyNxnVbeUrBMYHUxn9VIMtaGizNrZtocZezZkfNw
hm9ae6v21BIr35M21tbMqSg18t4O4cmKVXTKQsngvG/xzEZ75tkHaqwJzqnVmh6oq6/a1hwN2eCy
nHf62k1I9WCx2cTS1moe9b88Hf9WoyB3wcb3J4rZ7jm/PxzzMTGLanWrYyP3+/kj60OESPrJqgEx
PTI6aTM9Mx88nlNqeMIGaJ5WOOyOZxurgVDKN5DSJsv/snST3zExiNHUxm5cPF7KuqBAq7vWCHEA
/P6WJpl/VDdY9XYg53n7Alf7zqabll1h/RCx2T5d2NLl1sIQKFnlzFhs5odYIJOPZeXWh4y+Sxd2
RlP4BfhyzDRsc8MU0mFc1Ce2+dVBW8KUsxu+GehwMDejL+kSA4hV8iD0U4Lyy9EJhiLNA/goCwRK
G5ZR/eFaU5vOxu6P3YJHwO61CtBLyFnXAMwPvpfKA7QeP7zfxo5x50RzpxP+ILoJG+tAh5NTeXRk
78olvtHYHdf2JQ+BRsKfwbG9Lj8++GXtrY/DAAg+GbfNxwbsgoCroPpXlmPY98xxuCLHKmt0VGOg
4NNJxTOnyKPvE2Rezk870bCEVLqsYEJZ9tR2D0VW6xKHbSStTohD6/26HtMIb4loocmuwWcdQ5Hv
zHDehJ59Kthng//IxzGpyKqfECwe/7WfhFv0TguB/eNr4kpjEfrk5JJsXObcOWdqg8Ka6gTjqixr
2G96UfLCA/LtjBP7RYJdmU5Kbz64FbwZbTOSPIFf74zcg/a7clUHtVTxQP5u0oWf0QQn9jkKfxrV
rzOTZSSK/ZHIEQDQhwWKYY4wLi0E6Kat/G/7eX7AAA5TK1ctwMGLvHWMiiouyjQC7ANFA5AYZ35D
wtovj6PnZ/jJJL1VDnjh5pxCHg13D7LG+9gbHKa2OzC7Q2WpkxR8jCTtPD1jK40xSGh7sZob/w4N
EK8lgbWqlqVcZp2NwGrxWmBCZnIjl3Z+utDebwPL8qEhoSynAcVEXNDZs9FDCimc3v8Uh3iHcWlA
1FnyJJNHuPjv6rREhnkgyvUxcegdgJ3hBnO6x2rwIxz/nQ1CglVWDgwc1vvWtMptxWd2PMNCFgIu
3etk7/6NXiN0MXDAdUrKYfUcH1hEGHWOBNSYxoZYvb3aJQozCXDPzinW/onH46srOQFV8VTdBf7R
EbEUB9UkuAGZYsf7Grp8ChaDZ/eA93x8r1Dn8FAmBIuWXo3tynttZkf7WDW0RXjkpfc6GguH2v4b
RllUDrvFuqAmxqJB3QyPJ5gwx2m17ZPTzPJng5E1sCZB+wVy1FZE2bXhxHeZvrwrmO6xvdtr3EaW
qKHFYzeoAhnBGHCqt53s2/tUzoFtXeRLP30IKVs4XjHxid4e43ZacP9JjhEfaC3YhyYfizExPwwQ
xXoL6p1M350f+ZCx3Ztu4+BakD3ERLNytPS8T85f05hFSFDu1JM5Q0qvCRrMlrAlUUHEYULYh8q2
Rp1wmraERHnugeXUnq8foaSVKVoNlDp1fXeQZFgt4RJmI2Fne0pgX8ywQW+fXv3fX9DTw8z0YTbk
GVRvr/096Ja1gqnCAqiccWqy6kgNBmFQWcHtM5Vt1Ch+M//AgKngCYhfhOpUCng2IDvISLr7NwaF
eeRpRKEkOU3sZHn3nWDcbcQh47ytjY1TfveC8SM19E7rkgcgedlQv65Jmy38wRcVfg88t5fvaLgB
ZMDSG7hWn+nz1NJCFwP5VsG6AYArKsKZGuUiliGdpGC6cKLL4bhDpVjK5uPfqhNVPvrED4XklNrG
jtXYtwUiYPBcuy1JtXLvNoNIlUYfp0Z2PYEs2EXu7d9CcmH31Ms+pnruYHpKalTQ/Tw4RL7inOyN
xjB10rHMQ7lTlyH/zWitNzIklfknsJSAt60wa0T5W9Zravw6eIYx4eFYrMlJcU2S1ar8Io2D7/pF
OuP4uHrAXltRzp8Dmkc/kV+E4hssHT/DxMvZagskDKkcpsORgnOurHm8Jdv0g+G/JOzJR1R4LlRl
qRb87JOn1GsFbypko8GjCYVrLDobsLN2giIzg1kwSq8GRKd0UJ+KSqB6chF+W48CGAwMpVgNi90j
MtnnmqatXfdrbdSZwQ+tzh9DPcouqhFoaIDENx4KEndAHMyXrAjnTRqNV3+nUyXIRa3fKOsRP6Vl
IPZzEchHih7zhE/zfZ2ceiMgaMtCdRclYCy2/zg80d/6ZuqIUw3FrtiaqSGgL/K0vVf9gCkdOvS7
vQhmeQGFy8DVNlhWpbAwsNfP0eHlhRn+bnn4qvsmoHImM+YrIm3Lz27lzP7vs8h+ptIVwnJYio4p
cHxuU0wDve5ldU0LEgveSD2+Fx6TZlbsKRKEyrMV92S5uxY0LPKanJAW7rLV8+rrnWy9D12dSp+L
2huKwSn4GfA9hDpftJv/I3Oat5Zh3A2Ruvnocnz9w2z49dMcyWlDXvrOs/d6/6SqrFITu/zlbALG
SmDOg2AZ4TlGoM3EpuB4JLfBBwEkp2upiK5VBdo9Q4sd6YRe0pvlni+wQtRay1oMsz4Of9J7GoXM
1HhcIAN8icnZLntOrtSJL1F0bpjQretZV1/mUjyldLExk6mHvwCDZMUHewVmey6k6pe+CGK00bqI
mxLyy0idaq+dilVGq4AQNnmpiTCwZr6qPKi0inqqOWr2t3YP4feDAcRgoPtdT1jPX3NHGXV8o4y2
hhPvm+Gk3Q1EbRsGrJTCAWRRSfaNDcd/0ANJ+mXCiqnhzX+ttG2pedZB/xSU+reVjcM6hgAcOjM8
sg4LeafkowrpMPVQ1rDYxR4AtJ025UPDTCJye2QwrswKGhBuA7dbRWcNpCjYXAA2HFm+Lw1E8H+z
2zCxOzzneU3b/0wl8LmHB7bhvW0Gu/WxlEH7CEuYSBNFCBDD4UmFr5pdhv5uQUpteKx3gtlxme/G
eFtbCbX83V5mn6w6/L70MrIB2K+9XGTniJSEE5F6o83iYSF4T1d7v6Wo4tgjd5y4eBmD2PmuL68p
o2ktpZY9zRTDJvgpy0h9DYGxyM1zD+E/CWXAbM/ILs19e9fPNqb6G3y3xwtxgHYjlCmWIBTbxA4Q
ne0xoAL/fqSB4ZIbs3nzpNRcOoS5e96YOkvRULzpEqxmCeeUgSOq+kY8GOWRv6CjUFS8v+hMxfUN
F41p0KnsHuLH5fQKBpRmjzE/DowgmTgu30aOyApEaDMO4AqVXxYlpHWv83HWgyb+F73BFnFwMLVY
RhbmwRbMYtZch9xGY1YXzO2iwuIGEYqSGgZ4udDwib2wloayH9OODhD91hkrNdx3keflAeQ+gf7/
Lw0PPNzRQ6jb21+wFASL+31Y21wKHfZhR70Yl5g8JwyCJsyQ4ip2EXmG3a1P23pp+/sD6Dpus9/w
eC8uckQK9FWD5ULioR2oPSpwEy+LVvDhtn6l928/xkFmLfNAU1HLY/1l+WfFZWLYVSCzKHZa1GhH
56ClcOeWKCrze/LgjyZfDKMSeDJplYdZ0PmtFAPBRXZFWb8WmN16FRuNSaZdSvz1dRURLcXQ/pgI
47qBcJ1AAugkVk6wD6sF0+8qccnIyuXEJHr1Anj0a8XxHVjmEdFPz/OMl8OTIk7GuiDfBvCZ9l5B
O9nW4VQAgMhLWTy8pZ22ayvgZc+e3ZhhXxz6DL3KILZBZS/Gg3po41ZVf8x8B8uZZ5uBR5DRcuUY
50NfoS527+o0iETpP7wxzPL502HzXVMw5PdupLGYyTcxVQUgcYQz1vJTTjhNMZqUjxuN5kxssq+V
lLoGa7hqukI7IJsnZq+7qIxHRVC4kOynvlL+obe0eOGOX4bfUizGUraiD/2cDL2sI7zhfzcsqoxL
zFyG800laIXR4UNhtj24Rhr5cB78qaBqGAe6nF01Tc5kXKAR/e/iKdAwn+860bRvbGNp4PAUhjPS
ih+HVMPQPn63wNx84GQE9UCPnWi8LFe/iuROmVysFG1Q9lTSLUVmxlDrVU25ECOb2VM1aBIPGRPM
T11Oy7xHl5A7cd413DYSoFm5PmsuwxwziRLxCEd8g/0/8BH2cADQfB8eBXF82GKaZu4QbdcdliFZ
GTp9g0GqLAvXxAYzqj1iTxtLy1DZseNQph1GwSK9N9UmHgomkBbr44/Uv2bVbcG1MFHW7RLPPyBo
sWwkvEkadO/0fivPwe6tezFa/kBygP4nGQ/M3Sno7Spw2hz6nPlj/A9j4ZP/XIY9NjC5qEU2/2Fn
OSAO3HrP+Zdv8AIjO+2AoDIsJX4R2C3PyYYtXUoYhJIb6ts/chVFkzW4EyOrPy2MoDFdwS3WBnJA
8MNVidQqglTZ7VxZLoQUT/ovYib8CX7vIceSEtEMwMbTRcr3ZK00rv6V/HB9/3KBzVdMwU4brLAl
Xgej+9Bx8VKfrSY4WqI8Dg911qBxV7k8gqdkmfQbOdHUmfLeJlybsPRapXYSCtBPYlJHwGWloCYi
dD3DyNELeKyjI+aYQsGxvBJ2t8E8vJeCMhREgKXIvOG1PP7XTBnaVQmkWYIoEq3671QNJ/CgeFuy
2zs+yNJKLI83EOxg64QhprSJViC4kfakJcmpt6J85VSa/yiMyM0JtxEnZTMz4k1ZHEIsyYhbC1ri
qM32aKo5xxU8FvMvsBd6sZSrgE3S6l+NfOeXb/gaiPIOGht+pcy75YWOVfZiN7JX+v0HSAG1LiNX
MyHXvUwXUK3E4/fPKeSbhOYWb1O2I6OAbwr+6B5M3j2oBVw7XVp1RHCNpcMhQ78QkyyRM8o3jt2C
DjW1o0GjPGNusShreyn7lun+2z/OVD3LeTPqHo9lvxtxXOcTe/23AmKsrzmSa7SGdRSGJjJqlrot
WsM8Qm8Zvpd5ys3x4k1U+/zZxysrnHBtzY6eCzpbqKghqnLjyJe2rQa3wF8LfP4E2Yd96abpqwcp
ap+qfmWLoOu3A64tkwxqDvgrJi5kqH+gyiY8Ctj4kgMWUpNhISnn5h7GedzJelRQW1MeI+lcChoV
ihc4SpxAIsw0KdzX2Dj8QHFvKEVK1nSGVsjhzQYb57CFyFV0qOd9qM9vcAel8cYqvGj4KROJYqZV
ZjrX8SSh/IgpmatXsVfnB4HjxHspINdu03IuEMUemPXT0Oj5blj0g3wK9FhNgENWNcAtecqN1OMO
dIj5JwukGW1LGG0g3stWzSOS+JMdtZhsmTV1db02G6cj/A4br4Q+SxUP79g+L4CNhXkXONvJMxN5
ybiv87AhQb+v2o7Z0Fy08A6qs1Bi296crIDzR35aclEuuakqWfjdWLsB9x3Wlaz33Wy9H3HLOBrk
mLsJHSKqkLpjRfmdJL77tlXnjLSF+MD6Qvj6w44QinOhsywSPOazaFscN2wGGs0kRyRETgX3QMGq
hGVuAUtTS8ho3fvN/deQ11WP6y2qd6BX13SQgmwGpZxYken9Ib+Sql041eT3K6iTs7oaRgyTvTvr
4WixX7nb3IExiTxvWpjdfHCGJTwZl82CuWjl27oUWoSd0V94ix7iiRB6/v3dzbJxylxyL0UuwGll
eh8jNF5rzT9kRgScz9qrUbZPmL9HiOwWP9nI1ClllvIhboi/2VA5DrPU6K8LKiCX0H7p+lb6h6Ue
HPXNyj68ddaAoLUtH9lHSWiWey/c/Ed1GocVf3Xli2tt6XNjPR8ZzGM5qPC85K0XHa7rQwWqeaRY
iAkRygv7vrS4DzKRV0ZJGPUh3gmipyoud7DLo2Sm1HZe0/Hnt6Tl8SoOj0jpnvBi247bB66d38p+
9fQzzBFB9iJdmlrvuGHVYFnuiRsVXWRKDl/8oyxIVTxSs7HF1s6skzOMdjXLmbckUv6mhxaM3pcg
/8r3F4VaSQFCsMnCZzDvYulQEyDwPjY9sGwmCJq125VAAQ7ZiNafwqvDp8QFc18fHBYgIzuZ0EgY
7G+rsV5BKTzKpEADezjN3/UGCT9LiGFSWLqZZDsVGiLasKK51wIacejqQqE4m0tPUfF4qrf1SEg2
tFV+YodkHXRkNX1XuKr0kA1FyawPwG2sRge6cOGGTdzCfFpk5JGakO+TcYMOZskGoGGyA3ig94Ee
OO6tmAiGPedpciAN3AzuW2bNJK7mEU7OoWtWa5xU9VT0zhqQyWel7PxnuCOrqSAWEn0joFd0L7ou
J7bQKUTlpyy65DNwY4uKKB9QSX9IssNLFELsfRAl3S07PQgO6CLU4xy4oAHB5LZoDV00VKhsy4zt
2gf4ky8eiLnxbvfJVqSzYP41fF2k1RSpMOhqLLOqfIo6joRZcEKyn/EjWITwgbTQuRaC2dDUsgNN
vFOghojE1YMPt41UXm7+fngihsmaqx485M1HQkk61bD2en44YGdyAVUvjR+WOdJK44YiSNBQBHuy
PSHx3NkMQ2NpshVgrDIoatSzey32h2v2QpJvbztY3SwHxzUvmpOMztcA5ySNr2DLCmjN1d5vbQJD
aKQhjwzuaLhcHAnqaxUqT/lVTMBN2U3wJdILtV5kIqy3DjYsUhDcbV6m8K2RqgGqx6YrS6/wPDQP
Pk+neDu558Cnd3D2OPZpHyVVymG8bipYRQxFsIaM1qZfszbgzalc1qU2e0AJ+fNT9Sw9E0Hed1bM
tvxUzCSea4IfmL2UnFUuwIjE7EsVe3XBDZBYeGRSsWgXuZnSOXa+110PuyH+NXrImJ94oLqMkync
1geGQov11af+XJYBiHr0TO/WnB3WVJkoem2EZJSbso7NpnofOgUfttHKQ8YedZXkUDVKCzmuTKXc
UDeuSAnsmuWYozXQjpMJ144/CWkOE9y+K/LwJqkoBkltIuAUtUV4OdMPGjBj0c8cG8jF1jumPGvq
zW4b3F6dW/k6BLwwzgp090nB1JCUZxV4pb2LtpBlFE0/RSCOA3mk7VrpCrbrRd1sGReN7JTaPxte
ftdQpxFh1huF9e9+whOzjQwuFDketTZ2iowfka/0jtjxms3O8C0MOi6NumKY6kS3ad/6Z7n01NRZ
BUdkjYep/AyurT2HvYBk414fTchU6pUWiUwRXJ1OP5VkvqL6mjmpGWPVCLPqCB9XiHBC2Atl/PaT
83657AimXNQ2iqFORIaP0geSLm9tY4ZLuLEWmIA519dv8t3CFWYA3cbE0gjlqeGD73+lI3eD/Hsk
dBjee7mWNWQvlR3a5uR53K04HKWEnOKFmZkHX/8sY8UtJhjwMK/WuBd82uC7Obla6fAUuTUmgWAR
Ziblk0Ug8qStUUBf51YAQEoON/MqVnyhrsFQzV7VxHLTlSpkIKajdCW3achHzqPSClRSxgFfbwTb
Holg+aN9tvunFk2Dqk1N+XkZnKFsV/YDe20A2KSmuxKwhUhKKY//cRUEZfKuhivFnUPRNQY6MlsO
Ira22WpAeW4ueS5jMLaAnZWSm/Uhnz3pdkEq+XhzePJcI6PNs5D4WN0TshqIMXGR6mQLgtZ4A2yI
IeV5wwlKReOsd7F6z+qymrz+gLTPtiP/CvlHQNP44+sRV9LQhYN2sEUPIVQEgHdLlbg3ZjxbAuQP
uZSluvpjzzjadb4CIqRk3es++wUz5IUA8Li140RKTK0qf6lKWnhpzadTEcZRzb+Bpj1v6Kpm2FvB
t01fH7nSmXSRL46E3MDgJmdiV88aOYdAvdJ6VxcBP1gAR1l3BRST4SyRn2qWv+Gr+WGz6WMCQ1nN
T/OKAPdl/UctTBHEBFhzR57ZG8tl79v53wNciL0Nbk4LV0kyOAEXfRY0xDhpZguSI9s5DONdhtu1
SemQqvfDRWgQk2qLEXhD82rcihbSQJjuU1eicH9GawLfjAgW3zwCTgj7Mr8Wz+5diwtjXW0KgLji
vcIlmXStIJ71EX7nbvcGX/065cAFsKl75F5r5wZlYb+FgKM8pMYgB2V4xwdwh1UpMQb5OweHfjsq
SeCY/J4OVnFoBTIg+ecxBxoyHlawwxj1/wCzwtIciLJ1OhP1Kv8zpKFnUlbKttS8AUhShphNzQu/
XxK/dHupGWTMoFnPyh/gKEMlE9wigi83fKrexXfxhQHO8rDtzU/IV8yBfLrQQ0PuUmXNyJ1tARD9
X84nLURqn2JMNRHpJ7ETtK32ZdHyXC5gXAiOVLP17yzOkgsrzdB3tWdPMxpmsXAw12nJeYppw5/y
IJAbtgT6aJYOzVD2JWoqSG+XfKYrvRo/8HfODJibyJaipYN5FeO6+0TfhejJs5AwwOgsx+2m3Otl
bVeYc4xkuS9kM1euTlbUToPnz8BhJD+4FJVDWNjfuzN4rG8yZlpGYpNweF9oCcQWFcvRQWjXJSDg
gcSDrF4BpybAFbE46HGm7GHG49aHsqAUIrBJluSTjcD8lEJwJAeAiXC49peUERulfp3EdpNyLWl0
kgygLnuH7zfC/DYEStcdCAj/UanIuY6dxHDaHMkNcxnAOCQGr0B3f8joAvKiPJVWdg9BWT8wFv9F
mb7LLvIOwilWX2UWFrR2GGMPGEPAic6Nt/8gwG73QfzZTxrOGl2EpffWdft/tgzLUeTLPE4VKzar
Crn8kks0VvdB7tS7rPLezPPuaUlQNJS3C1DNss/96TkhsgvOB6O6f+ePwCFAsfrNmJlB1aB1hqhs
MtnlYG2rtv6T8z4eQd+/B2iT44c7UL8G3T4zaltIYg01RSmxVhjsc9/8L2Hb5gQmW1wIi2424I6z
yxq/fhThbv4SdeDMQv3d6OHi/c5UP2v3zaSB/+wShh+PQoMYvmHV2uB2cZhHTI/cIrs7xR9pje0L
nQuz2k84xkfKhkRa4hDp6cELOrZ2uvJPvkY3+RCuO8Skx6pA6ZB6fhTPGEbp4bwkxH4pA7Itt/nA
7MMB1P5t7VIPMZ9b9Q8dxAfBwe4e4oBspTcJTbINkm6VSr2zbPElQIWW1Y8FV7VmYKohrnZCeJFy
KTpragL41nW6p578mb6njBk+Qi9t/+u7vQxE4keSnFRJEvjC6kdc8a69WUXfxI1nBLyVmYp0cqIS
a5afB5NICEW242vHOUPHFNJ4xUDBlB4+ioOEUHc8lF8N5ghZJYURMMxvsz2RupscvVh0b/fn9R+B
R7Z9uEFgU+da1Lz92v7rfq0KF8hpH5kQ1wYkm5jlcXux+dCt0XdlkW56/HLIwBWPHHBIzMJj4cKL
f6ZaYyL6DoVMTR23lzGErlKGu3ooyo0Ratbkr3sbJk64J+s1r6ancarNdJtG+WguFFXT2Kz2tWgB
9Kp8EkwcIAmy7ni85LnCePz1HUobc6aYJAbsWCBqhF67L8jDD/GOlBoqoc7g6QimDz7iHV4N5puS
inyJza8M8wbdz4tdVBSNgSWTQrSCxXd/4QgmeCPekuan8Pxas8F6dLtgvUH07t7CDq+ZeeAQ6M5z
183vnyJ2l+xxafz9W6OxBLd7SzsSR2Xd/lHfshwKqYtagl8q+ZeHWGS4n7eM9yOG/BrpqUPYebdX
WCfxIaIZbCKd8g9MnTrSBuIXTVscbbcduST2o3jVKwSHkGkZKyMTIBxYBHZMZ/WnGMbvR8GrCQBd
sl5Tuwd+urWd0sK54+w8HdqLLmIhqFv9AV+hX8MgIKkrjtzpAjYcib9Z1WVS62nCUW1MuWoIH83M
/JuE8paPWXifGZaP/GuNBUaqrlZ7fz02m5dtw80AU9UA+p8Z8YBQzb5wvx5gyYWvJ+cubGLW5Xy5
lDt1ElhUBy7ch6Lu0P3faZSiOx1oeChZuBBpVBK88Vpv1aaB11563Abzo0xcrMb1jywQUuKsnSTd
3A9JlkkpCa1ty/7HZPAZW42mNzImOlDnPvBXchNcuWvTQpv4A2uFymBXrzP0gvGQ/qF6tU63UDkA
zU0+7TfL6EryUuWMBMf+JImqXWQ15HyvXtomP0qlUbrvnsKX2Tmnal4QHZnKeLHUhGBzwrlSrjmJ
lSELEQSUCCvlG55VRPNE04gVC+Ftep6YWn1pBZWUQeyOjvDYte0VGabzxpBBIRTyOdjnXpJFHVZK
eWs2zW2Atm5JDvifx6L7R1dVqeJlnocMugJdJQEagk1R16gGsa/b7fu30y3LPnTm5vzJOJikhS3B
26NHDZTJgm2/8jZ8czPLocsLNC6jHSLETOrBwXJLXmybPDH9w3z48+xAODTLsNMkAog2swP0XNND
llPFem8iIuuspVB2U8YPBkE0MxfachnrJN1GJDBbu9SFAib/iUdvRWzsRL8UwkZorNQVVj00Fl3m
VhIdlSP0gOfWCn4z0oL6bp5vsLPiE8UQta57gC+YH/d8W+cJxqAA7vQbx2GU7E+PsQ7yg7zWhyL2
tsVY4VnpaI4meAS6tFflJTkrh7Punc3Z3e9JuTivXlv3SoNt1jiK0t7H/yEi5SUusNvp87f7FwnX
NZo8uywgs5v5wQcrZ1gFj1tKstZLd2h9t2XiuBllNMsYKq5bQkKqzqYdiK4aJ9E4AKt4rh9UK8FB
7QWoMB1ufj7zJmuEjpahQCBJtk8btYGZzrdai60SyTO39rDZBpp2MT+GMKtsPDY19eu3SvOQJvSW
xe3ZfrHsFZsMFS+LJ3i1OuMxCIJqUR1nt3rDTXX9grGpZJwxggiFebAhJW/vuwEoj2ZHyQpu8A7c
lZ9BOKOWQHxYAleqPrTX0p25X9SNydTxrKKtMEgm3loD8MvNonhoZKP1beaHgtNGOc1GNU5n0WKM
Fc+3daje5A1YZTjyfz9HVjrfv7SPF1kZFiIMwErbtsKPVU8pHiTklkrkVezU0svYd/GYiTjDev/r
KgnEiZaqYgC3MruDMGsdwmEB9BPq3q8qV6FUzk+8Ivnvr/LU4oSB7HQKbC0Rvig/mYvUuX6aHrkE
vXzvxorXcYVVVGxnVXsTypWbGY/3rPvaZbqw0JembHUSFGQ4y2vrrNJOUu8dPrg/fRc6w85ZuJvQ
U3+iM099JULI2+UQr606XM5MfjTuJiUQ1G8Cg4/WFiMDalYsv9MYVCAMOzfRlT6lPddguAF3inVF
J/adkP6JU2rbRtEqn2MZ2bN3fAqqkBGIYVuG/h7RnD8KiLy69/ckXWz6BOQ6Il6Zz6nMqDOKVQsb
xhGEF682EVGZ/j+qYMtE4+o0baqT11+o/WkpYKlFJmaIPd+O/RZHumw+rBTahXHxJASgLJXyvuXx
RBi/dhuPe3biBZQ9qoQ2ieFKy+ZMZ1D7OW4l0AUTXzhPgNxiQO1mINSzjc64SFn9dTJeDycmUD90
dRVtavQvQASmrfTPLEHL41i+st90o3Q00ECWfaX0ZynnhY4BpEJA04ndc1ECy+BBHRPvoy6LY30d
JJ3I2P1/tK6br6UYb6Y8UOHdWSmkr7k09FIblHz8iy8g5ONLDMUaiD6sq3p5Mc9j5CqZenrC7RPd
RPDtua8fWDOl7sO64YUVXn2+XJcAlnnVfdacuFx6ssJNzyvO3ABThxRRhSoUB4kQu8ivcZMMkKZ3
ti9rkzPyXM3ugUneyHXe/TBs1KuTBtKrO+F5Upszrl/pBm0r9fMCddfWlUhG2TW5KPNLRmmugTbS
RWmO/YFKcJYactb2BMTO1/9zjt0HTJo6h2hsFOEy4GTfPxwb/6jWkKoVMVlOGy9bszX+SYyWTJJY
3qcDwtajx2hJluHhkWVbjcv9Hpto+7+PiMI0sEbt0CH1+lVr88AxuVJiRUHp40wfq1RnMK2WdFJf
E7QrjU9fBuNzRXk8muWV4E494/FyOl4FhUReVn+LLYYqyhjsaoRnwambK4Y9R794U8QYbq9r11GG
ePv3XZXLM6pTacUoy1EapdzNQ9i7Fdp5+kIUwo/O+Bda8fnWiYfUDNbe3dwOqXPT3AhhZNJhtgTU
f/FjW4pHV85Mt+A/zwUQWEs2Ix/27TEAD2PR8WI1eLJIkqeqBENgIN7RjAmHSfx1UgpcDKF810E+
vZsz9CKnewGztmhX5YAZkxc5po30GGwWReTDgr4QBEz+r08nTUJmo1BBOXWMc3tYoP9/85vwG9O7
Or4PHtlQIU3R6mahLZXLby0Ot44DYXSBKywNm2HvnfZM7ykUjUHpYdsXnf7C2jULW/Cw8VjQY7YE
npH7neC0lyCPywSZnSl/d7pglx8SVs7r9sQRZp15acdR+cNlH1y+mDMeavI6opNFup0hCAZ39ByJ
9ti38VMdKuaCvZThdzHHGMGer7GveigxQPDYfFoJNq9du6/USkjRd/M1Yf7GCYSff7dP/rvhu5m/
tSi0tYaM4ZUI7AmjTp8fNpPrfil+XpymivREbofqs4wvfvnQ9cnQlyqV5LiA689rctBs/DTMDXvI
6SHFvj23HaJfaXsDe7Wqgan3DWV4DmeBzey114wmhQ6a4n6JHD7KvVh0p58hDNXVXNn2jud5c56H
fiC+r0DiJaMkrxoGpjLLZTXcT5xwW8NdM7ETWyXzeJ5k+Sg67FW2Eg7jElqhkTBx1r+suDHQoL0k
E0Zxb6tNy1AhEkOMyFkkfpOUSBr+Mezxsv8ZmRgeQGyS4nwGvYZw9eNUrc0c+wj+0nbfO7RJmQcT
DAwh9GmleQGzwBFdRZ7Vg3BJO+eUzxLwicNqSixWGYKL+Jtc0Fhzis+uR7I2GcfWDuLBmRHenEFs
VMzQL+5mhrHF6+gktr9kNhfZwU//OzsOVPR5vG4cmzvXjNuiVTy79EjTioiRQHSSzZ9e22Y85gYK
2JVqTBO9/NbDl5w5FxLQRmRcKj6A5VRyWSbaYbDIBhCAGEza5xAFq7ZFKJiU/WXOxHtl1b7my5iV
2k/YNb0RuQPJ33aFrmITNc3OtLv71QV5ivyuFHIuq/p7cxlpisSs5uAMcESggVFYRmD1/RfMpzKw
nMkOyGRAqnolthageZvLWuM42YvEubnHtim07hy0FDTeH5T5Shje6Mut6ENY2T85/DOd2v2mUM/I
9O+hHRYbTjMf67UyE7ZKJScPfn7RZJHvpYrHWVd59pxk4g0Q4swCrke7iY5bFexvQpLvCqJygnjL
/iVB/qhg3jWpt9DHbbm+/bygfxm5TcZUdXHTGqmTpkNqAJgcCk1dr0xDGGVYu9kJlJndxoY03+YL
g5hA4q7tm6aNrwr8C2ZxZa1bw9R2ufAMdIUT2ARltsDv/pIvLDI8iVjQzLWv42QX3kBzutz1NqBy
nu5BIPf2VxUJQDgZeFLcfjkq61jWxjxxrYCWLnZjYebb7tJDAAv/RAY8jo5SRsQ13PPwSusfSGhB
KpzMH9OJkrRkDWco44xW6tjNLI9VMecNa7a6qR5qbkaJMFvilt5eoS8gVlAOkT+Pjuyso3gd2++N
UEUPRhEjS2a3Tft4ZkRf7BrYZuc+akNeZChVblcb8WXMi9VF571MZUUT0ti/OuNkyIg7OYEUlv9F
c6foYmoTn59+/VCLRB2ND/ZiPdHdILN3DivO+d35cNIxY6gXdf+hwVBWY/HFjN0BvwyXcn5UBVPe
lGT5Y+EHXbX6GdlGMA3GIjLe5iWx6htSCon+boBgafQUcMKULrNjYVepLWtmZSDu9vzKPKEyNNZ6
SZVqyerK7WuWAxdXW0Mpj8R/ZtijUj/n2JyPe8C7lpkw4SVijXLw5SZFqhjrI4an2N/KLIGZleTU
kbwmwlDOr6kdiCzFxD2IAVBPNqGn/geuoRc0YhEaJlo6wjgCYQyxgsw/E9T5h3eKaeYKS/HHwQ73
uT4WnDQ401Pb0OfvnnLrII3TP4KwcCtPCE1LXvobWryS5qu1/5M4W2mB3SHmWzEOrhpiIEukQlIK
MeMhFiqYoQ/H5V4v8cI8OJXKr7yhQq/X3qtPa1Whs//Z5O0Ztg3H9DXmZSg7sJ8TTDX+WXZCMG0L
KzyEiFkSaPScs0lGfNPY0oU2GHeOGoi0ht3RlVHyMF2h+ZOB+nJDtIjUXBxqAShRKftLAqQqqvLl
DZg2sLLQ72WeUKRPKBQGS8A93QjYtugMWA6+ttE8F/Oe5Fc5t6ZPXMLb7MSeDzpmQJXqKq63uSIg
GMgoEDEtUybbzqdVTqVY5IxDsK2CHb5l9CRwG+ZnYZ1B/cVhFqyRskeJC06Tcot4s2pmIzwff4YV
jg9di+3OMhiVEw0GkFoEI3T0CPMkVvBx1GyfBMEArjehDr3CNJfcNgzJ+/WTBKZ+p0F6XRyQFzPk
bcSENYLpISbLQTCMz+seljOtXbSgiCaW6/JYMa+xNrHXHYBP0idClqS92DSxIZ/kly9aQIbAcieG
i61NkW824YqBGOm0VXrpv0cD9GX/eWGIWYfXvjv8wa/NuS5d75JXkjvRoFFySkSRszqYMEBgPa7C
fyimqW1UTP5lLrapiXO/U2a7fA+L+3SQ70SstmXuiK3Q2BOXT2qiE3fa3LXV+GPMeqZ90iHMRkKZ
f1xaS2l6Mn/Q19lkbszwgcxFGlz1h0GL93E1ArLoZOwxkX8vygepI2NRemGr8Pip1BLqwB5fYlEs
9rbigrwlBCeUwnSS3YTWOz62TfNjdc5894dmddhafOyF5nG4cdivocnyHNEoKjK/CbQ6WcnP9Fkk
jBz5OeRd5cs3WEKlqCAg1F+o8CsJ/+IzgkFJlqQV797dDXd97QVpOrBkHtwqwBzcZkWzx85wPf2V
fGH/KueBfQ6Wo0AuTnASsSfbzCyvHimGWrm516pAsTaLNlGYZ9pnm3lH53jhMtAxorg+aS5yV8cn
CzKz0ux54lU+80pSkJqy4BEkqVWXDfTIeC96jIOAsat0wGbwu2PTLuyfwDtmD7HKamoqzYKn/d3O
X8X9U2SCiXpstFIIEbGQbAYRL2RVZQd5O3tbx3dezDgUh7Cf4wwS99cpwJnRJLI5wxVKwb7M87bI
pGzdxeyUGM5UY23z9LB6eIHz71CVrPvHPD67rmjBSamQ9adq08DHrXzmfs++GF2hYuXhhxKtmRtv
rcGrjewrLrCjs6Whx7SfFLqnGBICAjRtY9KYJjaP2y+bwBuJQ0gOkD8U/IhCL/hsbbgjn4knhmoh
E703RH39BdtAaoAkUceNMxcgoCQqEokFBtLT7mTOkziaOqMcTb4I1tR0rtLKqgrb9+XpDFIL+UC5
IuLcV8OoJVy6MYuYAUEB9c1LJz9cOFx4M19/tjOfX64Lr9EaOuAnC+fF7L8RFx4K5l7F/l7Tjuzy
MrAy+eqOECCAZGP1ZF7bCkgU/VMqDIekAJFJ+EaWa89W0b/GqxF2Y8idFzfWMUM1PW0/si20adWm
0CKMbOkpdbbZxxXqIJq1N8808/7roPiBgM9bptK2mChcFTknJEfU4Gj4/zssmzbmWrey0L7sa2r+
cC95HQhGGu1FRRZMdsKAbwqGG+/pZ2P9vxhrtdZi3v4RgJHLEbKE3197MNXWQw1zL+lu/KN439sQ
j4eDjPOcBvfh9lXjbYxPCW05SJEpqTOCAlkGXHJkxtK2pOo9bzBAgZ79xWimA7IPVyvpjjP2KjyX
3uNM6j3kcdJw9Y/HDOyS3tVncnuRs5bkAEXvl9xLQmWaroV908jEXcFPPtEjdsUia+x8XwkRYo9D
9eqWDJ1m6qCCZVesn3InVsSwUx2qSIN/7ZzsZDzk71nUdtVO8kAQtYEWeFfqqI+GBhiy2O7Wp1d+
oQpyjw1kbRbAyVMBoLY5bL689V2JezNFo5GKgigvFQJpKeJZdisr9Xsw1RFcdGJfQCd6XXkZXFVH
QKNNADsiO1iyhqfUV0cQyDO/sxislKZcZVYNt1gFAx9urZEvANzXjYkv+gsj1Z/L6cRetB2pGJW5
SyVxHCpVOSvdvwa1MOqvrMFW+98nGniRQlC3Nmb/6E/4F2efHSMpzSgaeegciL5QDrEFvDKqwZp5
WZe09rE8UyZED8lEZB9jEyFU2XbgWVq8/HHLkb9w/FS//5mxAld06SunNgpbgUH1LSJpRFhry9qs
SZkAv0PXIHK2hWm4O/i29s3ZcZjk2FCnvOTGjsBwZxjz8A4Xk7z86+aOehJf4gEAjorPu9Ze4X4l
HSPzVz8kEOcW1LFFCrK6Twv4bgLHoECNgjju/pRcuXOd6p4H+fDLSz3j3g/e1CVYsDNkO7Q15O8W
42MV5fj1mPGujxsdPkM7LfSZb9LpPpUadTEHaFfxxIwyN8XdNJd+NaEVuh7N0/pAf9b2/IednhyW
FIyK/o0ciJ7WegRa5WqFN4PRJBXpu3UMlrxiNmqMS9gOB3582clrfnDw16xx2DNS/LYCfRRNJRu2
aqEVH01GYXmuqW3tVMW+456sA/lVbllm0pK8BGXSNiJ96kBGpxuP/ubpcJH1qSL5ziDdupTUH1dI
54TcGbdyZ2AW+MWT7vi0p6emvOMLKD8ZMuckHC7CLfmXpOMot/n2sKDpXnl+558NjeyaFAETDTiB
wQjaNpFafCyxIBn3meH+4tm5pAAm6QzKONvsIVQNYP0cE8fqRMYduDBBhh5CPbRrXAFgj2lp7XbC
ELGPuRAdcwNlTJ6BTeZ1Pb7rZicCeFa2xywNWgHnZ1We6Mm3lWr7hzfy1nvofhpHbSqadi2GAjgk
tJmG3mJLOyZvK3LVve03H4Ra++vbAHmfyIoMSto+NwzHVxA+Fq3i1i5GZEbVLmGf6a66ZUjx+krO
eEEhyZ0Cby8BGeiBGePEaJ3zKSrW/4pBxUoVpMMThUoodtNyO+xc3YNfmx+g42ay2XrBHpjUUiPW
KdpQTDriJBL0/vFTJo1JrbYb6sIX6gB6MhPBO9vkOx9Eva5CMlKeLEPEFV2AOPzxwc6Z+wEyHzoG
lLQNYzJ/rQJjKdSGTgF8rWKF3e2HZmcy5OEfuLLWNN5C+7sJtzuI7PCd+Z68Sx3PodRDaDnSdhcU
FiPBOUciMpWKwbQMZ80ViugqTetk1xis4Q7sJsM8a6jcVBcHZXBGRU6ZUKPthzsmxBjdZTJqOnYs
rrZpmZEkIWUNsEDyY7AvksVim7FGDVa0k2S1dLHUtmtY/nKtohD9bXLiXQkC+WDIMqT0pF2WFIh5
uqjVw4XpGOn74bNB57l/oyE26yJTuR3aU/kWnP6qShhGWdoX6nEbzFPPC/qsV1ngTN9PDX+XSYsg
6KzHgpfCJEGjmjsfvuWVPGghQ0/PAVaCHq2lIJ/LOsXGgocAFvdFrFxF6AS626ax5mkdw9Akz88s
ShCjLkwfKS0PEKAfzUAxnW1SaoeQu1L4uk4o6s0cWnn+J4OtBdpDGilfy+uDRdE8lDDRGZraP+YH
RHz4aJqagyOABJtBnkSpwYqSsNACY1UlrzyMoq78/q203Z1nx6h64HIafxbvwv7w4kU86xoCQ7PK
N2MyznvzLxL1Z2v8DHmxpFlIyqgKY6RhnM4bOsS9GHkSth3NOB7WCO8V5Gd82mE14uW829uKrT4Z
GGZYNBUDdVPdk5bnEn/hmoTHtWWhxuZbfRaog6YeRDO1oSKSFhdSmlmUYpDg8aCEkAWWDvtBTN8p
pSrziKZZ4A/G5ueCkOkQz+WmvDsdy2mT56p7+fIslpiprb4zXIwrsMVscIMU2grhDe/GmFsJsPrt
MOIlIa5ES63SJhUfb5a8wXW3hR7Kw+4SuGfzkJtf9qiSkc1TUDubdNKjDXPLUeZLLgXUS8ME3h4V
KXgFpcSw0jWeA8DeKv9wGeTZLaVacAsYrlfS0faUblIIVKGt3KB5uO8lpmmja24wZHv112Q3vQ0+
8pwmFFAU50IwvDfP9CbNhC6VfSO52pJWmKGxKXQHHPYRpQFtXjc0jeDK23ao3CEFatYSbRDwEK0y
43Ohs7jAIaj88HX3B24xmjI+z6wLH5I7Xt+OHdN9i9DSHbLJ1v3PvvVkGwM0jwsgFLRTPO55BgAA
ejnhpBmvlZqBf8sCGpAD3bbv2KVbOsI2GwZzTtgAQ6DLPuiytFE6qzgifGywlHQo6E/gd6XsQzjO
QlBM8jAF38aFEmiGlIEmpIyB0Fvrv28GeY+JezhfRDivQUvEnES7laJlrZNgivWDk+gkmhEHWNde
HtsWlPKjmo7qWWdhUhxlfhhMDKTO6PfMNJfpPla2HZpfelk42mRHqckT5mgu9ZAwC4gyrfXbw79z
x1XHdDja4EuqYA87A4sRcMwB/8s4TAQZ0FhrQVSFBZF85ochTcWmLrCJ8XaWVLOGe2Ee70O9I9nQ
iErxKngQrosRt46XsrrhU9NoaZt1UtYVoTHEppUZ/QMQq2r6qr9x5yAHUk61DeUVFq+SbX3edfgI
F1ah1YfGD7PJ53Go1sltg5/+kQy5jMctcAoOvxwfnpxS5FQJL4ncQIAAla2kLEkXLUz3QkgA0SXh
gVqiL0Bhv1sxKt19Cza52p0qBSTCT4VDHu5zA3CIMSv7wk4mBGqyldH9hpdAursgVrMiuqXT6Sny
ll3d5e+ZATQtjWCjh/5lXtLxmEyJltEpZUZBi43g4Zb3aTcrg1nKThOBc5sb0qXLxZ7Jxz2CkARC
tjlLuKHdK6vEtV4PQm0wDGH5DeytV2SI39nZ3Fmzz2TOP3cWeZoCdIAkwQQ0K93uR9ApvzFZy7k3
5Yj4he9/0HHh28sMjkaJ0XmYLmxO+KTFgYZVd0nDIIyLxDG5VsRebc+yK9HLtKG2Rceaw0LwuPKy
bYtWOIjnPfhtPGrTrdDdkJMqgBiWAt7/JS9rRPJfIRu5Sq3nN4LfArLNqvj76Dncez/fyOWIXDKH
fcucsLv0BWNSIpxHviMfSc6o7OKmKOcuptRV8W6edAvMwMaQ3+Wq1AeBM92SiFOVRK/yllCB3pTe
gsrAxJwpWaxbgwNXZ3Zrn4+BLQcwQD005GD/RIeZ1ZTa1YUF8DjJ+qHdxS6IX9Vg2owS6isWQJQw
NJiMD9OULUziRSZwS5dPrjc1OI9u3sz4M456mUfVVogKDjvohWABex9kczuO9xJB6HBM7SGJgLUR
w3nOMUHt4T4Aaw/tYKF2r1wcaVzSN3Uf9zXjUCfLwV9j5KNElef6q36UywZXxyZkDOiHebrJzW2E
I8TNWHZl1GyGBjcQ5gqdg8p98mp9aa4J/gQyw3/lc6XCTSOt0LW8wvyN/feSL0FPDzy+1ROOPORZ
z2yfaFkC1RirNfDe7DUBmdTkfizU9Tglv6cfh8r1bXyCkvM0jzrgdlZJChGWBqSODnV/FTtLcC4L
iqwLrmnFIJsFrAZukfox3b2HbG7LGywSqFn6LDJiWBM2lQ0io68w0Idjs0V+9HGhHniOUBuBS92b
T9HEwoOb03KtHWJEZ8F++EeKL8lrbm6XtVXCoCXxdkMEHLB6dNM/dO3GNKQfH76+n2UuL7k8I9CA
SSsXGMVH2jQHONaxBW91RLGugZUVwJFza3wq511CWKeDpaY0BYxKR7vOY+pOhU77r6Y4Y7JwralX
jaoelWDDlBj3nZye+dcLs1Sk9J7UQecBX2njgQbkyDGVbm79w1X+mKU0ulqFgCzzbUPqhbj1vN9u
7ifnSrrDD53YxTwIMK58whjYCV4cwx8iFxeHh2RTDPuLHO5eR8lUvxPTQWR2ekuXut7OTk0b4tCI
CBLK2fhPaY6RBQGWMP9nxFppfQijYDU9niSAhekXwLpQU85fxgQfDsIBarJzNO3GPw3GQ2Cv1qlu
Z0+DzzZvZxrHUBCg9sCvL/U2FyUhn1dIV2Jwb5dt6WhvsJsAi51eQqrmVU7aX/yUZKbQ3K89dxi0
4u5BfrCmYduTO50sr4GvQnfBWlV/eKpDitpJJxAPrp+JeoARwaoksbq1ezQ268pcabV+2myPXX5m
mpjMHQuD3A+uCX8NRW2VSG0xJW26090lhUe4F02j4cvCX6wwRwso3hvYBIWtgh+C5VVbcvGj9BVw
BeKsTAenKRKyNv9WiCKckv28Klq6WTwFZxxycc+vrVNtL3uLgdcQLGWw8jKg4Qe5UU6e1s8dxj6B
+6TVlW6mLQS1K85e4g169YDas5rw7lSLs79J+0oLyzhDX41vhXqS0zYYtY1qyWtUKrHPABxYCynf
A5e3/EaEfQwPgVuzaIRgwdXvfwxQXf5yGVpc4WmQcSMKkEv8ZJt6IMbh/YLeEdHUhOhk+xyajj53
qoZ1rOW1k0/NsSQ6r35dJKwCpMwOhaPhbiAac44PlfpggjQ5j6B8JORCTsuP4EGX2lGawAFlbE+n
A6MGj65rJbEDS04dMB8hoKE6B5yA08uwl7G4BKLpkz1Pv44YgBH6nwixAzRz2AtLSbePiJJTZrv1
bebimO049GFNQeNeti94hfCqhymW8X1A5dgw3JBQyV5pqdSH8XTSdXLrWkeQiLdipR11jOeeDkJ8
Q4Ckr2GxIN91w99ZH7vO0nnfAJ1IVWb2bx2qeZwPKmdF1vYR7DtIqOxXonCeOqkMRxUuFeGE9+Qn
G3BDZP4URjEFmgEZd6Qfto0KJdICsm8KjLVFW9VWmQ3cs49LN7/IsWzO1iTcqU9h7VxXmpiCgdrO
eeQqhT24npqay0cSE0JnsRj+0EsDwADG8P0f0lmAURM+aXrTbsk2hnNYEalpqMEf7sg44r36H5kg
gqXiMWP7BpiDl87cdcCC5Boyc7YG2auwz8+cFBtSaTdNZWU2GfLua9kRodGKRVCejXxCdZteHrSL
RQYS1aLLNcjGfBmyQaATWmGAmoHopFAL3MWQAHjP2ZxyP7VzLHh+AdU9LQxw82b1G1XzSXl6TyzT
H3RPFRrDNn7RWrgTrmfumatFghQmJo2OT2GcqQNEg+tU1DCqHW/YTpBrIG+G/O5UFZwcxkH81cX8
IaY3m4u+GoqSpMXu8+SR4pdA4OZ/aOt0rpVjlj0AbEmH/hg1YVQ3kN9zeB9jIQutE4EVai3nSYIE
+dKkxqJZlzugvErSXmaCtc7t1QDkUZLt4TmjgTt6hgZeqRhjZ4w/sdmgzbEMozWYChV0CBunB/1c
18EvswQXtFinkv8k5vG498hPLBNN7YFzcqN3i1o0y4OfuzEEVD3zhbNkAx4EzfjhYeZJmCR4B1nm
2n4j65kg/kNeo6wKrdJQxs8XV1nUQc1NyqP4RRmjPXICPVO6uZQBmYxMBDHT3vSmYvFzybbvAcTD
B/1HRpegJLT1idRdZCt61lXJfsQYnPryv+A6PpTlIcNG3FREbT3QCo1ykmHvCGpJQvBGn4K1DUpi
IQCENdMJERmEqeM5DHl2RXx2nNYDHjJmh2xWVcUDTGb8WUE7QbkZpRRWELXb8qh0/AOm3QL6VwEB
jFKLeFOALrBhLxenrht0RZ64B4cO+Qrv7RXYMq/Uo5MOdduZUfZh7d62W8/CtjcrbP5Q4q729698
iN1+c1VW2WXxrHW40RVQmGmN4wH8/BUVsixt52kCCA1aiKW53MRZTUqAJaDYfDoJm6pc2Fk3SI2N
cLLdbda2z5R3QRo+4+cNa2jLlzkA0DerBViyiYQB8Zfb+8xLBl5D0rikY7eQobVW/W/zL+fTaUky
DUGmGMU2Stri/2FPgPzgKsVjcGyIThWhyB9bHJMQm8btrLeb3baleqE5rSYn8r1dMbR2cbB7mEQU
yOLmN1ZSgUNItw/1SxRjcCNR8QOacAezG0TrkukFEE9W2CVCqiS2I9/hGx9cIDmln8rROxBCeSQY
5ApglrLjGM7M/DdfrtI/E+20PO5lkILk8GZqX90aVbrElcFNEfG7MIpyrrtZTrmKYpVmKOraGws6
LYy++Hv3jGy4PgkEzPd9qtgRTAzgvO1rdwlDVYoYysMtnp/gOKORarUEJkfxKJCnRujwLCmm7c9y
ALL4QRrF6cFB3JKcbQcGarvNusG/r9y8LL42mQ+L4w3z/8wdLfBl2oLMQIU5ceetaMk2spn3nlUV
QJ+88SoI2E8UFYWA4oOEPBjJOBU8nYkr3S+RvnxcjXdLZNNCCsDfNeteTw8QuUY42825p50NssDV
7oBKr5C8YclvV/dptGFtRUAHvHoW3uPqQpRvLlKaW8xuAhguClOBcHjtYWDjhyrJVN20GTWTZbrh
GVTiaD3Atf0LEF92YVTKUH656hArRVfAL/5fnoNbdyPtJ/trFT1kiNmYxdmLeErt8hOowbqyozbt
jodiPCpEMKCVRTrtS71kVsmNBb3wZJzpnzK7CM7WIY+CPp1UT7iqbFaV5YAMz3u36uqKLIzxZ5r2
lArzKnwhw0TC+BH90sl2hdh5YgQpip24Q4HNNk0FkYo5uZd3N2emn3cpVBHb9somBD+u8T9v1Rir
mBTTlwZ+Iw+jmnBIXkieO6Kc3WRGV8bdoNNla9ZZJ4n2B9cUR4FTruIPK9GAb7IpXgjLq3wpnoAr
oiIetcYGhvv6L1/3ZbEIfY2bFQRsj7g3nXk7ld86+qsNzcWcF1/QJ/GEOWoJdlVAOHsy8pmfcB1q
nZSKiUeNpTVh/+toJT5JIof0WoJpSzluBqTbxe7cVWZ/LC9RpqdXymTwXecxN7XgKni1nvu/rvfe
uuqQYlZjyieYjUvlhgGrcO3Jjeuj+d13qVFojUEVl58pZpsTkGpAgUxPlxA5tEXKS1bAgpiAe92F
8zW4PeqMAX6kiRrpZ2XPVRGySCUB4860NCaLUEcWzU2q/REwi0Ql3otJSW2g9ydVcGlHk8y5Gd4k
nQojcDQ7z6iL+/5ffp4WSBS69sKmRU7DVRRvz8A0+lvpYqh9I6ScPj5S1USTMpqgQ6ZFJBMSOu2M
S2as3sgQCNRiCLrU5rxhecvslaWnMskgfNkc9WXw+ab3DdnH/XfIwQoboVm610jfBAnMswtb+mW8
hKEkiwV9ovehxay6V0IGdEHhMIkb2oYqZIzAarQ4LIlw0eHAiLGhq8Mrii+6xIK+gLPU+h66ONt0
9gRTB8TiMyXPyHRAEExpRhEhF/b/X2E3EGhPfE5UqxLuAJ1qnTIQqgaI5owuLLXl8P215aXiiKS8
6a6MVdA+kZ8j0JZ/gX+ckpNrBuWzwtPBqmY/cHP8LHoLRSr4wNFJNC8oe9cTr64DMvfqSc5WHVw7
77XA2ufR4HfaNcl4N6nFNjKBQOsdEznOTH5EokRmZmRn62//bG9155zGTou/AL9T6pYIqopdqrRH
kr81oGBNjJyL+SM+zoXYy7ZyTO8nRLWw0vYtFCehcIEQBiyySySn1mJSPZl1oRNGC9bybJHqudod
IrYNO5Pz3kcRe0dlz5/dxdiTnY4BVDbH+PFX6CGKCu7iVFC1+hPqPhMCUzkinUEt++o2uo1SzhwA
8uwv3EV3L3yEsk5mHgb4Ro3JzdIR1unV581jH61lGvZCBQS3zT5RM1aMh+LtVo3BQC0Uljq8q2EL
qCtvXh+svmcVTU18Ajfb85lNgdBGpKl+PD3auKIIdwNmo8kUjubh9NlLewpSNtYpxTd1QJ73R4sa
RLqwoCGuaKsazCP4UmhaGgP1HRG2h+V9vxv38uAt1Zonz3tIMud5aDNmj5nDLXtPDqPIcIVZeW5G
8/BSNYAPwQAMEfs+7pBi+89XySJXTIek9hVXxkT0X5uLW1h5/VyIOMoemhOJiMhEVyrYyt4O8dpX
2oL9KMieXW0+BBJtu5rmCgtltmthJVFTQCXOfO6BmvoRPwyF/ielG+bRyeLBWZPmH+ZFCfFwJ3wF
7hO6EGsv3RJudJnzj7yiBWRno+xxpot7pimmgNNykev6/jmpKi2FE1OYy39+IHrL6mVnz3217UqV
HRi/poSP3Zj/hy+TTKEMrK6Y07Bner9alij4LiRYymtGAkm+8hhAM1fu3b5XaXgDL5enyIkyEO9v
pNs4nPwgIQE6nA189yvhXZohX/fpLuz6VuYLZke0YAcf9uG2h1FIWK3ZNPl3N4GY3uznkz1+Xdp8
vDUo4B993aXdptsMhx0IiX/nY2/bhP1RrOsEUaslUgWcD38tOhnM30CMe/1iZFkXJOa7D9wz38Ta
2fv6d7+ZmlYz9gKDg8H87lNkSBjycm2sIno2RR5vA6XazxmmMfMetstYisd98jDW4VLLubBAvrSp
bkrMQPPDcc2cPdnnYPRZzWu7/jH/BLc6HtDpSetG7iv1M6QhHKQAXglYXLbX8yRd5NgLC9+QKhuc
DZVhDf6D8VUrg7h74lvYRuKpsV7eCB+OV5Q/1Wznry/WC/MXr8b5kF4E8pqSHjaX1/u/WtSLHQ2Y
5SiTAOrIEyw9OnJmcNUjV3aMHg3A3yxihpdTQAhuOsZlyPeMPRqYznA+9ghmLsK0/nWQv4lP4LTT
qJbCMPuBzytPISths+4bu5aoNhxjvy2nRY8hiS2DRHGpadT4/yb9KMIo/dNr6nrObpnMf6dlLafK
FMt+PbUb+PRECbmYM3+LxLjVC+agVCCktHiYg5vylmUmOpJlyXO2fZ1juR4uUlEOvUcZCltSJ3YE
VbL3/YlScrSUx/yQwGOiaiLcx0SGTB38C1gdU5Nujkz6gYq3ErRXVSgIB+ARPRzaNL4C0ucu72n4
M0WJvqOlFW8ZLyfCtuMf7maGwLI+hlFJ2xdY60EJdKWSLo4QZJAYCzH/oRJ47D4+Zu+jfaVq8N2W
sVerXtiAqqxpUVmeDdljDGoVkdDTYuGP5qNg+HJ/bVeWX0PpNC2ppyCd1knTisA4EaJqqipN05lb
NSxVwCc/1SrhTnZKSI5XPMVZGJFvWRhfKv2LlikHsDGdbpqXLIFUOfTm7NZB6nndReiVezT7xpS1
0rFPV1ndtK3A9vwFz41N1KsJd6vv5ddQJNx4UevpAaksjv7iiierQtwBh3FeEab0bCar7OFqnrR4
kmcJywqXaV27VY0wBOIDNN5p6aLaJ3DEcWzGU+Mb6PhfTDejQUTxZDiQts/468q3sxmIRC3xtDGg
f4pqdUPzUWpFHTGUbD9lQl27NrtXc8ywyBVmoE4ummiw13f8AlfJ5M2gFUjHZGgfBiHYHi12Xtm7
xTzxbytFwrF+otJ7a3TLsrt/7ZNAWX649n1L6XvxHFJBWM+p45j36YruEmxOKZ3p7/M9FIM9dA+F
u7iNsIA9xFcOBxrarMYRYO6tgf5is/gvk6XwnKAZAX0CQfOBDGn3LMUS7fO51Q78CvWPaBogRQ9l
DADoxRMvtgk3BRUYDTbv9gMAs/BTOPEklv4BgXvkbuEP7GYaQIE+2v6Jb1L9ZZzcfz54g63BqEtF
j5CZ+47FbflADMgfCiAxFBvXfmuM1uFvHqRBTzUkFZ068SD3fEvxQSwDnCa2gNDLwstT7bwMaGQi
MkFTCdhbDTgGc1MQ5WHtP0HLh/ixEtrEGm4hYAEQS7mNuBVt6n3Fw5xxNVp1imzEdnEmz7LyNEBd
AunO8oNZHjamhZfM4sq8WRAko1OsHNzTxWbECVmSvOzt9yUN8Q+9ufvhoT8ylI1AMGawm3TZlOPz
331bmhGPjQMzDejNXcLoKJ45BmIQz8JFpOMI0jllrfhqsHpHZFEMK4moIEHjvqMZRAPUKNhexWAl
JLcpHqBxc/G2PLlpiBcmVmLK43FNrXwIdh05ksfEFyxR6W+jz5Pubw9UsNzzfpAQvfvx5gxj+p9t
7Uzd6B3Pezv5qnwTkbg+mUJNiXN1GAXIrVxGglspT7AU7tMxaV6cITscmjdKpH9tZoz9OOtrtxD3
l2Hn1mb35jENXWHYlqC9kCUe25A/S7UaXq5jSWTwTHjexuAn3EJaJP/CtNN2OYakeDB7a3e1jNN7
aWKNfwayAWDEFYeXRset/B9O3PPrU7tb5H5bO028C+TUZniUx6Dzh7V2OJY8gDUgKFQ7/gHRlxoe
evyppfCscR+mxzbXnXF2dC1eW0YKeM18N1TTt07cmQfgl4wgDN+SFeEnOUlkjWCaZVW8kCXopimp
JJgq3kJuJKDPGG52ezZ9Zs/nVTsL/pUxv8RzOhkhwcu0qQfvrsd3gBu7NLDJ0aUfzVcBtbONHCRi
MMDYd9ZrXAHVD+71Q5o+TxOM/cde1G9/DjJANbd8NYhc5IqdAg26vIAlrm4ppyd2nETA+s26bYyz
bbXWg54I8s3BisqJ+VKTEb9GNJ+2jer50dvNggR660eGpaPzIcE024Ia4WhCgppkUrAwCEVRJfUJ
/5mYNm8DWD0m+yNEa9sBz8B4q5xpP5m/v4DopjHw0M56g6M3t3Z/ee0NXo34oTt4lKkYQnn/7usZ
skq2x398amR7o+CAZ6bW9KyRJPkwvWiH07yA8FCsNRcodghGuQzdGDg5dDw2gtGg+xqE+V6T0E6f
VwCYO1IHXOKnSh/MX+remuowAyXFVkoCcu9AKEkWEq1YvdTaysqYuR3a/POLboueoOjzhRxKL56s
wW8UXDXxugRnlS8szifpVkLDk317xLTnUlGRW/X5GEAg9KLgqvrlmaIJ/gLZW6GBcKI4wMITQiFX
2mz7aYzElkXg5dC6myq4BdJXeVneUSKBiHT/+UqtXnSmwQTZT9DDGFipM9GiOvkMKsAedExpdeaC
BZ+mKLEMFrkZEwd6vBVYvrAzH9bgd3mytwasKGMqnmG7wEkb16oue3RmyhAbqm7mhXNx5hdvoUMH
rdQiv+B9NFuiEioFE110uFyO9UOS3cJ3bhlrV8Ulyiho1AeReE8BydqX5BF+n4zYfNdeBpl/S3NT
lcvUMl7ypbtVpbjTySiqBwlwUquul5BGin7YWWJG3bs12+k2+P4BNRYDqPUwh6PG8ZBcaXtWUtck
TNL0HGBk33anrztIcLouaanvRONfL7jjyzperyqNbNpaE3tjai3T9D3vnzzi+RTzvCDJDoEkDG4r
oNC1cNAgzYcGuCDbpaE44jutQf5fKsllxfWXuhIgTcUoV6T7zOlPh5qY1+z1iM7/CfopXBa0THUI
wsRqZnT37ddZlPemX7tg5AnAh5WU9iciUEWjPDgeIJwB1XKr8n0qr1pWKcxEzKVQAfGKUw4bCg3P
g7EzUdQLpv8d4uCZIzeOfhAYV32L2CaODbo/KN9p+L8s7NEdEyhVzvNYGGKyKsxnI9wmUV7/9uot
u8KfCLanY+44qZErj6RmcZCIBj2OwiHzOSZmPqwAjC5Sj5rrOJyfj8huNRYzXTmWIp87EBb7K8I4
txQlPRltm9/Eb79xPr101lvuUaCIfdFt0wtE/9Oyi+7cjKuBMpA7FqIOFzNRzJpIk/DurN9Ixr8m
jDvTWgHyLnT+rbZBidQ8zls2+3pygwprz3Q1hGxeElfHVV2CNG3GJcrGikYdK6Lt5tEXdcTJOjZG
MA3GEiF/uU4HOxXsLxDoZ/70V7g30dzJqZChbQVPXdmPZXh4tWfO/2etjGMuMQi3B1zj7gycB3NV
EqWmqrE5yLfQG3NZp0oIcchi+iY3CCooQfT0mZeoC59xENHNSZ3ASiLQYk9Hs3AxoSf23qEq1VNV
qrIumxi5bj/1/sCF4ByjPm8BkEaitfT14wSwxV8s+lbeGXU/hxGBwSq0o53c6EzbDZdbDgAdO4is
QK7SmQ9B8nhA/3VnpUFsSHkHvYXRZM7CbAiFAmO2KhsZEipwF0XXwkx2m0HMWqSlByHr33z2VmZu
YJWeSSUUFW3V+gTd53/9eLcOPm7ZPfZ+jYigbx3LS0f3g5gIgWvYAS5NUrQPq63cg2msoeZdFc0q
QN1S4KA0IOiPKmJOgTOIcPXX0bZbq1ZyqzCIoE5zqvWnuMwpsTZY858vWE47vdIIdNjAENXn8Bs2
uergwqIfqzdSofgcsaXDlVXHIC1zMiEDiCNQc4elvIBHYoQ2w0zcIXU1hVsCZtJflYdMp+ouoN59
zZeTLADc6QDST536qiiXWevETvk1YQVx4KJQzA2BRLCHJuUQ1p9xo1zbQqNOtEkGQrZAzHIholR7
JibRX7vALO19zL3K0mHs/ARgN+afVpY+ohv1q/xSsQyzzHxzGhfEj8fIYHk8M1fAAPNi8i2pNVVB
Gwsf1wEoX8AXIyrTyToI1Awy3os9XHtAg8NnvoFamsvYcn9pCQIplnUbcT4T8aXIclt6BlU38dcM
bN0GAgIyI+W5D3ZLGkdGovmRkHNYZrTGUak1/bPlxD7dl7SQO8ROLJAEIimuGveH1ZaNj4ORgBRQ
m9/j9dYWY6F4PognEWsyKoKdZa2nl2Rf5DcE18hs86jlduTbdHrUwpjPqQ0qRkFoJuTvZ0D7lwj8
wJe3pINQBXFiLDjxSNX70AiLrufQum4FfedoCO+tScKHJHrp9rnQpDkyUGyQO3hOSuWyUmTl55Ev
78NfpI+TwpkS5EQ5+OMxViV5OuNHW+i0nO+rL4/JvUfoy7XvdPAElfdnuCEzDYnxWx1+qxv0g4XK
0Lon3Fpe3iNAVxT9Wbs5fUkf1sAlQpCh7xRpqRrS9Ss94G7Ypi6pBXCXZiACUcaBDRVWTDS1wN/9
qXUueo95mOemDZn3G7hX7B4l4PJqx66NFLLbJ3YebTyx1b0dXsF9CBr/cEirRcWPJk8zjek+X7Km
C5aKslCQRGT92cj5ekTKqHZzDKm3ytTxr3qWT6y8y0FGBzZhE6dR3jP5QNXibRZul5i0q5unoYDJ
1Co6JsOwOSG07L4TDhgYwHWVKcspzjmsehxFgTOsMtOI2KP+LM+cdCPQmqk+rwCdtlbcV7nkJBPZ
AMeTvmy80GxqYlrI8SgeSDOwW/Gp+0VGb2clz85+50vBm0D6RYnRV5K8LIyDBjsevDJawrGVcalB
jXmvFFG1azDA9zQWl+/fh8WkOZtpn6BYG7OhVzXgNwJGlIpvlJMbHnaTWj/EZK2B2eSpOya0Llmr
pHv67E2Sp4WAL9BdnubZviw8b0YgkF25KDtqWofgyy8YgHMMkmA35DpGJxuKbt0bRLqctfqVL5Yc
RrPetQVrr8GlkagMLf0KIJ6xQzrFahTRePrGAK801qBr5gU9SoVnSNoGNpbk0WhYWM4+FDYNlWuL
yeopzqM9Kvz56G5hPGxE68M+t6UcvrC7uTRnsFPgls07DVwO+K0XYw5PJGLCJLBidZtVDF/eAdWt
Yv4i4WMgOS3iGkXDxdYdWzemu9xChwfCytrPc+VkYOv/WOxjyC9OVzX79djttxPJMOVBaE2NbGy2
5+QzHUUpG5Lzys9EsHpQypU8iZ+jXHx4xM8jKbe3ixSCgw/OJeRXYttiZ4hh8gNoCDeXYi5rkqeC
xctrhrUDnyurJFeNT4cdcRZEFSj7tWNyS7BaRW66pHJMq/GFQrGRpLYzgkFqBCELX7HyYzAeQjBA
WHackaAWDF+8p7FNGdhNct36oo1IpV72YhOFup+cxgx2gv1GXPul9IB0H53MAMJxlYr0folFePau
geHOuRfW+jT97PYiahpJLi8R9ebbMfMuAbDuDbpQIrOqc4Z/HfHXKki+TgKhlGa+z3FEkMDtXRUS
GeEwpTrEFDzYB7BUUOgTcaG7fGLENYbHXy7eClHuiTLlSdpNEOASYKxqR9cnTMrjm4OGAldL4Flt
juxzT+rajzP21e86ckTZMDYIAf4HUvXm8faiUUcW7Za4gaHCw8n68ZGOulLBo/9+Lpc8V1a9dOfp
b818tqBAdQKJU1q6Bhxf10s1XRACNxDLfY6ZCHzHUdoX4MM3ztvl5JZzkOb/zsw/pgjZzUofdacY
6FJvSNwzSt4Q5Kid66eBqXxpFPRjrVtQHtgDNgbo5bsKsAtlh3OBLoIu47BmGyxD7IYHIowre3XS
aY/T4t1q8eTfHdZwOtXyf2zZIVbCnXejes+0kstsbXLRdse6JBUVuCjZGmYrJt4kdoTOveCdE3EL
TpZUTcQr36FWMCL9mdUz2ZJIbtIzRi2ogg7eusfio8+fXEBdAD19iRyoiZWEJf8fl+pmz/H3eIYE
65dEsbJmbdlH4w2734O6AoeXnNLuhtgZhErE1pmN5z+LAUwtLtUH+f4rjj0y5aX3mCZCbr+FvjdO
iy3VSSk09BIJPiJ//20e7SSYSZjMRFKgdrkiCmbUGaR78JUyzS7ClxjbYyKJj6LMBNddK7jxhG+E
7ya7TS0w1UsbOv6I+8JVBJvUBD5IkZoXVDvMfx3zwbNVz/hn8isBU2zeCtCp6BPz7fAqFIoC7DOA
Kn8MaWqA6Nu8H5sTzCmXOMe/yOSu8GUsJNQGTHC/IxV+MX1QXtNn1Uiq8GMkNuXn1wj4WXNk+l+3
w3XS/0xGjecPrTAor9FaNP5BOK3fWeBGqeZAkYPE4pnEzKOXUutPa9se8F3NNofgc4R5p7lRreRF
g6OyjI/i7aUbg5eHAglvDVd1cD1nyAIUFfxq8XrNNhKyfACiXdd3wJnMJAOTc79uzjY0ONjzJbpC
WEGLiZ6golLXoqi5AoHjNuhzXZSWLT1lF1nZ65zt3pUl5LQjCgRAs42cV9tMlXrblxTx8Pluv0H6
hgde4gs2ourXg6B32Dz11QxZdT6bX4P7DykV/fR3D/w1LeDRGrOc4WVtE7+/9mEewBiX7iZfs722
unb2uKt1HswFX1YB2KA/NuzL2oTCMgZTboV06XYoAMiB6WZFjASN0sqCT87nM/LA6jueLfjWhV2/
WmT7YGmT1feLViZRiwqZLy7VjBY458uGLeyaEbEWI9cTO3pqEWq0r6XzoOLAmE3qeKfyVKIMayOT
CfHXe0rqoCo5eRU8j8JllYBvjybwbFzq7IT/si2IeQSEe6dsFZu4GRo/ZynS1lO46Y2pHlpZgQp7
wrrtUzd1qpCAjrpEtebSSwN2P1R7X0uO4qWnJoPTFTJcG67KoKq89LeQRjQklCvErd4XX8oxPZsi
z4WNSR3kg+NEOpLyNMcHdwSmF6xol1r0h7vS4zSTGlYpiwYIsAobOqp8xNepVlZ1d3NNNxOVCdop
BMlsqu1YWNfD79nQ8zdb9FQjJvTRlbV2iQtz1eJtiEr5GrS8zMpZ8UyHiM1xb0k/mAyYT3qdcCvv
3TsFWyKDJrA7jPsHOGxT1qJBHw6WLqwZwetckH9jsRTGaM3WO2gO5Ac8KQkdCRsVii2P9xj+daxg
oYhjOp32XxgRgDJ3VGYmQ7VeQ6HG7etdigX2DLPt5ItLEQfJvE7RgXhz3C/en521TT0ik+U6TyXr
nltSra2qHmOaadGpq757SVidCvuPLflEu9BI6Va3X1GCOedoto/LLhE/7kcxP+N9/uRGBVGLs2bn
sIbiw24C8kG+CqqUA2BE/SyQPIx5aANp6qEEaaN1A2Og4eeP/Y71sfJADj+O8YR5BO6cW6dcfNx7
kdyLEt6PaGl9SWuwibC+AiyWstI48vW7eN5uWx/npXNJ/j2yhd3e45gnq0nCrI556cCAeH8gXeje
QEqBli5wsA6EUIo+3JUObQIKRl9wr/N4DSR+PYZIUiOCbIB8NFQNAROcXrKUyukHnFnlcUprfUos
Q2hKZTvZOChK6UUkywCfFHMpEWhomdlPHwnSDf7nMiEW5FsF0H+wi4tVRMCZoyUXOagiHiG+nZ3i
95QHRxeAsP9MW9jWXBlJhe7BARBHwe2tTbwNvVP/p2beFIeTYMuyDpmGun9wEOo0lm74YO61mfiJ
q/nPFLwkesMCyzk0xLtK0YY+MeFfgp/r8cxQ4395BztD+cnbGs4CEYks1t5mIE2zmOs9ICapb4zN
ml+wxsmYltoyrKuTCjIvV71hL7hZbPrxqMpy9q5wlMHoi6S6WTJb+U5I35psG5eSgyrr4FL9TeNH
1+NeYtUDvEc0kd043ErCfPg/K8clCXTbToJNOUEnoqFksGOyVzG/RAJnPN9wyDwYh/nzS59/6dA9
mxfKsDSQcz9oEFWMTJAcx+HHLScycg8hIn42KxQbxu6OfqTNZ6LFjQlkXXwmy0Ie8h+WsqpLwiQo
ZG62qdu+NK014yEOwnpJafyJC9ZK/z5YiUbIXvG+0CpnNotjpLPMGlwrG/MW3jn748qBWLI4b+hL
4sG899XD3804vvu7Q5xB4LI1qeXy54DOTU82D5dlX+ck4eT/t0i108qOKjSio892/UR5K7BX6xSH
iDK+OSHjFaPIHEiLrO9paa+Mrn9sVSQHd86iqqWQHswp2cwJ+kAGDgOB3z9Oyj0P6QGCPgsLo6uL
Ef9BXI3uKeD72fv8cJ7DOo6lq06GJMB3QB1NfNTIUDHUVFMrDajwXNToccOGMRJJsErDCeNMj7/Q
4C7/4CeXKzVPwgG4JkRjwdE2NB7K9C+J8ZVis0ufFDG5NEd/LLg7RQxaJ6KBlS716NwXKjFhskh4
Kxt6ng6BuE+Em9jpd62XDzUD3GjRWzxtw7s3/05Rzpx5npNvAO9m/x4XMceJq/94ey2ZhgVgnXZr
Cht/aFTPXEuToKZ99nEsEmxJ7W1IrJI5AhbDO9Bc84JN1OJVT16R1jdDD6shgNAWS/M6CBfUd8LJ
XsM+Nhea9RZkScA5g4CTkarctALnLaQ5xFh1Hn8YWnp+NW1b2/ssmtQS5KdYQeVr3qcX9u7jpzXV
/iQfd8xjcO8kObCR8Y8tPIIO2AC9rNLTQF/2LAi/Y5g+RmNbdUoLxopDYOzpSrFCU0vWBLdBYyPC
WNdGsjgmHelFdiO9dNvnIUfRRDLA2tTnwMpGpU/sYzy8vVsglJWA3Oj2OprgiI4Fdi7aII/wsnSA
kwn7IUmLtRP2Jk/9l8se/oWspZYU7m26Xx9LT2FGaa+bgtd6S037+aExtWa9iiFi+fxXrkVkc8GX
Cww0yeKqkjjl+PCQeINiFXfd8TBLITlEUPewoiX5cTTbq0I+PCH19x6QSn6UKmzMMa0aULwD87tj
fZP8szcA0pniFfLfV2NbnKRNZKFjWPZZ68ddGn+0h78m+lOAJt420VGQ72rrQj+uyHoIfoBrNjs+
fWBosoAUxcsviG8v+e2YGLv//oT/XfYhwaoBCyoaeR/Bevcxp0VKvy15BHlRPbtyMQteQYJr1VEH
GhwT5M3T0dYSMblgeKsosU8HNUnbyS7WSyUXPfCiizDe2qe2hO6B81pweN0nz40qTf8ae+RKFP4j
6Citl/4/TchudoIowC8oaeh+VYbFOvXenFNIh+KuBgkkMQlZYTE3mTXDHYPdHR1ImpW0lUXN6bmg
POdHBPpLmIE3QpyCOiTqea4WWyrnf001ii3gsPXQg8xwYKv1HP7yRhKFNaL4hmTnfbNDGkAO+cRT
NC3HVeaz1LIiOUViREwAkdocjZcJdxq18TCl56SYzrzQKvzr75QxnR2UiylXIZHfe7t7v/bU1K2q
zgv6jznwuPVhCrgpVHhldv9dRq2GTrHOPtPSMqpTvENPOKO8T1VTNgbKGv48ZBlh96gBiWcS+W1r
aw4mH7lJQm52mUZmkIxeSH7JgEMwDCvPdXkKNk7StOL1guM1PYmGP0YOwDS03cENgjp3aLVTyqa/
G86kUwhU8TzSyCedEP+gJmqAqyBZGva5RjET+pHgvyYL5YR43KVOQSQvJVVJk/JrQlIsgkGz2pIl
O/Q59rBGlfJvFbgyeAev6upZEvCIvS2xyJUrffsXZIKlR1dlQ74cNkkO8cf2TQQGk5sNrtwZRyUW
O8kszMAwEse3GnPQRsaBDzIjKWKBODToF8p5QFbE1JzHLy+XMGTeh2Q6p8y+OM7mb1CsZEAvbmHe
uGKBACrHrO5Q+4EXtsVGtGYgmuXv7ls/4pAHr/uRVoFXgv/tGYm+yug5YOsDuRU1JT86qadmT7Ki
+V2hEtTURVoztHX65/5rzCnOaigdhSV6wEH2c6HP5b7XId+1kjs2ZQGgOb5eawtJpK7OecIQdyaw
dasKLybfz4IL3uAPlaoLMT0xjdfVJMAoKdQ2DwCiayiZQnuFmR09sz1UHy314KOQPwSEzU9lKuet
O71MsDAp/sIU60oT5IYgFIpLff0BD1V2978qKmr2zMB4M7YuG+BulB5oqUD+pX0z45Cnjd17MaVZ
cRKLgBAXzAeuZ9+DZsCv69NZJ8e58frOWA6sld8dftSof++cIuHnXlEsFA0CvwFOHymyNCplsHB2
c/MI8Pa6jp0IydX6n/YPNDyFr8MzddvV+y+TU+MFGk4sKx2nRuYSavtI1Xvo+sF4OdDAjUewVX+S
2g1GSgOyCe4h4kllPh4Kf19fsNGQXbkBwNxeNwXlDOAhhgYeZ95+r4ntSjVq+6uPn0zvI4k6xkFb
1zK9SCZLcb/TnFnQnXGvuZiV1H9c5aix8riLqNYnUia6i5ITubrvOkMUYuUwzhEOVYG6+26e6YTG
a4EWimub09hf89so1vXt5q/NI8dSwKCCfGXYSW7G7lr8G3jR324Z9Ew6ADDdM93XJs98jYJCBB9z
OeIlDIP2VuzLDHFP+Fj5BWrBeivd4fZbVfILH4QVy1hmR6WQJ7f65tc/osSFfKQ1sQfyKidbdAml
CN9RnXoJ8j9YnGg5rYGeo50jFZOCIcWwJsVQeqLE6zO2d4Yprw2u3OAUgD4kHmGaS5+bh2er4zX9
zO6XcIo8I9OJv2s6Vi9Malk5i9hTWiYqDGmTj5FXaboYd+Owoi/YLbcOTGCC5xESV+SCEGKeZr6M
1stGgPjExhRhIVO7sZgdbqY2WDIwsgAde3KtUBIFifbHXOsmqwXkXT42io0RMIcUTgJDsDV4jqmJ
ftqjz5MeoK+F8swqCxZmDZjonbXDWjfZg5yNhE86C8XRMh20tDXA6b/LNlxesa+UhjNAxZ9tRpBE
7ZMJhO/irxMkYvtSTs2g7+8SrtZ4eiPDRASmRi5djziRve7u3BqlYM3iieE5wSMN6iDQuTxMEte9
T8RNajd8MWWrD7cK7c5Khh32wwZQO4WOSZln7wE67oYWab8wj8002D+C9IOuNdalwkzFG5sIvnJ6
0RQ6o0q4c6pnT7AmMoyC5hacSMTxVJy8kqqWD2SqaO1rzoKzh7PcM7WcGJpZtNxlUCh8dmSeCccM
APtcRwPS+rGMfJDqjwHNSWkExb6ijUxwdte4LzpJxG6xb58I4WeikoQ/9kg0rA4q/5y5FPf+I4Mf
7/A+ZZGWS1NNwRGcAeZJXSOuM1Svj6KqTgieucQvMFT0HZTuQ0qNdrFHdDZuGcwet34QQskFcVJP
6FBZX2IMpJkoGpPvKQzh7vf62hfVapeihF7tLE+bLQ6KPD94G4/fYyOeTWx9EiJ+e4W6C6m/0YnA
AjqszLVmLPYHynDWj5BRdQWIa4TG6Y6OXDEh1M5qAuxdjaCXsvgAugaT5C9S4G7IbJ+AJ3qlES94
LN7TSryBhzMwowsee3Koz2mBtZ717qy6YxuqafjZS+R86B0bWXX3wqnl/JZgvyMSE2b6tn23w4G4
sweh/eB2Wn80fSjkJR9wLkLxLx2OECJcvfcV6MPWZDFGVa8EQ2/NwwsIkGhcqHsdySKMs0zrOMXY
P8EfI06K4xmmAh3nc3Mvt3qNQFeU970QQn1xiw7SXcUnIQSpQAvgcweIGdv1i5gxIuf181qwEb1R
gkUGZ3h5EFawsspIoFJ2CSgUwqfp7I8I9AXjMNVqRFVg6oklkySjlszq8/jz5dTAJ1utr5vs47MS
fuAiWDjmrwjmdH+omzng5U765SS8SxF4kKeRft5JFNeUNKXJqJ4mKmNqClG5KdJX47zQV7T+6KI/
PLe6QD1LEpIZjLMMa2+LDSxqBMzxmxbh5NkGngTnvTEWZQhR48A9mS2SDzAUsxWLUrHlZNOLGK0V
FLAU9mZ92qh8bOcE1Zw7xgAKoK6aAhXxH9S9Ri41nFEMk2O/1KOc0VDy88HgxB3qhHZ1muI4jGCF
0vtT8vGh1f1f2zVjq3U/w635rzbk5PKdpWe+N7M977TDZ88xbTcVgSriHwCXAS10bjLJxog8HGdg
BiSlZ+Ui47TEDF7BikVvxtfrhxRRWylH4+3jLmkLNKUruTPM5w77HGO2g8Ng5wf5wYg6xuKtSfj1
iReNC6W086swDJcUQhULEjMurxqxve2XQaPFxxMwYi4yeUW/7nAobIDMsOC/wSxfj/DAXV6YOFb7
ApCRcKHnP7gk0AIQjN2HvYqEzSMFOamj9A2Z0Xuj1zZpzdFacrkCWzyxOGipn+sqhX6rNGS5nq9X
8VDN4+stOKLrvHwj8DG4x3q74lxaXOdzUOE1d+RrhFAegTdQMryq+IAWgQuxOyxd4WDZPRf+EGal
EOnz8nw6Z+Uetg3Iy3ojRqgrR0SHIyphpkOqmPKk6QTlvPAHC6hfjt/CqqN5xBKmQXbrOrJ2cz7H
hA4nU+Hi3DHtfB2a+33wgMOsQD7Nk7fJ4E/3R1q6qCPypNm15WCLfL+bK/UJzrKjkNq7pFJGflpI
9FBaTkcS7/BizL5w9adL8/SfAOysDL0fTm20qmUuGA4tI2C2+P+BPlI7Nk1suukie0E9cY5JIhl5
uy4EN/zxdzoLrngnIdkFj0g/vZdyrhXlzpfDwtDuQmeOSZqZV4M0ZdSD+mPqDYcbwShv6/tJqP/F
C2s1mj7tH7w1bDeTrRwYln51ULMC+1jZmyLnfOFzCKSIqtzlEJKeKmEvzPXnTU3RviFuhPV7337F
duG3wc1YQyYrc+l3mHIiQqn0DuXe9sfk9GB80/NBLap2VDjpthC4MKmBK1DOa+07WTymXSyGb6Ok
Qso2ptJqjXBnndYtV1ggDJMuL8zxBPaa+J96gObsFMJc4VDBbFJwY8dXa8GXKyEWIZp32RVUgquP
AXcO0TalKYEHyjnU9cw/oNtZK7CQ1aZ3QpFPJAKE7KwFx22mW4b14gFVg0T1PhQ2lsGVl7uIfeB9
h13DYmlpBdMLtO775wL/rIBgMTvFD8bvHNkyfh4FKkYsLa2PQYM9LgknFxiCMI2aOKib++dJ3hZF
if7tMVj+XK3bbFimjSvb0Hbkf6YUe+Fs5Ip1N9Sw1q2+6Ld82UjwUCaLuCJIdW1q5B00gW8xYdJX
aIyUxiqRHneFYGwqaK+G34HydBAHlwu67v8yoNRs4109U7jHNuROk5bUTQYjkqwYBAXKJVxPE8Fp
gzMA80MvU8m4682xgi6IfpHzu6lRM9tUuxVrv9f0Pb/qcYg3cxT0Ww9VZYU4BXJ8sVR+nFgb3ac+
F0R8fp1VXxxKPHUbuALb8J8SXiGOM3cji9iW6PMjVZLYbOY1aMKsk0k71cc6gCfA7Cay+nT/2ux9
zBTSz8FM+KI1vYXzPNQzxYuO8X4Ucqi8MtHM/ZPNRZ/HuT4i0hbk9O6+n7yo1sd9Mxurm7xU1aUp
iTLnu6oE3w/bUfxESQdweFBb4K8FVMsJ8/SDcgiv+ayf7BAFeadPcsToi+XhKE1aE+1cpdpkpzLd
t8dT+ndN3Pa/Pg5j3+BrqF4PoCKWNlAf+NQBTjJwrdq64xh2YkdXQ4SDKjf1RnruIZgDBDFTthUZ
vJ1Cak26fymfwo+0xaLbL9I8CfT3KFcXdqW3gqwk1nKgtmqkDjiBUvtgqWLlhma1E7zn13HtM8mJ
PieFv8BJsJ7rxxC2/y503mOSZuHQCDT1Xap8C7fCAPTf0kYHtYdvM4agHDNwsaie2NbyxQi5b54h
8JyKXjWwFpLp31q9dgJ9J9f2p8nmpfETe6J2HyW/82IkEwnZIVvmeunaxgBqt8WqDyHk6a7jqHdY
Afpr4PMlD1rh5TOuL7plbIuUheU2Um1rzvY1kcxwUWhXk0bTEQMn1U+IAL8Xb34QIHfa4wLo4QoX
oSWBygHfMkJRgT2untXNd7dIxHRDzT63qOFFjiHCuxoKAisf5xyiZRgr/ZgDczDK8UV8m6CAKmUF
w+artZzrl6YRdmniS4YzPsueI8r7LBW7jlWhH2mNJ8X+8oUzPpE0e9FKzAwLdK8OAwIA485yKq10
SLwNDBgGm5TGnP/HwJbyC2y1nNj52LSgfcOEP0gLtr/6Kms0QVWdYZdQ9jJ8P5xe5Z0CQC48YBvI
V1jbIAGvrHUaNG03i7WAvv52FdAgveP9/rEclmPcUtJ3IsyYWvErxr7Hk2CSyXxc4RJGbTqEHvPf
/F8Bs8K+dbcwrFEaejEv16y0MJ2Q0caAqQK5wzaHEW6cTHdZcwqHT/JIVtoP37g/1/fnFcj2VK20
tKgjQUyWXY+nmYZ3jyLyowknGPlenfbcmIiNvfqBJaMT4w3b/KcKbxM4OXETlj1r8pLacLeX2ptl
4PaFLzuLJe9Ay+ejacez5mfrdT1zZzOqdojBBwC4f2j+4RfYNhoQzojClVucS+Cz+FtC7qv/C3E5
Kk2pKQO12hmSv2p3JhA9t89lGQH6oRut9exdQE8fsKzmzdgumfbYEiIFUNXQA70wpH1l2ocFXzND
4OIEp2fYUD5qRkSqp/B1gRMW5jQvG/+5AKn6if4MHTkkbx3erV0eEMZzFiJbXCMxj6z5PpF4TQI4
V0CfKr7OOa0m7bQzL5cS8zpmOrv2hwSitpJZUYQYMQXRrMvT2Kjs5hBgVs35gw7zArRE7HvD9C1l
UbdZYS0/ylIri31A/xWI9v7pgQWY4LvyhQHsCNGCDve4HKETUdBHPQrTBHscGL46Gh3/urcUheGu
LkwFVj0AC3R5VF9jcOQP8J5rcpuPl8N1+EkV6Ux3tL1xKWsK9+zsnEcX2mK+QPyMlmykFsmOXtZa
s6VhDUQiaS4GdrbH4tgW+05x/9uP+MxG/GwA+xEt++Zn8O+QXappIjwCL7L7NYWP6LOZr2b7ZElb
gzaCEUdrNS0a3Vq4f9fWA5IYalOM+ofrgtKSVNva9i5mI3Fag+VoebHOKnZHRCvpnDA+NsiSY0Em
bKS3xd7Y+B0GiD1kYagtPbeQT9OP8aFFhvWZbL9Ke+xbRCV1RJYBirO7bG8//W1b8SCznx50fkWT
p8CTA+aI93wYeyBpJnqJTWP4K2BldE8pdLtwq4Iyfp8pnzemu1T9c2jcxI/a2z8jjMh3WjyxEKrI
enyKwL/zwc7yuwcwnse9QbIN31VxZO4m40tYt1pSB4/fN+M98nu2XNPDv6c+zXZgUnnz4gL6W2C2
7XDiQES6JEyuiANF2WJlwQd+OqIn4in0j2MmfoBSHk/N5pLwGiiMQAJ0e+8eEMQyYhFA4kRrMf71
1IeJKegbf3CZtCw2TLGAbT1EoRbxDEs1RcLpT03XmJYDZFzDbGsKwHaW92iwwon1fR51Mrc9dlDt
/vfenySHeUZ/GV2NWdTNPQHfNsSl62YwTNgFqKzperA7WvDtyGsbENw5BIVKb5Y36a/cWrEprqo7
dsWJK5q1F4h8aVp3mwOA3sYmO3Y7O3NVhhw7pgdCfY33tq8Te58q7NyW7vi/RcTq4lES6HDjcJg2
bnaarCmG/IaITMIDM+2sdcx5zvUyl5wIUHsFNBVIonwKu0Lb/avyhN8aKtlMr+isojUzGKoDHVsq
5Pdw4JKi22+C/u/KJYmALyGIoexIKPVeRW4xc5BQiVsAHp14pQnt7YPb8kjcuF3pgsuhOfVC8npi
h8wuq1k/QCBVrGjkOQL+x/Gwtop7Uw+6BmLpWzq6in+pFqCnarTD6Pkci80MfPnlwJsBwjsb+7XJ
WaPZYrDkVpIukJbil42qxgoEIApTOCarb57Ga/99EH4Wt0Od14ou8PVnaW/0xAYx1YkT96wHVIve
7a50iXPWZSk6Yy8Wtu+/vQIzuk83M8XBbsyCn0BoEYz/aJ1nV7Ax75K5/SZbLfB6TcMd52dU+nSq
qDyPvGSIiwgnRKQaaF00GIjcsFlWROFwDe485mY+i5yCx4UBRPX6E5DdLwAG/FyMP9H3op5Xwufl
Zv+wC0pjGUfxp6Ss6xfkKD7HCv+08byJzPtgrSqb0YzfITPdY/5D+R9l4Erf2sQXeBY2R77F7Pu7
BiPfwM+09VD6rUP0tt8Vx62xeGpDf4HYehYkzXB6BkGDD8jCXW5yk3HpF7pHR+XIFxjOC6i7WAtx
MGNhZHtuWj9jJZislGaoqJtiR++VDw29HKnsjkhrisJMPySaR0z7cLOU5t1AwTJlxeTpVMA7gfGI
tE4q4Ozzn7x3CaLizz8lYhpcI4E8oCWwKfexUdx65KPzN7F7eDr7D9XtUhnYwJ5PxTgKvNybPcaT
033WWK4qiAeJ8dOlNSRbGZ81XRWv9ADnj6BM8x3XHl83YIOO6fg6z9pOYWgxQGw/HZ8c4CZQfrIH
BROWBdgd9TaeXgruW/w29YMwrOO2OuTvTdUm2YiHZunS9N68GdTAA4XzzA3ijUYV+l2RNrQYnrFy
ev8k2TvqOU+VDj0wVP3C2bBTFay/z1uab552f9RdNYsvXDS+GmpSBkjFYIdK1YwWkU0OpdCGaXNC
73kWDok37hdEARAGjn1CQHX8iqjco/eh1bF41rYopzDeda5uENQ5U7h6xceWw/EQpuv7Nn5Fsde8
1Hh7NchgRWMygQVp76rTk9cS70ATEzzKxdo5y11+MZmrHWVUD1XB5HivjC7mxRLpmiTnQ/7Kjv55
YdlVvxmgDYnJ5e3I04UTJ3JiEngcaaBmtyOEvqrpvlG4Xs4qG9qQwqqiUIDq7TIXOmc7hFPz1emi
b1js6RWtSbNbN9KihTJxIuYXQyxHnrpkb817w5sYnvtlntiaqoKuJ7Bsojk3CC6jCzb5IdtnOzJ7
qufq6auFAvn84k4YO66sEMMGmcCOqmk+c6jJQER69lIYyguBUAWzby+eX8wIv/v/Hve7SuD/76MF
PzL7VSrz6//qWjsugMF7OKlPMjD8nr62OueAbaN5Suwu811J4Y7IfpNEdCPhO95iCUlKd5pGMpPF
mZrBCxkBiqEhka+RuE407O7d/eq962LmVBk3EmiP/ZHhq7x9lnXLizyw/df4BDDmcMsrs99JVcyF
IKyiAvs16HDv5irHbLpJMFG4bnri+sJNW61tuIFIzgwVRzxvplnF46p3219LRe+7wT6dYX+gbsBU
RIBlHYC639J1o/hvoG68Rq29A1mJAm/d2Pz/IzKdSidbDznixPWoUTtrH/uFN+OGSK8VPMgH+VCd
IqgJJAfERELwmOiQuoCnmTBbPkH6RlMgf43ykG1v8VoCOp+YyUcHaelqweTMg79K6GmnwogiCWSK
VNYqXxFf9f0bBCsPpIXpY+F9A5N3U777GiTlxjuonr/ja4JFW1U5x8LeIG54lnDczLwIZ9TPgAOe
nESABml/dl9XcZY591uWPDr/ZBMqe91Zozi1hrxgfaAE/VkFqD1LI1u8QlLmTlkezS7ZuVFAXWhN
Bm7MOZZY1p43Vq1h/JQSpCc4H7bNO7Hqzi69H4OLaVeQhH9p+Z6wqsvR2nqq29We2FS3ojeB5PZA
i6vz4CPE9II3jsqzm/JMTJTlTd5nAu789m1xdLwXj6v99tTJdRycJIifoQN+LQ5dFiSqNCt/ylDj
OEFQlNwMwPRkeaz2QszEK8m6pUD3SKFA2Qdk4g0GUC9PeX7M3Pb44Ux6xlyqC8dNCwMm6HwQhtH5
7WqT7JVbaS5oMwNByut000gDmDC5txcdVO8Sd+tIyh1yDd6iD0HIZM7qmT+HC3Tkl0geYdVJsSBM
MPIX4CG9bexZFLdZtlWbq8MZCfOvlxyQ3ywYvt6CG+NEfqFSIUah36ZcPS5tcPsrWhravdyyV5Sx
K+v63/kZbtovFdiTo5tvNllXUSjbLym9wfmtRt4LqGtbJycNzEV4xi+HtWzCs6JRuFPeHRUWDQMp
Z6UBcs52Oa9zZ9K5wZTUHuOLgmcEUMiMyxZ/MoJQyWek4aCSnIoSYDDhZoEp8bpvxmjQPTxA91v3
CwfYzBviJjWNL+00p61Q2IZku09ja/dyv+DdGq7t2u3nZAJFjbfomnyE6eDb4qFJZazIqgJzBXkT
Yf7hGpYFmrolLCKREyJQALThzt7w7s0p964AiQIdFyVoHiQ/B0sbTz/pyibKFDpyDi53vJOADFvW
EKOMU0rSZovHoXm/Sf2Sa1r1fLZ/menqG8aoBjBaDKobVJ5Ny2jx6g/3sTGgSbly317u+WOrI0Fs
NVBVUnLArivFt5G2S1KgjLMJ4kg/Y3Ka61MXn/l9rzodFG3edsgcc+DCIH8qASdYfbUsgmgWAE9d
YM/XCaf8Rh6Uqppib73x48+rY+aeWw8K/m9OWE60hQSi9FtUmkYktq1P5QHw8cjH0PLfozo6Y3sg
pN1o2fiHLYOmXhYjXKXR1ufcJoaPSQlR4a8qRxyrwr3o6zsZMh/WvweZS6JxK0PdzNnH8i2Ly6SV
MmKfQXUTehkFNf4EYRQPRnTLc7yJVwDaBHr4sHSkF5EKx4kDjgateKBrq48ICoNwbS4VuVQd6wze
snenpUWnNd+gJS7BqSWSiwqBrbGIlnlSVQphoGzf5OBfkbskM0iuvcIIUUKEFWk6yl7l0U/pImcW
E98jj1Zn8JDrb3mn1NyORipfcCtSl+bsJiK4M1KMA5Xxt6leEneGaBQDlKL576jEbqO/YU3KK0jr
9yWeN9psbHVVa0hueQWK52LAxT6obUiZ0z8p6J4RRZHIyJyrrE2gaGXZRRn9iupOSjUEc0BS2Bi9
+JLU7fHd7AP4RZ+0paUbNMy27Hv+fDb6GspoSi1IR29RYYbcvcn/EVBjsvCFR0qz91quCs19WANU
MzEvtF+g7mVElQj6QPMlAE3ctszOG1cHZx+JpChFhhBh9pt8aopr4KzaTgRlDUn6hNusmrtwDlz2
BRCqCd01v6ew+sRphy9mDKRjisBH3mugHQgdnpXF8E6qa2JAKoDc//AtQZXizJ3xc5ij8ai1hdxJ
isCDB8nA3lebx4/SNNxYUgwcTYGpbibB00/Dpc+IKHGjKPzfnsgCW4hUXefyzSHtm7esK9cWNAzT
5Loy9OJaeS9OaROBSCFxjFwUm7Wo/MAk2V//T+pcoX/zorv8KC/ztbhAf17uf/y2MLbSjZVYUtV/
mS5Jb/4T4HFhmnI1+sHF7oKvkDWrU57oOtlh5H7vLtNOkrZrEDbUEtYDDuqe+mjOYSOnHKvh8usG
7CKFsjk5qY6KPp+nQvvJiL3IeO1OzV94iiTyoAdhTTGx+ktn9G9Mx8OqrlRpHe++8taOqQOyI2wD
vqj+cZk3SijJdihzbtlgOOybOlRuety7G96NEEW6Yun15bHgxqb0Z1fd/xQNItbohJYaqe4OfKlq
rW5bXeRhuN9mLlgnnoBuB4e8OsYDCXINfxJro0bnyouT/EZLvjBLYJ+NFA3v57W3kQC0uKtU0c6s
w4XPVHwchFSzkWa9eso5BW1i6nyzKbRMp/EkXtGyLJ6MZCUvTbbOWq0M6HrrgmyiQRoV1IQL65Zm
8rkyCDrHrtuzwYx/cWyixcLA0vkI7aorroRvyDB79e6kSuYVmOqgDX1Y8yrvMcwO/UU90VVWBVzt
HY0DofjuVqk4L6YnYPbrKULJ0mODaHBTXsJzwJ5nZXFPEjRvQojJDMHee9O8iE6iOtoZDpCdhtHr
mpm02CUSTSZXsl8LZehbKfhXWU8enYnNHEeD78Ps7kQ85i1+REqA7/1u82vMw/7Lfe7tGC0UrUVk
pKYmtWkBT0BrOF3J/znCyRaG8KxKIfDsc2Q6DHpxRwhMXrAQXqpgb/F1OfjBxPci08r4ogoJj4la
jqLpOx+tz72OzpLBjnPb1hXIXOET/Qw9jHRt9VrWHVgvcv7hwGUllovX3MMzhmWJLvAlqCZr7jjC
6A2ck+09KCG26GgZI86k89ZAEldJdwl5Z1ywql/5HGKUbwTEs/bfaSx+ZAQZvO6RKX1qyD/+n/Tu
/D8D8HQpkRqZ19UjRXsUCkJMXkrDVWIaXIvdhvYSAFmQBgrCmiquYVTyk3r7B/GLDIa5IkAzkTvu
KzbexltgBIFUJaRdEiZVZroPod47KIzJpK2dTckPe1qRDQnpKEUHU+6/15ZXlNcsGCH5KrfrSsHU
89qoE3aGqQx+VJFz7jqwVit+UKeibCP4jmcHz2OxpdZpTSyAk4z8tJ/WhTdi1BxRE67t2Bc2oB7V
KgMWWq4ucarowwMFUyB9V8uUgfsWbkmFd/hYYI747fctNSmhUy5R6rsKZCZN+uV2UwqvW5ntY+Ru
htsgjBJhai5sg/5JIP5i9ZBtXq+TpL5NLtP8OIV6Qmnqvi6c/GrqR+K5ULslC36beBYDCLIpIOIF
vzs51f03uTjXZwmXKbPKtw99zsNpGBeKqqAEUsbF3jE0UWgln3YCQZzfrj1xRt+gd/sGko9kUaoN
BGPtOwYxES6r7glorEiPqtkPB5z2yj9v7XxtI6sPq2Yz9FVIapGNca9nvkLt0aDCFIrEWiBvDaDW
c051TdwpX14q6KEzOWL9vy0WRHwwOoAv+Wxreb/kfT9Kh0ZHoYqQlujHNzxKSIMXc9Lny3jOl7D8
mGSlueYCwO3Q0RIj8YE7nBpwyiOPIZobPDEZ47zDJ6jzMdN2lvHKPVUbg0lmRj5eqtikw12oKMyc
A/ggd09ayR9u4u/RVsSMQd6VIR0Cd9MQZSkKIZgmqlHifVhJZqFZCfDYk5yTsbXJX9z58NaV6P8C
qtYl/lPAX7eQpdYejjD+xlhIwP1M7LxP48t8wY+ptcGEpaguMlUs7J1jLxVSaiIujl9Undmb+C5f
n1QY7jSnHcr4n9C3FGuGaP7o3643Rs99FxWhWWQ7EO4VduZlOucC7Eas/xQipvLbRwULt7qUOw4K
8UdJWRVVIVsspNJVV+WT1nUqvGqh0bE0qLbMSK7gvcdOIs4eKM5OF674eXxw6/srHPA891d2bhEg
nUqGYoZYVdn7MuMNd2Fif/rVyWiKTLjudWlIy9/+DH2mPTm/I57lLuwNM3lJlRyzKTR3BQCCUTCz
LOYiGYRizp0qdMJMhDOrFIQeoZWfiGT6y6hkvlnSgHkk+qXF757o93NCulhf3ZKR04A9v5Mk1pa4
2hZ4orbvyL3CMAyMp1PvGgmmMxfPKyoxm4fIhodHtTuqZZmbD3osZoRDSaDAagrRQLiXiqhMR7bC
v0c8ln4YxQdoMgXaXwnK0ZpFXYJkh8tNDnVp3w3oMdEn5YePM8yHVMdZkZJDg3Uz/JjrIHtnK4op
ONcwRM4Xr4lsEMX/9dGkoDvsZFT2f2o38OBAE/oYarkrxjGyeu8d1rD5CGWHUBoOJAJyocMp0VYg
kjreLTQuV55MUA0wviEkANIwAJ5ofHLXFXsnMT/l3BeNnWSZI1SiYZpl+f+qcnn4pB1bqWN/X9c9
UfERxDK5OaEo7TQ12vsBcpxR/9wHeMMWmw44WwOAcAhh7w2oW1qdrt8XKDt9NDY0qghk087PrZmm
7FR47ZKwmfmXZgWzQXLTWmw7Ml+sBa847sIdxg7iOht4aiYhZayF+dc1/iFirHkf3g/r7iHEI/5+
II1F9/b+rW15dtt4GkBeeXdg7/VbXR6DrIRa5lMbqXC5E9fB+4T/JD079Rlh8VdsAZrmFz6VgBRa
EG3UUXoa7pxRJdSAPbSSbaL5rjf0ngQsi+bRlG+1pFLWXWJPXEtv7Gi+QZAt9roEv9zvQrRFstma
dMGzlsq17tyb9KiKjUb65G8j8MiwUqXA4RTmugmUAf3yaOsyeQBCfwNyAvIEZjBU8Ql5kQBFLrEK
3XfpoUPph7sDDuwL6gzrlaiP6EZSY00NCtGaL/zKJ9+gdOFoGJ2HUNp++neztwiDtSnZYdOS4IyC
PNkO3CW6JzcyZlz/vIP+Zqab2TZH0GEb+6APqJ/bUq8DDAaRtT7mstYYABNWrYgfoEpE++EVOfYH
4NJTqa6jOMxbYFUms253A5NLXS8w6JTA0azkM/KfQG5BDoRgRyOhynE5FpfoShI907GjdTPYLXbV
dn4VrmNrGdfv10ioBsJo3VsbKP9p2HQgW1hrT3yfMZN38OlqpsYCfW/Kyf1l9HOKnIyQqIV1Tqqu
pW1PkVfh14rMnGWJtwvpyrL9PO2gEh5/pnPfhVNFUd2VUqcmxg2rbgTWnO1kmG8Ycrm2KjfaPH00
8d3ijq5yl3RD9HPPcuBKlEW4lVacEbwH812WdJAWnDoyfKB/WJ74ox2Ihv2Q2TaivVtTMMWfDcma
7dopojp5QOwyIuPhnwSnl920KqtqYq9IvTJ+O4Z4iKF1qQ32C+QV6poKAS4/+INaK9AEodJb5SkZ
2NAJYyOGCVUYY1K2ldpwp8qX5CoeE/DUkgaHNJIztHVoAVSbgj2NCe7lZJ9HNQ/0xGyidzHhQZkv
c+Lv4s5Ydvy5RAk1ZFx1EtvlTx9bRPQiaX9gFGBdJorJ9OW5DkV4enL/xPNXbVy8lJai2RM01ORa
NqptkDDhjIMtrGn+ockQvkqKqGO9UDd5QHx/bZPyN23j+ch7NFm8HaOaGPn2DYxYf74H+VctcLCI
fu59q/PiY/87uc/7MfT30rRNIjtHelFu+de9iq9dO7i3WB5+e5EW327obNH0dKC7/mAOCxDVhqVd
GnVQVlwDFc3gJQqujr7iBhDuWzcGS02QP6CPBPmZ1wLc1fHpNxF/ITMyS7bg/z2h2vDso0Tk81jT
+Ph0U9SxtPPPjC7kTfO471qs8NaRXqqfb0LmVfRn/pcpNXSM/HbcOTYiGX9axv1TFeOwzzEm5Sqx
B6Kq5A5zPxUCh+3U8e7tf2Yiu9H3nICQGBhEC6KgwB+CC3la3V/nLdwspVRQhoI+TK0IXVySahOM
dNW/ZsaGhzfYtfvGMND99XvpLZsSJBqrwXEEjCaPLP0WrgSr2CfV0luLOxOghYfZcvoOZ9fIM5dl
8KGwwULMzso+5PvByOA1EKAJppJBPSJL4MMUXfofqnmbqRYhVCMImf7y2LBQY/9NrSh3TjDbtRq2
1OLjn+0xYBrGlcb43LDnvGB4lfESp3rYPEBA5lnmWreYGC1Ef+4frejw+8jOYfKXcPFPR2wBloHv
bC3vvnbZK9Yj5eSeUWqfBqU6WCycaAPqCDX0BOyR1gFjwsGWZdnC8i7sQotMZpVXi5XoIOLk8ESN
bOmkBTqmxuzl1SigmbDldfZizMZd9PmUsvNHXtQPDh9/cWiOYGqiBV7krPnTd6ulzmHNUwMnm+Sd
lyhrtQdRtQQxbXXxeHUjsCCvevM+MIeQZsNnEv2Wj/dIoNsTaPoIoQP1FViL5dlmFDwQy/x87V0p
kAnwam+8HsgbtYLmrv5sGXDJ4OMFPVv+sUy99KKf4jM6EXzlFAnMSIYUpjVvL4OxrslYkOP+1jBg
aTj37nwRN2mMo02Or884YkBupWXQFLFf541IiIM6SYJicZ/SeaCChLf4aaMVSQpJ0o9RWxu9+pc3
YQDFvtcQcSdvIYHMpSl/wJ36KfYQ+HKD25dXJtj5M+VMezv/MaoL0ujZvh7IluhcRAMa14dQS76z
N06ksBzu3LQCa8FCBb5tRKP+6AY9BPm5N/4LTbK3SEpTNo0l3n0FuuLBRiqjCFMti2nI4vn9Ztsk
+vH5r/1zAb6kcCX99XsbPE657DHeDcmn1kxxsBnjlWpWfaMcpkv/KZeEZc4eLMvY3JdWeuzZwTuk
IEoDKFaHtzKNNTgIs65rwzVVwKLiJN7rX8QyWoiq1sDgxfhH6R+zHCpAFDIqyNHKAXyT1QRAA+DZ
OI5FBvgHZPSYAizfm+xH+09JKtlYeeA6QV1JhOxCZ0D8YMsxEfhz6Lz0dZBz2bZ1VmBH4YhABx4u
XgTyGYJQhEZjNuETyRs8feDQEc9nxviWmgvunYYTR864LYsPHvdXIUq/JnOSlfwBuHRWGM47ipOY
B+D5iSAv/Fen2HhkjltL5ISO6KfmYh0eChrbkHDyq0ju8xLBEbodfdWAlsKJYro7VYePVt817TGK
cGbt+KEpesDQlxQ47r9A/nBfdQTpWFPJNoa3iGetqVFM8leKvaLiADsVhwRSB3Z9A7L80I0Mxm+z
sbEbHeOYHjL6Bme/1n50+qRXgfm77SL6War9b+l0P+rVRSr5Rn+wXmE1rxKJevljXXCnW76XssSA
FMSAmflOdF223bhOt8fAFz/M0QxrZoLqZ0jhoyc0vsAXSNjkjifMljNHxM4fOlJXkeqx9UnhwEly
W8qXbAiEiQ7pmrXl/jb+DKOfx+e4Vna3pv1Spkkp++DY8dxnRUK3XXkC9K5KxWuARWCpb3aeVyIp
SYTUMGWTVPfF+qIOXyi03Bf0di++HiDMoHnj9BK9PHsPWURiCWni/x16kkAQwNwDPLDcxcG/K6yk
Qb7bmOK/M7kEIo1mdh8V4cNAXmMXOjSPg+EwV1i0pDbayTlv8lbnuuTuGR8mS7PRXHxNwrrhJHjW
dsryQUL36kukRGPUOOQala2WT0sxAVu8FNCVTTV8IRx5Auyo2lFu1V8lecFo8yia/R9YyyfQZTt2
uUv9X1cd5e9q99SQzLx/DOB8b6OAtc9IJ8fa/l7CIdBHwI53dmsIqf4XJdsVkFsIVvKmafxx3f/D
n9pwXvvYwy3lBc5q3A5fkGTIVLbu5pkQ4f0Gjpx2obmFvFa9ON3K+UQ7sNjynictuS9Geuk3twkJ
uPjbZ6h0xcy99tecWasDRAQTlmuFv12YEwbRfCtwUZqxu06bZJ3mVpFudsbm8/lpccNtubNMmgp6
GMZwc61loB24fMnfFOy0icXj5oEjISBF797M2+40RXU/81VTygby5psxOrI4QvRdUq6hL5J37VRn
Ao5/3Rk29DsLFtdXgVnlsxh31lAh1KJc2pfgyGIJ+AkuhKBgRu0dX9q9Pc4SMmIqYyDQI2PE0lH/
0Oz9RMVdoXyWEAFVuvp3rjGAkzIzkpWQtNJzomieSXcAOeIzxNbHmPI6jKH103RUd7kHGaayqhFp
rJwY4k49rQLVxbr9IFmDrFOcSXZXwuMSiPgIxBLATyBH0DCyBXbzd18F40ejj1JVv4uqYF1ea2pu
4lv+olW8Wqq+JL8dhYvjuap/u4drr6u1mqUrnYas+iRN5qURqE1GkyF4vrAPeYd9b8MK0YyOGm3B
Lb099vW7gkUWmlfTccBAmO5Uc0Y9jQ1YdMOGVOVSmSP9LHZbQ8tmnUYJAJvIGW3IkwHYzGW9zmM0
g+Yj9VNU1C/mCvOXborJGDIXqCemlI1XaCfMmS1nMAmTIKY0BnArsZ1awHAguW7S6wISgWR6mW2d
8VFVai8QHOu7lrusO+c/DzzKt1wdIkqsBZbgQ7uoF1bdUBsBqzHXqIioV5auvVcyn2pC609W+Oc/
omLz5+Qe0Wgj9rFerzsVVx0YN08qss8d2ynAcl2BD0gs7znVpcZEGhUODhINJAK8vVDOAUDGuzlW
sWYSwQitfy5gcZ6O7q0GNtbBVnnsPvZ9N6Q3B414zO90+Z4WLC6EeL4PDfbP4CP7B222y8SYmsIc
1RGaV62dmjR01KAK2ZYueeFtndQ1slrrPAG9wAUpTS+bZJAdoJfy3pjmvro8BriKiJj9NMdwNjGv
+C1WElUuRFU/bTRKclW5JvxlPqTJre75jcExNQL9uAkEQrQV+n29mt2OMma6zmgE2MLTz2/8lFDk
n0CzThuF09xHtmGKd+eI3bl/BaQ1b4+l15ociwUiy/mX8S5XN7DPOvzq6y3SV7HIwvb9DolZ8wd9
R6fGEJjKdt7g582M7hbx7q9NV0ShaCCjf8pJIB+80MHHGH/Ru2msn9Vsnd914z5k01isf6PgwIUd
lIVKCbnHsZggXR3PpzDg6BVoa+uJEq0QHPxGdc5L+fGHpC2mFGMFuTj18y/qAULeRVv8vwPVqN1T
jsffDO1ovaKy6kpuj0EHifkyzfh5XxRoPZ6gZcg2MNoF4pFl39m91aY9JklOEfmYKGDnT6vaTI0D
9MuvxMlc4tjrACg4OXyj+M55L7zrFVzwFy/LEI636lRjQxolOdl1YSW3xF5wOnCF0CO68Kdc/Fqh
2QdJVTEa+UzkROEfMcfO40+Rd2LCc32c1Aa1qSaTJJUmn9gc/0aNxAGpyDwB0Mdqct7mEXWz2jip
EN8aqN3w+K49iLra3tPBqVBHtbfsNWeTvxZ6e4l+tXW13s8XW8Eetof1q4BJf3zAnjUkseW5m6jF
BFn4egW/sm7QyerVEFCVe2MuaYOr//mgDEWRTZArZc6IuUbx7aVU6Rq/3W/bJll2+HCy+w5Zair+
ZE2M/isNgm54YhEvZP5TJWXarOb1WOMbk+1m43xFtBcCTCG0Qx+Ui+6TP5A1nJdvkrqBph6tyxCH
2o3R5tGWbPVpzFOKJACoSxdHyEQ/EdH1DemeXWIrDKCwEGn/v/l5Wi8WXgFfo9acmyFh3HlaN1xQ
t3OGsIOoH6YTZ0YXcZo+LwGGm7TAv83VGyeddAAagxU0b0NT5lrdb7n1GTXLiZhctrMZOH6dYKRS
bplBVDq58L7kPBTvfUfBnMKs8+/UqFGYOdmkdmry0UsNh22YB4eD0SmCCMOnAgjd3W3AlxTdQJsW
0gPbUaRxfenH6X1O3GdP6pCTHRxgtCRt/bJhNPnFv92mR50YccR56EocIItX/H2nkfExPolzEbXH
ZAcdcsLD46We0vgpSIlH2qQr2eKHs0V5Oegj1riyc/0Au5W1+mHPx3yW82gj9BiDgQG94D+Wuv24
jD7dYIBYZvjwdE4GfWdnELBU7psy2hfN9njrDJWAe9BAFv0nRAGGlDUIlOOwkfOcY+YvKuseidvc
nkHm68ymByyN+As3YHX2VRxasV9OWm+viYcHVgRiGdODrDWzy/dbUL2G/XJLRhjrxoVP6mjoHSWV
pFpTSQxGhaDHlQ02rYOdtcGkCLDDVeEsDbYpMt9df+iW3PjgQMavNmiYqFkgno2BkNFbbhPxW9+F
8P766m0Kyg2iAWm9zXxAx14zO/ICjtmFR1zLpELPnuj09T4kCMJVSpB5KKeoq9McOqN0tJni/j7o
GcQhOXVxmnrdieQpls8/GA80l10TYJ1Xsqqb9yOx8i5wADLUqUwBWWJ/6M6RRIaJUZVVFZpjtTsw
yFQdm7l2kMiASaZYpi54xqeJCnavQLaKxxxzBAvlSMF/VLQAMj4Jqsl/XHRVjtjleGhs940qQ7uO
dXSXxf+UbhAHNNRqjqyazUQFyAeVCr1xVRoaswJ/MzztyTu78LZB+9nBtnzus27RZb6d8ZWGCoFG
g+e+I41hyHo4NpBpvyvS53jBA2Qq9IsdvC9WH15zMs3PTlqFUCerQYd3G6lcy+wYqsobyVbGWd1w
f7KIUXop6gWf2S3WCXZKdYVlv88yVr7z+6Rcyjdhj07lg7bVHX+PffiVgPARqrHL40ull9+IO2QH
ryzk0dTt0CBwpzKb6nAFJr6kBjiYM641Q5elt1iVcdsnLkJQ/kFhBJU5T/u3g96sJVLXYaUqsIL/
9IPIY+YeZGyXOVQflEsVokIPneD74xQm/BiJZNxoemEIKF6aA117KpdmzuR0rkF1A/7IGrbzHS5c
WqVjNTG1GYXP2jFL5xDH2tMVVC8j6Kq1YlznxY8+7ydQ+5AX8Zjx4FX8qlKVP1XYXK1CtJ8VsgBP
Z6BtJYiBlSMAVbheRQupS6C88yywS6HrNASOWLuN9PUSqbz0QiL4fFxM010ZnVKnZvZQMwBff0jr
U3OMJ1HEC48/FKLMrKuRQQL7K1RmXNIHvvb9f8LLTS0Wx5ImGx1v5dibUFPRENbJSTet62gYxg7m
QJl6Q0dCIXL6/I73H9nS/y9ieM+xva8EY2hkfu9wLENsn8Oo6DXKwK5x5Gv1zhiZU8esmGkomPOu
6OAbnhfxrARJ/VT5q90FcoVN/l4DlDbniJ6dgNHWjHjg8jHxNl8CyhZgV6LX/74mQHA5PMXrTK70
I8odCt73AoP1BR8JVE5P7P8Dm5hgkxAuOaW0ViRSpcenSeR0zXf3F5nQ0uQSU4M9oqacvabo128N
b6VLcL3uhWmrKJP/+ilXDfej66CBx/rzeK5eIiss9JtZkPLICtY0PK+ASxK/sKUir6SnzRhtoHh+
5OoD/CZjwb3JineP5wL/BKWcFkohdkAnwgZPgP74rAS0KHbW9b0c9CTZfLAhy/Pa7FJI36YchQQD
kEsm08yKsBSLAePC4bQvxlT/w4T9LBaQX0WCBEv0zOcy5jSFm5gF2Gnl4Q65XL53O8vIJHXr1VQ8
mEx1WkXt1DKFjyyQpMuMAE/il9tgPXjPBQhrhqVvt8tfqDKxHOIAqgWmMKEKAFU8VKllyznGwHcN
pwXs0siLl5roOWYZPRpJJeowgTQtp8YICoowR2r0mVEAWtQ5ybO4fY0wIprTzEbEas0N6D0m/+14
Npg3fnO+mJw5hM0e72ZPn/F/6uLXCQ14P+X+rkfs47vrgkKbg8p/dk8TQUwa3wte0++ZD/eLlzPn
orcVUUT7KQV3NStUwcQTujaVi+1zzqhXMSGVdXO+W+9ZnAvqwvDpOWSY08j3xGXBzWMQTdalAScH
Fd6mlykre5gOZMh0ayPmJC8alVkB0dn9UYZ6GlvcC7OtxwfEcb+VcQpVwZrlkafRYO6cYtC0H++J
nSx21D1hChbG/R+iuTVws9RTF3HR7FWimmuUB0eK/MD2ma/sDbXZf+c3tmkqv7Knqx2c5odKGU30
Ku16jZgIfqEgYmBUh4g4YhYKPlZCmc3UjSwQwkOrQkzqv48x4tiRkGCGQ38r9/JGMMxDmqaEB+Zy
Pj5WpA+NZN5ElwQtQijPg5Wma8KDFwiz8mMxkT/4tITE/f88z1bLsFqWIOwOjAo4IoZeAWBknipM
Ter8MSiAKciPZyoeN/KUOxqYh3e8XiCIg/aw6w4lWqMggtEzzF9fSPy5Nr68C+qY2etaHZs+BWTp
MTChGw4DeBAu0owUuKZ4WXchhdNvgaraVn8HvAJbjUKWpiniM4iRvtobFyOAPjizSqBTh3znibq3
YqwShxWf7yxNQxh65t7v1qquigsueruVze38U6Udi8iHmg0IB049kWIPz407VcHwTm/jPEz3Q6Dr
51Ia+BgvKwEVSE7NoNDxn5bba3LQPalfXbXZCeM1NDrQlWdUnq1Y+GaXP9a3ra7CwWxZqF8+dZSH
VDihStkIJ6dwS7ahGkR8w9c+wbLE9gmSGLrY7Wu1mIimkB4B5qDrmvwlxmKZhV+EuH1/Yv+7K68l
1apaDkunb8qTxN9G8s90mHCVdfOwJmetrRI6vmDL7tgU2xu1NAw1rel8IFcpiyHNBZ6RB3l575cY
hOuhO4Jjgeyz2/LsptlfE3LB9wvxyRGKnz9o3hwAa5/Rha3pXG/X0DzUj2OnTetbZOOw2lTwzI+w
2QqcQYM3a5dd3IKTFFHYGj8SL8uxhpxueppNsN4cHTuzI0QAy3Pf8KbhxuUFvdBcSrAyItXi8hNZ
5/i/AO3jtjbDK7tEELR3VfjBLI7d0FnmeGVK8JId7DVVFTybo4kzjK5EAnFmX5FDvcC1Av2qyg0V
z4p4M2C/y0Y1JCsrcg3BPSOcN3AuC+fKNpDU2CHF/56WkF0T4kl4CcprxSNieln4CuN1pvQOWm2g
LTTQ/ZLg+fK3UF1ED1UcAvbAiYsnEa3SEJFFQJFSQgx+eUmkfa6ITTPpprsJWdbdKSZnu+9nLpIZ
VIm/y/HXFfVjf2tlR16FrFSDQ+dR7Fm5X4ut+HEzsdE6ahSD6I857+s7ISSytfZCWTetB2RQUnbI
ldf02P776cjET9nj4FpBKMSczBTzRuikuQHA9QiW/V4ywIr5DqS24v/hDkZ6virowmLCFuGAeVVr
CcyVNILeRMxMipaPFiZ2rm+Ik+E6Mt1f1jHJ0RtOyO8QZFGexllyTUO8QZVjbdG9XU5MDUPZojK2
qop9/GLDqsCzti8ioQkRN2h7k3xboChUBWyDfyM3KVFkIEVz7ac8V/vsiR7owl2KMIhuRNxKdW2d
WMy/htqC44w62CBLXfv9OvSq1+Pazfuy+QiRFkWew07s2liyqnigoiLoHcCOYcsSUs6zBQGjE6+t
4u1pTWnENdZm6BRSilQExyw3hZSie0fcj72V2vAQlOdy3HY9PQM5EZIGu72rJMHVM4xqJMO4fCtG
k+BCGzfGSBZ5M2/WM/GIK/XJiopQjZkiDdFcwTsCCmkPOcQCTpmzArD6aYmkqdu0bhLWigwtv/bz
x3JIozhYFqv6XW42ASpSuAQTjOwUOoNbpdKQ6wxq86QAkoG5c+zdIzVKBPIxOr8aCk5A61mlK4aE
oDQpEgguPzJQ19DoGIhtFhMmEW6yhoTrAdf1bY6Mme5j2rVPcmJ7eTpYjWA27Crw8lbo0pNCll4a
qmRTmXoEzm/B89lHBnO2JYdRd9vD5DK9YBzSVsyP47tRQNwL/NSC8HWtBivuJjgZVJswgsWMPL2a
NIglZB8mU7iK5BzFwKRhGUlv2SKziXByQhbQ/W9MBilc7jYQaR05R6GmBJMHvjR9YxNjp7YqmGtK
6XfuV5qnmEYpwhfPICylaj9vVwun+iuhbIeMSodVD4HnVgM5w3A6FYYZd59LrQp+Z4Hyk7YTT9Id
ThePoyIPuCMqj1KUgvpJ0oHpW6iWrGPpii/mt18/630gRXHvJRVD0/24loXizLMUyDy1CiKD2JMW
RkuyHdQwgQYsHds0Lbr8Ar9FvoG6n9AiZfeP/IuCvs2d31KhSaVnsTlt924ZY0BlzO7C5r8j6mTb
BJevRfluQ8k+Ji2V6EpWRSKKrfU8nLL7eQEKtabpOC9YOpwuPuu+aaxD5t4MGsbGuESyFWDyQ7k3
UtLG038fdQk6uQ2kLGa/5jvltos8irYvsULQUMUL5X1DuwogSgoRRnQilgXYw40cFvg09pd6UYcg
Izp2X7wW9ASktmzgQRw8Uggh8IlOV/BoOx2BftbkBLESnzkp9sULvs81aBrHzaOXxO8yxN3pb6O4
gbQNn/EUdn2IhuB5Pj5gvGCMCFkugJgUjNRGbPg1s/IZF+GvoxKOQ+AvCnx+jlT2P+FBFi+aMHjk
XUkIb8YhMnBc29/YoJiMZJ6ueJmfCgYnJvs3TueXPN5N908b2ocCOL/vRiwqS1Rnuj33zFTl63wA
4ghxTf3khOuvAZeJ/fzPAMcDId3OzeoUE5/nbOV3TiZ7o25rk7wp08iaSIiADYRxKxOkT4GudjDK
RfQ7rwb/18wpEWZoj2oTA8hAvJDwC1cakpwlFS6/8bIidndBb0EjJlIHAO3qdM+SsDjQor+w/ImJ
wAGYQapN67iuTbqj8pOFKp+zdeiz/xfhMI511ACQr38t6ojujMldwaB9x8PcVnvrVAZgoCRCmiKf
zq+NVI9/xBlzHaJMD+y2YZgOvKdkc0rnCVMXxZJ9NcRgKCnnbETi8PCENQqkODxxNG1HAJyHSGKA
+hcox5n2lGhhRdbEn9NbjMeFeZudQ8sHRDT02Gmi/Kml8C5nrrnuMgTCYP0euwN6WIB9DukxMELh
zVQpOTLxHqirm3SpC1A9Wfuc65dcMb6Jwcf9f/E7LEnlhKxv5Xlxu9eXUXPhC3NMac5VTSyH2AZA
YF5vZC4fMZfE3bOAs9BbivEUmi+JG2oEy694Hr5EBQM771TAWdsy5b+X7Iiw4qTX1iWw6QExFv69
Cthpu+kukC8wIl2GkMGRbiVi34EM64ODo4SCpI+8ihADL5WJLXdrBrFROIFRkAXy2jUZglyQKQ2n
V4/VquVHYWfbZm7N2oP1jN9dHoy4lCfNSFSqfRsvt+42Dyb3bPRHIJrYWoWuy/vastIlKwUgPzxp
AAoDxu1DjAkyBF55m9UxahK5T8eKpMO2eRS1A+0SlsfmJEEL6jXsOT15vdxNVxtrqi8Mji+9ACiJ
0LYbv7dHH9HBMCD1YnWaCKmm0BJg7LW/J+evPMzE6vXLejoyr9jJUbvxTKn97+NtbA5zOg/bY5IS
8Fn3HJzXSULZSkctFritX5WEeIBfazVWX4Sj4ZFqAMK1MHNdICpt5Q9fqgusr+uB0uVy1P+rYCRa
kNWbVwyU/tDUVc6Xnci12tPsCIbqpQvSCJY1c13r+qFKjSzEDYDSUUB6itVuHI/TBV01oRKveOTk
QnL5VtaTEvzfZ9IgCPkVB4P7Zn9sFINVu4kJhf371L0buG7cyZU1TNDsv3D01Y9dOdEpQfM533ix
X/8t5VQI34tflGSH1jgsi3ww0iqTnwyDeOaEcs3/cgK3EDF5FGEISoiKhQ6HLUPeQvo8VZa9E0xa
Iy/5UZhSVXmXhqf/2NIIB09SBc0uiH/+EKGejLFetEaeIcaz0sfC8WDxkuh9WrCbrfqEwZbIAiW1
YaNZz+l/lxjhWsQw+SzqloJs+aGag6QR0mD0mlLYzuWiAq/uGxG37kU6rfSX6QOl+eWL6lDgx2qj
RfJJpT//jtY/4i2TGgFod4xY2atmHgc560a/838I5ObOuZQYrlBJJf8xRRR19bE0cmunLEv0IjUG
MqcFej/aZ7z+uP1dFhXV4wC9nC1kj7seXV55rh/GVLvuu5w6mvEp9YMmTcN2S68yWUAOmirGS7WZ
KM1FQ+lERn2BpnfBVu2J4qwIWxZ8+YKdL5ujc2I8T6NwiEOz4GGxbZ3tyew3OtYmAMWGpJJ/U1g6
Gne5GBZDF2h+/sha6O3HZKKFFqTj3ye8XDI90OpFjOaimeiHdqKsSX1yr9LkbWhQYJnKWEs4Rrxx
SluE0jskkkoRJq5rs5+4lif8qNpX+Z/UA4x9spHuDsLKaesZx9yMEco4GwdKo8YF36yxCMeqFwmR
gH8MKEMALY60XCwMkLzBZX5KJDp8FQfYVO2SDuw7uzatMgATG0vNk08dRQlvmaCthacp9FCCp+LL
8MWrHdYfnnfrTfQyszU6fNnOjek0/m9+dE73E+b1SarYYTPlmwpxwSTFYGyJFEg+Y62LV0KlRihK
On9DMVhdJtrlH/r/cnPFsh4Y9Fy+X38/3vMvyNiKvR3NGfEyy683cQrquZe0mOFs4B7nqhpyyLm1
16vYGTSiCrk5EyCr1mAd7ggmsszIKQSnd0/Nr4rlhrVb8IBiSp/UGkaCPN/HlEO7x7yEzsADkjfL
Kp8Gbjej+Mdl+Na0Eie1ghVD7YttdQtJL8Z4/4l9u11BlxBkUrP2qx5OFW2Uiss/tiWRGfb3jphB
jz9K3qUwLHKhqY2BfenxHKfDyT7B5KyckRZ7iaiWQ29bk5yt8hNeRybJRAoPzLqnIApW7HxauhCA
cHysmTxvw/nciaD/MbXCF0nPE4nVfIz2lwj7pF8M4cVQqToq7FPe9GnXTiJwpOh/nehly4b0KUU2
AYSpGb4IcRoSqVW25uOzB9RllJxyWuXIWsula/owOdxYtfSv6JkK8/4gyAHbay8lom1GrFBpIrea
DOKzxLISb3nldlO+0fN4RQ8HV//kD81rg6eOb6cCqw5yCGXb7EHR0eKGqGntVDiFpdO9ZvfYjjB5
USakx418Qg4ERYI2BMeo13SHGalfPJksM8bE5+g6ZMGO3zPS02MUyJKG+5wWnCO1kRQjdZBraiQa
ZbA7oage2RFo7Vc14NL7bh5pGHycZYoO+jX1d/JBUg1+VC5CMbr0wsWJ2c2druYbQQOp4O1XyBL/
9GfisOxqpJi97cH0+rKJ0bx6pGHfQUba66ONYZNiM+jiuuFo7ZhS6o3YSLNYqI+Ed+QRUsghzQk7
KmrOuy5JpmKqg952eks7mYgiGqO1VMKNMuNjTJ3999SlDxUEWed1+S4d8bkZx5D4RZlHYTqjywrH
lu2uxi8+KVqa+Z8t/OaEI5H/kUvzHFaRK7rDePg78+hrHwpUkP1Fon9Qk4vPxIcG6ir/sNlrWYy7
QSxWG1xie4qjHCUwPsAID2joqcAKI+jlCfeSVISc47JeG8Ihh5JFeti1rZJonj9ZfY8KZF6qcz8a
NmJhKERJAqGNe9MRh3JVx4uypDnUfYI6x+/lBiz81+2nwORMKfeLuD6qydn3LEIU/BnNdl5ft0xw
aQFQKxc/ZjoKHPdX4sD+0rWefe1RL6kxII+McjNprQLloTPyol2aquz6D/cbjsTiXS4QpbypGAOX
/OOtuLdbb+GahTyQsAYuNcBtBjXFR/mS9Ka51bm/SW2+lD6tpVIlkPuL/lw1DBwI3BY+fjmXZLDp
XjDJ6xxirzgsY05Hfd0us5zvArvr7y+VzXAUBq0FYTMMLelXNo+VB69kLr6Ic0VSZwvywOf2PQLS
jov+7Q2U/sRXuSn2lWBrty15dDsYLMd3TF6PYBxf12hfNFCjD8LnvQFPJysY9XzVin2lxdNb5WES
lgyBA4/cs0ZBnf9mup+y9AptF2J4FfBDyo2R3Dc4+YZTUPII4KYZ4teZZeOttMODeb/ldmgFUC+L
VKYFASXSmqmWcdnuY+MnUgov5KwbsEXBfun+PwZ6+zBK2U+7isKH0iw14dpctTkmU3RHpKn4hrL2
ZB18IgB5+7Iakqx0uGYv8015LZFT7eWTjX5RLrClP240s0jsb2Rx7W9Btr17JuygZfGHLqFq25Ig
A5sMRQLr0yMoIRGowWIOyl1vE14gE3BNuFfnBpqcsocU0/XqULWRgewcQgT7Bt+jmRY0f44k31uz
hGKCYNCeYA8xOQ5izw4oR1cvfTRqSmqwbOnSUy66aAZG0x0WEQSqukPl122TcYmxv9gB0JVAc7iK
XkZ2zFEZGJL21seN2LkXsEqrrBsdpXawcwV6+qJxy0hbl3/gCIlvs0zUq7pS2WRPSYnRmSqJWkmb
PuJQ5XQuftdb/A4RvChOafY8KpW4dkBSWED4zrG+hR5d0YMqDhYSSpQa2bdr/hNIY2qyQ5q9+b6u
FJ40sHN4HX03fajeR5Rhfq86lUHcn8kfCHaU9qVhqi9oTMw2o48Tcm/n+YmVRgAbdpkHT14/oj4O
mLk5fIVF4iwuiNh8InVwOE8NkNbm5llIhPZNavQ+CtfbNjC9Egs+fB6aO3WAq8sG4zfpBW6n3qbD
HIOx+kazmeRZTNP5i8cLM+flxSC56v2RakQCs1ClcLSQt+Lge3Enx81NlqJG8B0PcjSwLfiIGgb2
YVCEwiu6mj5s2m7WFpwm2FB7IfbVtJFKfa91Ncrur9cVdnPoGp4zv0lJrFZln0gJJO0I3ro87GV1
nJHG6Lmov15SJjt8VliRWP90TL02EQC3bJblGu/iVZ5aX9fAp0398DiaHMdH7KTS6K6gqBXUnp8J
nz6l1Df7f6B6Q0sDdK3pZY9FXoHQ5fvqXskZpk4a0c046sEJxXFO+G1/44Hej9Je5Z8tk6c+B2n1
pMSoiCttv27zVE5NAaBRHe62967ixY2/SbTgl/vi5zrFoBt+o6gRo+yzJtZUi8TX6VTNG22gRAbP
mZTqrQJUb8fKQHN6131ux5kQ5njNN6ckdDtBOOpuWgEAH/fVJjCTraU6L6KCzBoZFEos1zYzPsR9
d8JZXbqSMAL4NRyAuQlQgR6hIR7IqjxRu4zCgDHWEzyCXL034z4Mgk1VHee1XmwqW/XzAzlukNNI
VKricR1L4rts+5UYomP3q2a+1mSMKybm6VvbM8DYD2X8sx6h3aJVwUiBmUsSbPEg9v6GKuG1z47a
xYtxTcFIAIOwSp40weQhmoJNqp3xkD+P9BtFAiV+euiWmzCuLuBzOQDADdJf+VYp0XIkDG1B9aER
w1P5zKwysdMg7cJ5sMLCHwvfYwru3BQ8GzmMC4qqRoBVw4/lCeVtD+dJ2cH2Wa8t63BB5ytPKPt6
pwe/AM5EIB1/eZBU9YlH5bjPnAOJTPsr2mWYQoCIi03x4YDEyYMF+FwtbNxCmJEBog4G8zSg2UnO
P0j/3J7PmcmNZezC9onkNEhUNwK13za7ISuLptBxDNjM7CFA0qPEYe5yLnnHW7d6+AtKDnntuSx9
UuIsIItNP5gjouL99JZZvkZkSu5/MYgrE2zQIzEsXWSfnXW6YT4GS4hidZu+BlmVcrfGAefWdaJq
DvyXtKDb+/KkI8L67wbnak3v6+dyssMm2I3+qAN8+NqEEHi1Aelto762YZRx50WTPpQWPdwd7uzB
Efb2pZqlUjp7TtoV0U7AWVm/GgMSJPitpTTm7/mmPycHmuhLZWNBIiyeiJ+taYmZpPf33R3tJi0L
C57IoWiSAraJCjznJIYEyDGCy92mRnW1ZreoHfPHpl/uZtWpJ9mATw7+nlR45RR6rC0aEilqHFyo
sEI4wP+kFu//9ky7LIXOaYHCQZK91bBkVo28KR+hUDBNkh07F7NavNk7kPlzhCxg5vNFEcTN13lo
xZeo61rF5hLT20rlXc27dEYNuofrqBFxmlsR+PNu/VfsvBowbC8eonQIe5Wa2+KmUarfQeNz4QDw
Hz0fHW6zF0MwHOBf4H5NMEUDZgyLP+2hSZw/Q4oYKVc/dP+XlUK3k3WXwakT3+0CORM204GlRQfc
YBuzLc3hvT3suDm9ByRxn1vegRNrYcVQQ8imisCQtt0tU/W4Ok8fPlgqNLAr36s91bY+AzQ7WQgf
0zWbgXmN2ulYLdfJbmOeFXudDDmCdOkueEoRrMDwLrK2hySro1Cuzs3k88DtZTgHnDmZI+dI3gSM
kE1NKq4s4jA+3Ma6qEzAsO4x+JAygJk0bDrSfr8LTDJZIqTyr0LwK26HPZm2Wbu5IJDg2f94UvCm
GgVSYdVkd0wH5zfc3QPNyceVN0HV5gNXDt1GbEv7RIW7sA6McPh4ei8zI+GkpF6EL1CRZ3m2skV8
89SAnkBUA6mbzzTKx4EtkOcaCoBXk9bXH0/yWQvGKwNlYOYPZYLJ7FWIgZbW5rl/5gA1TZdnO5N6
AkwkAwJfS9h+xg6wdyWV3qQah1pbxDDeIa85ZKhO/T7llK0eN98lzCXVeI0dXhoSYbgiQghx6J0E
xXSowaUYnGAN7kG6n5vBKHU6hbaT0ZyvmTyyUCL/TENTd2KHsmfr9IrrHBL7WoqW3mneWz3pn8z8
gl2QJbAZevXoUsh6Tz2RebSi89Aua+0a7WKimDGHrKVjFm/kRano0Nz6j7/IdmINb8G7/tdaBSKW
EsED8dsPyHYeAhlRHNh0ZZGYQy9ZK5xqcoPAs+dUhAyeCxGtteUhDTYPjRJWsFJBSDdmLGOPtJa5
+XKuUNQZoWOVJnX+6R9waqHUkDrnDcrxNV/0iA1lmAyS7D7otT4PkxeAEz/bXYwykOeKhxjyY501
1YQTx6jp4cEsCIP+RTA5VhnZpqeQfQIfkkuPSJ4/nB3TZnJHYiiip0nhe6WPyrxBINoJ6RQP5d7x
NDXGKODfLHhVLqWeq+eOZvbICVnUWU/JztydgMPmZdj3lUkr1z9uSO+OxU5ktCkUvUUivGr5waA+
1tKtAtsdmB1NHAYsY+rYrui0eJU6gOrQNZf/mCI5LVLwr7otxlI3hR6w8cxbJBS1uAAbUu7VxkAE
F5ZSil5IqrsE3WJWTqEhZqfgyjxFd4v9qNt3imA8rTVlXLm3Kw7HTK30D/uuIxXsTSbs/QuiazJx
/yg6wCYw3lXjINkeqrpoaI78PQ6kE4FcsXuqWUPkcPHX/g/PxxmObLTntrfY41GSV4Zxovf3WUFO
t4UMLDVYihE8OvPUpx97z99swSpl2fzmDzcw5bcsqDaHwXKw4ZM71sG4ZJsIv6MFsg70mObrZYCg
2Gqrp0C9nm+PElQW2VhvbIDfv0rL+XM6VgkRyGKolYaklCFzhGdy9iHa6eamcX5r3is6tk3rmnFt
AH+Hc1G1HjGJdaLHv5rx1GDA6Cpgk/6l3lTIzW6Lnz6pGLXJN9MIeAiAXBajuBESeXGFiM8qGoxP
XGMd/8q19n+UcgzRs3Y8YGy2gshvh85LGbV37THsFuLYyCuOvoTUNGKKW5Epd8Xnpxdo27LKmu4L
2D0renuYHk3Fs222DPYVIDMcIAMSOhduUAmcGwkRing2fqKghzo4yVfrJGlwU6KvH07Y52nehKd9
o0GBi5BGhtk3gX1KzevLDJ0O0WGQJV8Wv76qffhurU7Jb8vmQg62UNK1RccSxE7now2u9vhfthC5
gk4ODOwYlwVmqahaISDj3kbGWchgrIwfCZChRwqrtj0Fy4rw1aCz8yTHDMeLklx7sDoXdaf41rW3
AYqiEG1RcJ87uCClj6BugGTkX4xfm1SRe7+VI8jtLwGCvRLpFlX+Qgdrvhz07AOeNSYLl3bDL8ah
MLcF6PkjqFgbCM0HhewsKRx1ZG7Pu585Qn97fNUpsiTwVeiKvgEVI6X6Lx2t+3KhnVsOXGPvg0yz
pRuLdPmxm1Fz30xMLrK5ZeHUyVBUlTqK/k23WxuGWszpbDUHs1jBQwyP/70KMQ/yZJ9hpg+X+o+L
SBJRjM8UiEO2oGhTxiDbeni5Zkpb/Wte7de4b20ganSNzuDa4F7gnmGzHOpIbbNpEpNfovfxVazN
q4rawnoIU2E9s8JHbnVWH1cyFpVHRTviepzN4NwySOlAPFWa8/s2k5MlPe51c4ebpzc5RT1fw1iu
WrHEDGl2EHb1YRA31mJ9KHx5lBHusy38rW1sjAcjMK5Pg+yDfmO6bHNWDreY1mcYWeArRjxZVEmN
wO9dRbsJW4DP0ac+eIVukNyxxV3p9HUdls17dZjHKb9BcmRZtlww69RLbpQQ/oIbENavXS10gduH
DycvmkLKqYA6p0RAipgvzQ4agzZ7vbhNX1z8ftQw0wE4y8U1Te0lbuhIishhj9BrkP1su9Nwpl9z
Cea7rhiVx3+KNcyfA9M4qIpuxK6vOgPLn+zWajVveg3Ym06U0+4be5jV030drEQv9nOxt8zBsPDM
+9ilhM4dwZ0xcoMe8M2zoacuzFEOvP70Smd+AGVNnjRoex3sLCtipTnIl49VYtGwwhn50wf6kmFI
cAu/7sDM+Ameqn8KiHV9HYC1HIcFdr/omToVwUgfdaSDSR/zOiHW/bShZQBfUCNXUW83HLMiPvfo
4iZ1Xk34MZnq/Ex+ZnNjki6g7rFg+plWOfsbHPJG4k885LTfENQ50PiJM0fLehqoBcelocV4A5St
3HJHbh0zg15lagshrM594o2rmJYxVV9KquIhLz9g8KoE6Am2NbCsQ2Gmczu3EPuU8uWEdg6ETeph
TA5qPdckBBW/fCNF1dLhbyEo7m24qMmbINMdjedlZVd2iurDwymIrPBNG90NOn88kEuYdYpI5WmG
eiWPGRp90fooGdbQDIBB7KYsJa2bz9DS0xKSM/GF4qnyRQ9v0jHVhZQbfJYZvYeQ/u+J/XoypP1K
BTXnQSitgnEQqi6qj6/BRBsAcHdJsrdTEo5MG364Vdk4rBlBv0RnMu10G1GunMKbv50oAhGWmssO
4eq0ikWcUSHMj9ghbCU6Jzi1rHtaLofPkyL+O5DJKC3v7LdGZqOCq8VFu4UNrnHBgNgSgDRa0Xd3
ok2QUvrG8r5p5zSWBqeu8EaKSX7RUOMLL6pVzUrjrWnHSKU5s/Yv1QWmt8G2k8kDhXozzrrgLOPJ
tm808tYj6ahC5aoVqiFo4oHnRYf6c1+CahOGJjXIkTv2ic5lXL6Pb/x8neT5AmRWfraQ+0VQmMtS
QH9QuEsz4/PnIClQcIJsmikY5LGpFEJkc6kX5/gWySueoZU5/uFWpoWok3LGokLH4TaNQCM8ln6p
naQMvmrGQt9e3tHGL2usSRINaEunKvfP/0vk47HS497IaliIMaUHtQK/mIabISeQYADqEN+CAPef
d6wMw9J/oPz1RJCCvrroAHymNONecQt1JqOr8FqIuDEiNbB6vl2nOu0LyFiTDjCd68A07GR5bFw8
7WKtvGgsuWC5jxmaruCpteIWUBRXhFyH5zCseu1MMbmwDVjXCMO+aS/+ILX9T14Emlo/f0OeDboZ
fSQfP1s5Ii4Hzo11zWX9dqkuTWXSsvDKr5JR/jPOX7nAR1qGQ/k7EhVL9rhwlR9/ZDiHBmb974UH
Pr/wPuT4k8e/6caUYqn3a6y2R7Gc1xdFH39E5qpK44N1T9cMKL/txMeDQXX/ll5fUJP9XN6tIyqx
oYFleM+cWKJB2vguXhVil9TaYsQkG9/T4KuXEuZQcsxl2jGL2bDxAsgicXDYlQ5ZuWkJi4davhiY
AK9YH6IULh/CiTUi+fpAG3qEytOHOb38y3boNndEG56GpykU+IgjCkMxAvxeDW9Wxqsa/avQ6m2H
+AUFS9C9AXLvLQN3Bggwcjy9Cz80zRG4nWNVXb1Ie7hyRxtAI6X0S1L5NB5gGZgTo+yuvbQaK2p+
NZum3W1TrEAeCw+wqPP2chdUT7w4dWmVfb1FcWB2Wguq+BxuCOybZQmo0+ItLmWARoXBQ2zgpheQ
Dp9OKz/7XbMlJ1x1qmrSRr9tLjNvovuey64nLzFcMRCDZLw3pYsrWx09PRRxf6x8FLxOI9+i6/JD
jRYonah638z4OYctj8DsAf6Ed/SAzcidKhfe3ngb8aTN9XLGLCVhq43EMC0cauWcdVAvW/MVCKPG
KTRjN11GA68P3t9TBQ57/bXJJyhJ/tH2usETf5btA09pt26Utj/SriyxtlOIUceuE0EoQhxl5idK
iixYBGEx/jrqgsHeL4i+SOeGjdRy3f3BoZBdMhrBiwcx4/pWrr6f9KSn+UPl2QTNaAMBTccl7Gaj
f1Sq14Y3yjjz06W8Ges8LHXZtzWCS/tCPA15LBKsaC45pZVOqSu3m34ozj+vdtm1JWrgfPs/YKqk
H8IYgaQINHtFZ6UBrMB3ARJ2Zqmw+7wn6DzilLklhMXRoXxv6fo725aZfEDohgboItCTqyTNxZHX
/TUoM+eUYDVL7rnvmScOdE1y2Fd7RxDscPEdHpcTKQykhyiFC8TOIwgDL4HJPO53+moVeJdWBlBl
36ZJf3RogOyl2VWCdknq1NwOvdx2e/47MJBVS3636GQPjnUmSV62G4nGl7KZCOtfzrSmf7yqeRit
3tHXYknOx9KfWtU3kxxYFy//CsJPnYmfWT6MBQNDt9koU6JnL1v/Rmp+nKx1q9Q32YE1IJZTsd8P
LKYij2gAO7mV+fGzr3nK8hYie/aCBBGJTDGt7zcNQ64t/OUl4NTpLILoiieg3cDu4ozjn+j+ufm2
3PphP8gRU0Moe8mUNzNRWfPGTpImu59vMch0MlkKxqIfaVaHWTVN/EBDd5CRO+qICy7CfVeOf+S2
mdEMf4G3MCniYhpcM7hqLARBxo2V9G4B8CbTPAGodScmH8aCh+ChPW/sRzmh/u7ECzPHoMTwSJRb
VRJ/PDhsxOPbeW/63BECzENUIJvOSfZrqwj8x0rSX5goTqV8vAjkydjY0Qr2pSp7lqlS50mzC60u
qodfkFEM5M6jtpCHaRMfJM5EZkk85LmPvOFdjXnp7/Q6BbtW/f2Qg2qR6rhVyvYxYAmfkwsusL9H
opRAQ3EmO9wuSGNh+jczNedBy86GYxJcSIixjOGXpa8ubG4OMH+18AhVhVcSGDnISJ1RhFWXQrTt
j2cfo/NzlsrTgGQg02vtyPHe5LbZi+35K9d4uF6rzWayIYDrXBJE0iUR5cD/f7sMOc91bdO6Br5p
Xgw1ybYu3gybX3+/Sh3NLfFSGt3gTH2y7FcuWYTlrgUIGxTe+lIlqxVhvSsQ6dFN2qc1jyadZfM1
ZehHEKIRN7mtZ+Hqf3IvMkdSAIjcOo8MsepOxRY5Zt49vXWmuU+nDeDzaD18bP0OaYktrmRUUx5t
abRbwZrU8OuTkgUCNlNlN+L7t1IZy33iPnjr7cSuFzOb3bCGZ/DXRTyXDrSnwZl8FlJ5nj2Uw3jW
KxsCyapmipPOagm/o/MBGXKlYHJSWBJCxPkg8QNrIAluSKBof4IDsunZ1vVZlj4bJlGJzt91SuJw
3Up4nEQAhkZJOpfqop/5nI0Dl6IA8gsKgz6QjNOELQ3KujLb73M7Fw4Sk6VKFZqSQ5oSlAifTLad
g7nqOPgzSG9oOT0a6+3h2N/g8o1b9tZCHVJr7Y4QzqKCl8LaOZHekMd6pZ4hfo3+1WrVDIHKij3X
i820tGOllpC2aKRf/Ij96UN2U73nO09aIn3Zj9EDRoGErsdCwmZBMWvwKWyYebeXAFGovcay0qLT
Nx5JLZ5mp52mVEfri7zfRSB5NDvb0rWi0ZipYBlQB0BPRxEU9qe5AfjQ2I8otKumDKegCdCLsCOG
YCpq5DKkcTY/rZhBWEU79SNknaPBX9BRhLl4U5IiZMTsYoUCsyJ7M8aHFLiGj2ebVSvTJvFgSGrp
EcVnTzZv+Wc9XUhSB+R5WKn9eP9u0bJm6XMsNEf2Luli+gWNqowWbEhFg3RC8AlNPUaAg5ZmwqwO
JQ7NBgVp+qQW7tbD4jBxwOfnkuMuDMJdNqI94Ry1sHTimRon5yFVRrVIfRtqZh627WdMWIYjVKtX
WOg+PZ+r+irPysJt1MnHYM5kyvIiPzcJ8F9uU+rveHq9dpTFVykY//ulgJiozCeFfW1HnGGXJiPL
n4LkMQpvoqjLjJlKAaNmsHw4jgQJsp5OpzxbtdFsurOOPBtTzQ3irkA5qSTRhFO+XA2ZPaVgTSLU
a6hY09QdYRLcydOySc9nW5EC+3A69acnpOd2dp3Ca40CIe72fKoQanv5or6NFZ1bzm8lMHQKTL+b
yc1ZOaLpKzono7abHgHgz2PwbVIcPJhlQndlniq3nsBiyu0zDRvxSQZTJWO10F83XnPWAsZsCmIA
e0jbltBcVM1rQTiT+cGoTYODlgo4GQvbCoMxY+Zvr9Oh5h37e8l7kCxJpxfCQ+HFr+tWc4Ojw7bL
n5x0HTY2s9aFUUuPTGWh83utwYbzYLh72ODM0OaqHe6LFCcZ+MelOBlAmJcfJRkmi4/cP5BKK4Lt
oByVH7AXSDlrfkHig1y/oktx3JZixU4phtD3aGR8pPry/EZemD7pJyfpPX0wSfXBQRjq3hEIIwic
m5ijlYZYGNkpqJ2nqTcHX5N/AZlEjBu/jfOQ+xp7P7H7OQQEgaFUWRYhN829+wAIDOzr5ToGZDs5
pY/oLJz9HKIrt6OWhQ4c28sqpwNQK3uevMYQEeAPLcfybxSFussffXqvGoQYdgfR+THQu0PsuP8P
uDQvJgNwlxPLD4u+I63kqSy8kYfEJePQFqa5lVgZyzz/JZ/gVIi1m3NZJtK3yn5stRK15Br94552
bfjyHTwzWuNvzZzyidAS5F5jUEusYrL7S35F/0X0JX4mh8p1gpOdPD8Uh4obPiWc1Uwr6BrGgJu5
Rzj5J4DofE7GtAjxuCW3eKTEWV9NDg2XW00CSvv6lRdm+expaK0rGn3CLUoLegKgkaoAHyYYxFZx
0CgdU/ARwUYPACip/8KJPcJ1B+97C8J2uTnoKROqwN2pL20YmRjXhPAqOballGbmMWLhy7wSTpmJ
IINpk2xW2xB90oW4U3I8XCUDV3FFuGZVm2+XLSYjktFaSqDP/00TWA2CHcc6NGqXv43TOB48qQgN
mMOk4TVk3tRsK5f4FXTfQRmufTZVqVuv64yco4DcVeC1HqVP1hL+CkVcz4gQHtM7u80Kkw2i/xbI
OQlPGhg9mfQej2IbIbHfuBY/eMzeLGE5O+tetSN7g+yR1+X1Ni63Gl5nw+x6xcLSjBUBdZI5WJJ4
Jp/go+7cb1wiNSPK6vTxl+gV5IuCAdxh818YJ6S0gMfdWyBC1u6TZtbeU1cPTcNLO7VP3lUk5/Wy
wUglpcp665Cji6MlVZgKM1tGWDCzjSOKmwCMd7iAYXt+Th28Fjctfqtge8Cuvsf7km7hAFOhRitk
OMMrpYTwo3XrrPmLJ0jwhbqy0AwUKZ/OwR64luAnx2vRKZUpxbHwmpiFepKZvXb+GrYpxlrh2lSu
XHjWHGrLAOwuG+97ARiY197bDCzietFNeGzvxP59v3qYq0aq5VEjWFK76NHheFVcrwWlIJ4f2Opi
yluI89zfTRCrLiNJqLIt0vSTkG5YmOy8JIkr2isnBFgtxk9QuUqzzART0VYRGiR45ZJD+LlK2XGF
fC9ZdRIvPbyzhYj1+q+pSoqdkAHgmiMTMzx4qBWNNhj0DbiSlCfnI4A++zAa3c6JDJo6yBJJdFUb
sJB8msBuBwXyJtUt9hyQH2gu08q5PYy8H54blJsfcpf5YE6VjrO55sKEL7vaw+JFHous3Rvtq3D2
1cmQzxUa0qOPCQTwu4DpyBSHkKqOUUKCcP5vI3kxJL6/ANY934AzIe7yw5gHo8Qej8ZQZMB0LbbG
8+qiRp+Y9gboDlAg/sMTlStpmehCLAT/hMIXVGb+9x4cSnDvtn6n8Fc3l0SItyqKMzsq27p4KJfN
rsctMjIsTyFVw1D/PnnptKujMbyYrOhlOmloNi2Gep66ovQ9dudGP5QE8MX0/cc9firIlXfX/fPk
9UV8KvkI9NAeTjMinc9ZZS7bCXGHc0oVmuE29AfiORzMbwVektYbUrYJtiIbLblZFiTpyqQyHQhW
r3LvTyxIEGvM5ZqqBpmjisBRItw05j9MFx2WkfMAp2lwNut/7CZZIp82UcOQiryIKd4IGxnkD2q4
Es7fq0aV6Tp1Hw9wsPYJSWEjjdcNOtGNJyAXR4q1ZJtGzSUFcE6dgglLCLVvcGsdbdWeA8afl0l3
wjGAHtDjgcfuwbUMve0ewCjz0gq2SzF2bMmZrXXrPJ1iMHSrPQp2XOD0tCl3n2EJti0XbHIzGCDp
tb+9iBC85CWYOH0rbOL+G0azEnsXcroSXuXLlr1jd3t6Un3vcSc3hgVckMCtCwX33RkveT6UslVa
HebGjptwp9keVfJV/kCCReUX4E1Yi2MjG5t4HzC/RzJdpP4ED/IIlkqx+odtZ+KVUB2FH1/dEcEd
QwT14mAj0ZmbMusEf4zaSVeD5LAy671pwgokajljrD9gnEOVStPZ1sC9evZC6g8x5j3Uhtu4ughd
cV5xoHPzeogcqjXJpVzx4Eerucb7Ckyj5v9zELe+FTWPjrIQGWQc/HHKn2rFufptcbReknMEUPhT
7xyobG9CoIBwLOg/G2vf0MMVngIyDD9KwVkHgJBNpiBbsrBwC01CJP2SZHAbGWsFRIAEl3axlqo9
5pymzJyWM2in+S2qEUACXTDp03kzFYgQKafdqtnBTDze66Lnysrsn1oNPUdizyvZQJndWffPMP2h
MXpcAwAmKstQMSjVUCVAlP1TsEBNlg8Z6TBdhUU9+3X5ZO6TzWv/I7L+mUTzthfF46PCkNj9uR5P
zvok9e8dXijVbbEPAjuw3jXeZ9TvnIGgySgj/D2n9YArwfTG9LZ/Mp+yERd8H9vx07eq2+VkEHBt
82KY+HdQrjVp6I3IiT3wRe15zOQQyb4BorQ3cPojZl0eXo751yTpJhEHdAS6Wc5WNxOBWNLZP4mz
bfgaDeEBdMiqxJVwGkqvUVjYIA+rR8i/gVe1KwDWi/8MobgBigHi8/s1jT9mn0at1BXlZvPiZdsb
f9yFcCeoRnFwJrCw+FP9LJECtgy2a1C92qCMTRe597mMXOKc10/TvT8ujaQCPd5xNMJdIkCyUbMW
U50XWJ1A3xNZL72+gUl64ZbVIWrkgEEWX0KZH4QG8NCxKGJfVqCIbH4jquTxn0bpGWIn1HwHu1t4
fCZNm9ntPqPag8UCc/VxRPnXX4aD+BVoaXvPTPsBqo6o3igaBr2ssy0W0PSGwLM7V2pYo6QVFKYL
UkTrqYJy8uT/p6cEUrES2UT9Ph7maOJMTWBELw/k+s0RcMB9eaHl1MFZRffGA9VMwEs6kIlhayep
PXMUbfShxi7NfITMEFSpMZ1t3fbRPaRgeBJ9v+/2zRQVQ4tr61TtpEaJgyLHneBErq6lk/xlIAOO
4reB1NZZNXPuOEHdNtVLRovd8unXluyvDh8eSQTbEVvw33iB2Y2dk58PneeY9phTfu+BouE3omcG
1Nz27vnLud3tezWNy54GwsCgxW+4l/gAjNhFka42JvaGyB/OmtPqlsLWp76hwi4yFrJnQWnGNRTV
Jmz45KfkaOlelRI1SDPnVGqgApW4kJGioni+LsyZSzPfJT8zLmpLJtaCUYR8vYnZNToX3DXbgL6B
HMtMbf4sA2ky59IUIEUBXVZOzalOicJOcNHuTh5bEUFkUnhrI4czMdVNwqgIkGiLBsErgrxzENZW
uKfe8s+4UomyTyf5qk72qHdG4ofkoIBjNpXewAf4rDrGQgAU0DBYFpr7r7BB9VhHhMhFRO/p6ji8
dpDRd+Tg7CxEtz7BH+pFG1oBcVh3eVjBni46LX9f8mNDXKkv+IgMu7gcXVurQvpQOw2HInoC5WGL
GguIgDqysSMMnT6B+LjTbpAZmKfZZZA6Dmg+L1aoKocsplnjrNrgaxeo2aflNLdQljCL2wJ4V0Kr
e4KLQ9tCZE58d14PCGh4LwS80ged8FuZGYiYdQlS4FI9eeS+Zwj2fiduvnFAO34xhNknVFkR9Otm
elkj32tJA9O5l1h5ZHGArfOsouM7r4GHYsM6q7bbi+Sg73/4RTrLitb1w5WafSk2kNhSZ/sTvst8
zMh3IaajfwYh1o+Ugg6f61vPqtktpZ6h2xptQpjFA9nk1ZrIrCer+YW1ZNi4luf6+kVxre4OwMRP
1/d8ShJvs4YCfq2WWeGIYHkplkg3dcUl1ioIin7a0Qsccs3PT4meFKC/I9o6xoYO2zSs8AzbqrFl
9k8DxR+5Y7tRbKUEmjuzPnpqG8SJmNJlHiTA8l5GQd2onyIK/B01xRKCKcIURPYoO+CXXYJFSVWo
UaBtXzHZOw+5vWwD63jS0YXq3SNODKWFeZ5jHW+dNeT5iPQfPUhyiEZnxPFYTVNiWFZZl48QQRb+
A5dSCKzyS89EDg24C6C3mwaRU5l09UWXG28Sh/xEJ4YcId+9F0Dydy1Rj4xzhxzHv/K8WuqdiAWR
3Q9YLEMzIu4uIjpzybSJqYPtpYL5TW9vNo2CPNonHpUVaQ6oAkBKLttFcKs5XoX7DaJBl8o3Z6aK
pA2ugRPcL0mEKE2f7tY7rwBg0aMgNKWB07ZvtxUOWo9HkNAP8ELvOe8Gw1wFw3zqnGt6pHKHrMSE
pc9b/Zd3tslMpb1e4CR9dDBgld9lotWja7JoCY59lW4S2BkWWTWwqwmDpVzsZeJJtuCBTgXoOHFv
ViXg7/9BAUVofYQqhe3yzOIOZHWMNMrQUyHnBFATaPn6NzF0hdk7vu8vz1aNSPJkq9Byd5Byivvx
ugzK5OZvrJwwbnK/uQtkxvOGryVD0wkKoH9RPJS/xIfhWYkFb0VJ5kXOkk8UEH2qG2hT7t9rttcQ
UDqDiJo0QimilKB4rTaVwijckZLVSLSdGg8r8UBp/BqUP97rts5lG7pzXjjJN0Xoygyhna+m7LO/
hGetrk4K4x3P7N1vpeDd36fUcY4PKtj5cnPnzaEsQsI7xXeUTVI9Zhfdl7bYoFDC9wRSm59pi1GZ
uZ+JHETRceG8wrZVlo5YGkLBdvLeEw9aVf5meB0jjQQODTQnCJrdTXAb+7XSi7imD6qjhP3KTiKv
TTNeLG47dqmAJ1cUHLLwCbpfKuOTUdYpcUx11gZcfc4QXImdykyXJpvp82qLLCBQlGLCNW3lTegm
O6ZdIWUnuQ3sYKj0DYAhVQEy4K7g91m0VSHQ8grL3v9RwrwWjTfQbgSoCcZDyYIO82bDpgLumNpy
K+Y4tllOCCrhck3d+3tyrgIxeaZJbCzFzHU8fkXTRq7cPTY3yps32bDciUFq8GT7xVjUh8zf6sTx
fIrGht98wil02f7knlXcUxu3trmpB2C00yiNwEJnt1hY2E5UKieGY5RtPrFt9Ixwj+u4yj1bgFBG
YrKv8H1/MeMjVEmi+Y06mnGgUy6yTP8PZV+QNmU5AsxOVqSMjB9KaAHTswWOV1SbkdstNB+GNlxE
i7KpEZJz9msl00bO50ec2172xD0X4crWMGr5KKULpGyWNceibeu5Pew1UjWTojxMQsiNo3X/okfP
Qe+6SmmYIqFzhfeq0KKK3sMMgH8cp9m146i3hG+YjKK9ZgnTlX3JW1DToaMWi0+mwnObWeqtN+zN
J6oqujOme/rLFDXUrTzVPdD9cjD+tHrQOyBVhQCeKiuK4dGjU7125iWOrcFhxwFIAg5IRRElTrwR
nxpA0tjIultoZNysfIkPLVLYNnsivajVNfCWD6bKHwRpyodT6IJRObM+VaeC5K9udSf5BvOTxp+O
QDNmYpusCWxM8/9gJc4x5N8h2oiv/1/kDmEhp2SZ0o+90sHht+1guVBmx7XYB5iksfsl2LsI2LLL
K5FYOKhVaQyaBP4MLt/Ow21WDtelj94WQ3lhw/74H5q90hUodsccBBr/faGIuVRaP/pU8Pa43y9Z
kuAd2fanbqNrfvGJh8sQEi+nl6erC7W+825TxtEx/Ic8kRXO3TEfr41lpCKAzjxdAAQAev/hQPAL
tR7n48ed1Xqqss1NPIGpbmLgLcoa93e5DbJvzP4gTLrPmZi0s9CV1PmJ6nhNX5lzpC5/bx1Xq/+8
QkNFmAf1cwc2MvfExf4UmXN1PKcRr5nDZvfVCUBRN2aRJJ2uxcoQQsIXPtNLbrCG9ccjQpauQvsf
xbgSDw0pBv8SnxIzeIDB5NzureE4co+7LoBFMXbZeUE3UhpV9PHhxZdL+d2iz0CihpB7Y2EwLQhq
oQO+uAZ7SbYDZAcjKdlsMHWjhTmcRTm3Q1XXCmyncJJGyfDnU/yPIxwfUA6TCr1M2wyhQIAKVAvJ
yeuLpaXzQOLmq8zDzccmHFyqbgrsazoNh/xZXv8gZWMAq6xrvojg9B7/WXtn8cF5VmR4tIaq1bzR
n0+ksICuC3oFec5l38w92UvIFYF0NLGlaRfkNOTvlAFxgUKr9ehZj3xZ/LLYmi57UNEAmeEHZf2e
b0W8hCYiFAGROmIlO+Hbzh0GlNgb3dbNbdetPXr6njxwa4aGqQyOTaXP9UPsVJQanp2PWqephx0L
DE+ttKF6TV6bS1ONCiV29AcefvDUDfhfiv4LbfoTEtPZk/pL9v/ufmoM5RAAfJpO3XEasQvG992t
Lf2AGVbRfATkdQjrNalCF5G2XhWk8rB26mgIF72bdzlewYtwGsH68v4BIRc2nYBAbtzDPq3SFYgP
yI0sReghAOev+sbdJ9HkDlvt0zXFh5Ln7Ah+r+Zka9juy9bCz5v0wOgHQZTacAjpcyqhR3fd391s
eNxrCvAm3/6TvjQOLZhNC0kNk/6P2KTRIxcEMEajtuppLJCiHwiNwjqS9tPTLns6uTuItYiWiQ+n
QiwomEKnkr0yfvOQ4MUwWfSIQzpJymu5RSD1+wa6iwrgOZ9/WTZbi87uXMV63ytBS2zqlXdEoZV7
Qzv8Ay7Gb04Xk4oA1FBRQn+hq8J+HoOdXqrkcF3ZqlF7f8tDwwJDhbQLgiUaMlRfq8e1azOU44Az
CeUjN91tm04+vqkMTeRiq2ithdNk55jFhtNuSLGHq30rkZqJrjKz+2Gw3rTQ8NaB7gtvxRRd6cSG
Y5D5Qto5CkzsYnjxxjuHulUIi3Asknf9JKxgCdq5AprJEFyfls1bZw3x38OqYcfsr3r4EykyS3AJ
sI1a9jNDeBRGq0evBtAQNDujNPUGN69YzZmChZiH47SU69yWwpnydkVfQ2iSxnLwbX3t3eJihf/T
fkROVFBICKpzQ1cOaKGWt1PtA+KIVzwTRd18SBubO9x5ujiGK2ighA+kc0PoG2nzyy2NJl8ZI4v6
ck7rE/rc+MDZdqFwejKxGOr/bvN1OjVJZjfiKw/Mv6MLCRlZIoFYwhS/hQKYwTgjLh9nBFdjsLqU
qvmZ/jXKHU2ZKjaz6pV6izc9IATHmpuvya7BBTxpPFFs9pZoHjEaQLmLJ++JM8srQenXJRn1dn1/
JQnKxrm0aPgiKxwBYcRbWwAilzD37CRbzxtbdThmsyogRJ3HDDXnxryq4QesrpFQogp4fmh6eM/8
V3mIKlwp7YJO5NPsWEXcHybL0nJJu45TlUCthgh1t2CPGisKAJm+YFigmBIUuIVTkDNTtLi8Fyfn
tWp4fCxxS+0+YE7jHYd6GnuTa/vxfaFX5TzYsOHmzVbiTWhDb99hoJ1VhLJzZXSzjDJMT3mRK9Hc
GsHTgpH9T7BBeNGBL+zv10iSkHKJWMwLXNrM37nu1tEzgW+hgKagKaK/QavPiLz4rJq5H3HyMt4k
5BbIJ7uV1kES6RwPRgC9+hPnXg2V++7auLLEYD2pINLnL6IERjTWszkArzkhvmyMrjRDeC8Z0ipp
uhciCqU3IlKDx78vuO5tReGsKBRPv1gPThhBFQkBLLKidPNyMCVfmCMK1VmE0xqfOv7qqz5rDpw5
mS6DXw48v/aH7V44TfoyJ7elIKHB5ZOavu6IRzYeXi+6EwMw0MM4peKse8FXHJHgq8Xn6OtzFt92
XzIxpmIWMF4rZDsRuJem/p8EIaWbj/5YcD5fBQBUclYuMs6O0W64Aeqp2C+ZoZAMHw3oHOpdl0wn
hbGRJhovtgTfjVTHNATlDB+y6tanRq5tOQaqPZzeJEoeV0SnXUzLI7vbE5HzgnNjbNxfbQRX+ZZ1
vYAc0fx1SX2zeor49njoMzJTeHDQZ8ZBD0sKx8ppx6wXUuaOyVZamyeppTEgEBbUuIasyp7QD08R
DVkODINf3Am0SqaG3fWnjNc/1dS8d+/R1ggWZjdG/sCgxiqoRSXWXqO3ZWjssGVW8G/872LzAYMh
FyI/QcDx4gSRDtoOui4X6m3GxY0sHq5NGyLxPHgTAQVXzeUCvExqIbRjPOMv4G3bHOM2tpMSfnLJ
tRBVPeYbCunY6XfZbiqoEvv1B/mOf65rw+Cy4myy/xBVK2aYzSBryDss3PxOJJWyYhpr1prw/cyp
75xo+Mzdt0h0Z3vLN6OXVPZw817jG04t4icVy54/XGV4mkPFZcHoY/9ANm6WdBPwx2oO/p9IWx2Z
U2K0CFbh3Z6UITvALLS0Kv3b7BjU0g2zFMJSSZw3ddSpquRT4KmG9ESd3YrnRA4MbqMnSj3a/lPx
bJ1JMlbZ9ChxtTle4N5TBeGbactbiYjb1lkiQBGSINYi2ZgFS7IcAoHMAzdSmDbCkO5aw3Pz82ru
AmxOzrY0qYUaHh/eUl3wQ4jjNYDwMd2ow8puSG7eYSryEYYhUCDqe9jsxKFY+AS3KzS1mwxCWPbs
Pt3uLrCZDTsweWtjfol5Nob+aG7xYyW5zHSYawn0ZYCywE8sk87s3eBUNhCCdBQU4MqYW6u1KeTD
9DZgFjlZE7YUDw0eTZKjk5Pc0cYfIhUVQBJUmYKb2bnL8JpDTAYko+tiARCUviXtf2xIpUDU06Jz
6qVyKobn+RWwKJjwRebWSDYrJyKQO/5KpUO+S+jT92Yoyx0aZspYcsvqoYqZNNMhT4G7eUwJq51M
khSd0r+yvO+RcfCrJMSRshXwxdZwq/ZCg2PdfLPZa6b6vCwpfnttz0oc6E53LGhkFcEsoUVy+/8f
9J9dewxvwgKBmiG++rckwWvgVxlQfQ1eQp9yiUBmIBh9GOFxChBYhRw4AdOMjF0GsQK48t5Inha2
j1zo/UHCzIs76wI51zgEeyCTuPMd4aK3GyTN77ZRQSv95YvXnEJrCxKFRpR7Lw7CgFHx4EvrwyK6
9BohutFGIpvEhGedhAaZnTdqlvyvznrqkuwkmHnMfVyWmYXrUhxYHkdTilVEO8uoII+uAbyAlAt1
wvBRQCcdu72jmNb+opKm6m72IrTUcTlpDEBgdmaO6obUyCeeFOUr3tCJqOpmYB31r822jyj7nCby
NRZBHfUioDFqN/1gIBGN5OfiugunYSWXf6hWhMckmOvHs7bcqqyZ2S7QcIxv5xq3CyxM+3+NFBn7
YcJEXyK6cbgZT/DaKmIUif6nLll6kqXcQEutAvnAECDXGi/D8Fuztn91d0m8N77LSHCRHTWxLzoz
D2FEaz0xOXX7blhdfhshUdlci7d/p9lLWtWFLiq4BDSz3QuaEExstFDSDQTyPxzsDoEgUBYZ61o5
wPP4Zka1qd7pRPfcAfR4a1foqN9Z8mhGbj4oGQ8yrAOq2JsQj1cCstl/NxAxoc1MDmCuXuGz0PSA
J0hU+SN5T6QE62tLiRb+gwxY+x99agbtRPf1VrclcR24yYPTpIDYI8EijrOO0Ihbc1BkLvYHwNYD
zzKGzA8uu/WPnRKkoVH3gF7K3w/tXImo/Pj7Dq3ps/ik8COdvItFIKu9X9aOVASHm2vpIqj8tRFK
9X9AKNIZnolmsRZwyPYYHi96bB4yIz6rgyqUmKTmRiRen9U6DfHE4HsszIjoiAoDijA+7IVhapU4
ySJAacs+2YkDSu0Q+dsoTpcwCzJSK/UQvc5ZbLzeJB8zg4WqTJU+LX0zqP4th/NJS9obbJCWZ5rT
mQsW3FzgdOo/yBvhS6WXLwUi4buda2ghW2CEECUCLO9WOTtqwqM//jxIXNGYB0CValE7cgI/kMaF
Pt/rgh0NvXcfr9wxkKZYwjfZ1gYcKDL+c/Po6Nlft0HpIcekToiOwOVt783NnGTNlmCN1g6+k7vX
lZ9WIMgSZbVgEdra2ADyA7+NrNVlsa3zqLoZNYCssuPeGjxu5cFH5JWICxYEIYma/WyHazr2JXx8
qHpNt1ZgfVMKpcXA+tYLw/DTJrJz5ssexyjvYOP405sC4qPtgRZa6UnlJL1qxhroPYtgk5usjsK+
PpfUvDEtT/QV5asQMZBYOSvZEtPAML5IJzT3MfeVlXReCSUlfDhoBRgJOoS1wBIrrMrnNUNpgl/L
UmdalU2lP1wIU1bdvIkh6A5l2URBB4I4vdcfOwq+bCgVUZlxxaQQHeg1v4NVCg3IzHP/S4pA/Efs
W5JklgL2L7y/998jrgZfJthZ7VWjkzLB/uza1ImDg0BPV7D3RJ0LKLgE99O6AOCfZPSOHLoMYiFH
guLKbFuznCeTU9lVMKAgXoU2U8cRSmTBYaFM5SKGGHwcblEPJKpm2JgqPLMO4mpm0yng4jAXzwJ6
m3+Fa4+MveVQdT2LXHWs8n8YW4uArtbkuDJkZrVkacutBi+TY8OzsbS1xpGmvafmf1oU3MINmn6v
2TxIm39amDnR2LbjLTGO0/Fh/piH736X3g37euWBbqyT/iRCaIxFZU7wpYZXcFs32sFD0oahtCN7
ucmEaY2k1jt44rKNurtV1iEZ0qiHSQ6GYvBp2FNVthl6Z0WWMxGeBjA8pfnXk7B9vJ08AvFub8S2
O5SrBU2Rg4KeIyMpI6WCKzVNvPm8L9kZiZgrt9IYTaxpo9IWvHQqPRhHlZAARXguZR4CrZDWsXks
FgruOr6RYqCyKU+lY47zBeB+/EvomdL0UsIpC3E8ThNSKUZXY2RGvH1kJtLtNDcBoBhL6txImA7B
saLu8EctsTKhnWumN/sAOC8A4V2XrWZX7oTsC0cGbQFtVmOwYQBfIqsqwJIIDnn4UoOXUhqvd5Bf
6FNU1rMVMF6WysOSFrJh0/ygl0iAID+bcImO5k/ZIiyxLV1p5x+aoEkCre2Bh9IB8Zhf41tVgeJx
J8/rPpr9VJI0yWgMCXeljRrl9ThnjRWzRlOcn4f4sq0hV6+sV//icRTvw3xLJ4LgsqCFcVkHDL/Q
G98SA5w0QZ3Pwib3eaIbCNFsCL5SyZdjIBYrX0aQFImBDulTj4FVMNCKY0ZL6GcpNfp4oEByWs8G
kH+ePm0XA2YNm7oByDKW1IvGGYsfs8U6WtrFZ1XkIG5BX9mW3XLctYB7f0/HUpG6mwAP7NEj/wSo
PRs/O+5PbX/eZQSa/jbYZ3p/4zSkyNpa5SNfnWkcrRSH+ZFcMh/aVWUJ6ub1hdagQft+Nhh0jH7T
ntqPpc/yvbjygYSZNhLGVYRwxB/DY3UY3EacdaFQ4W8cTNQK3tajyEtZI26R+ayWrBErORflBOZA
XLgTUUMSySyDHVGSpsnBxTCNTJHl1TfmFQX86+hcRf46rgVpzfe4P8P1uRO3PSjN/d9Gj9l2rS0k
PQRoa++sFn9+I/GR/996XzshVHbSfv+pGN+Fud7bt6RQBfE34OFtp9660EP6X2ehZf9KcvnBAr1o
utgw8+G31QCTzFnB5O2uvpuihrq2RebmAznGCfIwFmhUAow377JJvuWB06pld7tKDdfpp7zHItYR
CsOK2WRcanLLCah7ok1JBxpDNnLm8qkoLF9xYHVwulYv1SjQ+unMwEEUvxwSsXERyUljI3uaulOh
Xkuf9O1m+wUR7lAhJblmQmS3b9gscCFw73q7INnBS3GT62y+o5wkyBGvzfc1LfbcwuPCwg+1qAxQ
S8RBYRgPE6HR3bt0BAHzL+ALS6OBXOY0KQ1QEAW+jgTzZvoRxbcNS1RJ9n+qiRLswFyv+ipMIiW7
OlHdBsbj+/tpLvAMFnjtJ43yvTXdtXcBSEDt1+cW00VwPC5beBMPfZkG1Te+yjR3rEeDqnUYy/6d
ds43fFf52GPZEdfqJS139nCHZuWKQI3tBp02+6Fuk9ydHw1UixK9cA7k00f6gS6fvTjzYj23nbke
MhxEhGJ3PhIWIsP8T96JECfg7s05d9yEIeVlgfdquXR7vrhmS6gD3e/tbzhH4VxXYMwXRdszhp1U
f0MhHPoMfQKiKbQ45fa12nDbQaf8Exs5/jAXJXSUy5PTCZRUVDCNbbbP9mrro5b/mpQ6m6y0O5VO
70a9ZHfCbOrbe/16LXnAkyzX6Z3jCKLEia7A+DyKfBGYlTu4BSGotiRisp0bynP7qYJQ5AfxH/6R
WBgd996J0eqy5Qs89/k4oTUv3WZAJGA5rQxIyzG0GfO63m6GnMM5DRyG285H1WJoBNUvumdSfCXJ
Ikqgf0bQu75NxH+SO2QNW4Z3T4pzWlP2gJN3VuhXT8cx5wlwLtm+D+X+IrPnndDtg8sJ1gaAK+BP
QMJpXBk8D3WLPkFYePFxYBaSR/E+xaBuW7XRWUzV/VfHbha4XrV6NvrKOuFxnNm5v3ZgmVV5EtNz
c2LKlHPcwVt8TGPwLsI9hoy9TPVe27+IGAtZgVjO1fyXpJ1OWTiBdkmPDzegeArVw5vbezWWVH/8
PR1JmEswgucU48Vui6rOPJA+UZV0K1Xritx5CEe5zbD3HKkVYNUSdc/S/5ptCAH1GreDReTVlCF0
pW5iT7vEqsjHq4jo2Wacgb8+yf4mSAamLP38GunMDpzLDmSX253+PzzS1l+aCHi/pC9QibQhmqNO
oUu0OcQQTkReYvPSxNz8kNEUv0vUQxfjBhCZLeJ2PBGoAaVUqy1S9ghxEebT+yQBk1BEL4WxI0bA
LJ/jPrJ9/PXnWxk+IEeMqqJNFSY/ONs8Q8IebYqdA62WWegJ6IcyoFlmI0ZkJKWK1giQ1l8ZKOGC
fZpEA+NYZqeYnlpKzN6MHw25wCEWZt8kltd2kkP2c2V+svgsuni6QIT0ysi59T+F2eocTIn6J6w4
L5jFd41/rRZBWRsLZBMPlSFj+RCqqYKJEWsDjVT1tilIt1Hni2VfEfFrSuwaN51s8y1X2xj649Hn
Lo7X4KLJYYidXi2H+IHqA/gnui7Daikpb93cGJ1gkWFrIrKHBEnm2n7sUk/KDDj+Mgbzki1EngcF
Kv506EqPphrJX4/CA4Lb5/uCQb0fbRvCc5r/KYWhxqOEQ2cnaetpfLDq8hA2G7ZMg78ODTr2d4Rd
qZbqX8HIxy6JnzYma/PCJpVX57+tUjmvbKK+7nfOML5xVxufnwa6OeIMoZG/C31945592RFswS1C
C6Vid16D1sEYbw/N5eXErxS9eD5FrCTJbSdzTeHaGxx7aTiHFHCXna0uf+Yvq6qgvnSo9aS0nDWE
h/Z5gXNenbiskJ8hKJ9cECIvOwlkMfRpVVTv2T+fT4qVbSDSzqy9a0Dfv2IGBUglgLt3XiNWPswX
UbFQevJAmKm6VL6tZJlUuIhY5Q0L0AwssyvYX/LVERnPYJL2VasIpVXPJrG2XLgnP1fh32I4lHYz
LemrMMyFS6OazmVhSUWNbMZP7XZz94PuX5ptwm7L6bP9yGiN7lx+09CWOaWVtixkt5u4dsftPvOG
2rNcdDqdhgtHLejZpdjrhCNCypPA2C8IXOzUySV7/fhr5Q5zAS8n6hU5F7jqvpYrpDJgvniWlc4K
2Q9La1CFyDGUkvPRn2WhkQ96e9j4t6+DahyQd93RGtwRwV8CZ+4HWhvgQmxzyfA0AMWOSlYeyh4e
w4ZSWDl6oM7wCsBVTX5PafXVVCyhH9mqoH8Jbkb83mCjSttY+kBCA7kHLCupU9bf6gBduZNeSSlE
ePI/BfVZboH1BSDVLAWDVa8RZStI7e4l39US7c2yu/Kqt/ETX7CHqCUme/sWT3fvbDRAzt6nw2BF
eqX9MdimmyL6+5eLyRKmBGTphL9cQNdzem8IibHbrKNDIZfHjriIdIzvrfCDwP7BZFoxWvgXSckY
n1oMG4KwpnFi6Nw1L3uxc8RdZs+gSm3Z1NBN+O8qfGpveztJnu2ibfDHfB6t0mslNBKXTHVfgKU1
KxTO3e8yWKogigbr2imJBpYJRZwRRFrjhkgTpovgY5Pgwo1fVUZ8Q5KcaIM5AN0dWCuQaY4zZcx8
nQ03xPxcSirevD+fHi1Qo0zHDpEmPKw2SYJCI1l52cPhLrI+9o896c4cZaTaYF/zL584dt/TUmUQ
jlncFHkoQM8qbxDDf6+ZVDs3uQeYbZp5ipVVfI8d+hR6jE2uYVnlVDdlEHOa47zgQIhb1JiFNUxp
9YVJYEUQ3dMbORtLBWDy3BI9ni32gh98N+llS9cE8YIzLthXRxk3TfB0jMAb1FgRuR5QYoZnUBmI
A8sMi82XEeL9fgoEJA91rDCbrwZIhMeecTLNdJBm13J9FNMA12YsG0S1x9DmHxrXrZI6M49aNgMC
4bG8/zmT5VI9XruFLgWd63RoBWPkWfdm+WndWh3nIg2JJ3ct8iPAS5LF+SG23JUmUqNbpu9vjawQ
Zf7hsE5RrAg6lPWHxmPUik/L86b6h0NCUpwrTam3ttUyyJwKu54BljdJ8pHu9GiSIQ/ihard5wia
EisF/ONF6IoVna+/swuyMP4RoDfsPkexSpluZCPeix4HuNIH+eGt6xcUDypwXdx3OzRvrz99QEjm
pmYyaEx6uISNOzHq6Ze07+Gg5V3IrPaQ+Nba6SGaigG0geQBuIvCcexRaU3r+Ke7rH0KxPO3N9F4
I2c/vHh293Soc/V4yqgvbuhHKzCJgyG7qn/cWUaBTudj11z80D8HeZzYAk/zHNiZRKPl/UmNauQ8
C704Hfztov+9QPlRw4GT0f7UagtD7GB0+OfCgz4CcO82jpwSBPD+sHpTAZOv861xR3fwoJD3hD48
DYOoM1IGRnEOHZ8fYH/G/oUwwTJuFNDvbTbxElhEppffzW5Pzy1zijQ1ILOY0GSjozpP094SZU3x
2wSr4dhTWoEBlfSv+XBX0e12YEBY5cqvqsjpT5JQ4kQfsBw0QHw1pemuMbWB66yrDGe3uhwMbb3F
CEQ9k9+RzTCuPwPa7YdgkIffaEDwASLzZKKq+XUO13SevB5Qgez63IQR5zTco0Dz1mqZK1fcdQld
QVGL9+haw8GtH3g4hE7SztIJZSmtvliNF6Z2zrLpbbFG06XbDIWJ9P/ukM9wqf1wo30+kvDqBQIM
/fIK/aTH/64AgoL3FQICQsPyFYX6YRDx8x71oAdFIsYr/s9Aog/UGtzKMKGd+H/V/DKodm1MQ7XM
MAEsuyMbcjT3REltxGiFlLdj4Wq2Q6rnwRv+iAQJupYHci5jaHoTSplIZIuVm2u3cn+F3HZZ5sHc
H1W55l0NPbjuSy1Qr5QitWD3YTaSJUihjLxopt++FhCaavfY1TUOI53uuz5net2Y0b/U6k0Zmhls
/6ERWLNGhTEpvG4+VW5qAcRQ7DJ9fxEbm9/7cpv/BSvzQOVs79FCsH/bn/oMcUN48XMEfUgM5KZQ
X4CIV98QOqKQPnZoUFjLiHjJUscSqC+iq8W1k81sqTyP0DNmtaoKuRawRxCt6GU8y2E6FfkLZuug
DO33UeLw6xTRSC+DwmV2vf+g1SL83pXeW/oFhpuYw/mxh6+IH3nW9gLeGkg12ulWDtLR+V6BKUj2
EYexagdH99ALoK33mii5jzkWlIbvOmCPQam2StoNKsNPwjxDN2SOKzhG+7AjeJHBePDSiW7Llqr/
qFSJ7X+0Lic3ehN1Sex4IEG9DQbdT+6CEbUk4/IuPMn3JYiyz+0M5qXCe64/kYAI7bf5zeeLnynK
odbBQSuh/x486t8ChzlzteWv7LuggCXD2YyB6Isp/9Fkr068TU1nqPi+FX9NAYXZvj3bfVDznhZm
hTGkc4Xv/7uEh0SYkZcTvn67gja4RN3v01Tz9h1vkDAVKit9qdtrcUdttO7KDxDK2ACHsJZFx/Nc
Go70p4Gsp9oluAqomQqt3vb6W3flzN3YpJfNcROVj+0ECRa2sW1WfersTxs3BBmCewtGvyorzVj/
tZ9nlSVY5Q+tbwoq2RD+KmB4oeAoGwQfv5KTqebJY+ta0ahgt8WNZUh3mrrKGP5f/4/xmnsBC5mq
Eiz2HCxi4FKzuEXca/rpF/Wf7xlg+78TCNySnbBap7FyP/MijQAvPtitLPM+fADEu8z/ruAj/K76
rq8BJAeV62AYrFOQNWSoLP7LIE0uNfCYEeEicvWKNDYUoAqlNWhcOlnve4ni59Sv7F94NHpmr/sd
+Lsw57ghQthybhm6mAyEQU6EJ7A+qiwgyskRqauZA8cs7QQJDS12nmPd51yaXa6/+9TmJmLBH/84
u32CnhWJnQlmFW07DpVflmX8X8qiHfBqdaIZ/D+OJ0ee39GUizIKOT6LOwEWK1A5VWqgxdMQTc1r
TxlQpEG09afcytJgHbjXNFRKDC2v+Q7t3IKA+JwLbM+bWSMddZIZCNFJlzaRlbLaLOavSBfCmAr8
GSCf0bGPnltMRgd0AVuW23P+8E8phfn9duy2Q9YvpLTlpEwX+q1iIdbNmgZ0YBQfpSGBGRXKvT8Q
0L0b97OX0BcuEUxhekK1PdSe8L3wFgN1/5kX35t8vV/+2xJdX2mwtE5fcFNChYdhfRnYjUUuQZ6Z
WAQr/HIYegfjv1KH1JVMiTeTpk6K+DWg9l/9TEXPX1wYFzEa7LqnzJVaGH3Fw0e3wh0cEp3Oge30
qsQ8haoimXbIfqR8JpOItdQQY7HqShFfRos3ybX05wP3R4RXwXpQ41PZ90qFPpfzElMj6gb8KI5s
sX5FD+SyHglzlxfbh/TJ/38vY/wV+yBfY6NhsoczxtXhBym0BREdze50OHPgMGxAz6fULEpItL+d
uvRHuXDLawx+NFXzjw+i21/XeZ0V1PlO84Sn8oS0vwrS4fPyZHvxCN4HAOe5Osqd66P/3b21jFv3
96+DdLmagm18YI0EK1oaMWARrajBvjXPkF+T6SDEAYdj+OhM9xgY6WJ0uxNRq/AKIj0cPdeOZvaw
kL5FlJVbdt5V3g7GXsiOrIA2pwAYocTT5Yp8VDSdSEQD1uals6qNss6nz9/aMw9LuVhLr8V5qaXN
hPASJOVY9qQlHVWrhCRLWlo4rP73ojBHt8HoDkxY6yLFeN/l/ZqvCtCDtXNEHFkfAcCiFCJMsgjf
3r2M/QG0drw4RagC4hRghrOHiUM5qzftmYhRQjZnZVcMQOrXQkZwFaiMgLsAbq3lXArkLxdUEUiT
fCTs7Ng+9R+/lmb0gxJ8EsD2gysDorXKHjDkICnHSih+zwsFUg7zJQBNMQIEvPkDQQMbX/x/vdzI
xmfMuysgNqmn49egBsglTJ1Lz5GgRCZuTS297VhFayWRm80QgAem+w+2P263HUb4PnTM6rPGyXFB
DXwqhljuBu/159Zr6xJVeEOYKI6H/lx7kboyB2LMEvgtV2Y4cvA8z/ZEQsEi3B2v63BysD65zdcT
egp6TuyCkBW89yT+I9Q0aOC6qKXQH1v3V5q7LAl4rgmFHF8YRDOkSbVQIZxJAwSZ/gr14WJZggjw
udoAZ/iMb8yu0GUyCEwW/4vpp0Gg9N0cXQmtKPByRwhSn4ZRGvmrMeaaW99ZfDInJX6IvOsYTwZ5
bp12+Xe5rQvyp568QgzJuliWE7MaPSkw88NwHPs9mt43R4GnM8Lu4+80DVy3y08wx4kV2rf9GxW1
M5jOtEXBT4MY6i1fU/JIhM9VC0YdQQ5+q28OPdBzD4Qra6egHu8DWJl23930wrwkuvsXtjn+0NLE
uDa/7pSpG7EgOA0ifmOwJcQMKFDZ5B3+dzNarwxXQ7En+SRFDbYlGww1vYK8nqsYeEc8UJ0MxYMa
b2UUrYJqdSyCS7scM2WYd0xp8o+JSrZM/gCGuI2bERunNU04SFgbHp/ssk4Z6LKONBzNOYqe27A6
4R72vMkXWAtMCOArq8sREVsf5hVaDxeaNKGMQoMBy2r9mm8386x6HxuXlj0cDDXOIOiQ5rrK7MBh
2yzo0n8luuAICQsi2faqDZkx54FXPYVUc19nyzy6/+NGjy+jtSF0UC6e1PxiHUyib6wTWF0urpCj
yudhf+8i8mcDz2FQ0RItzmnvSJ7E7sb/Vp7v5eNpElqtlhnUDkW1N8t5MBIEXAA1M6xtof94/9D9
6X6qt9QXbSc5KpJHSgrpGEJXQj5YxnVrRBCONH/Hpe5uWSqqetc/u2Yg6hHWsIGSWTR6Xk5LoXQv
tyxUcL31p/v/i+WQuPSfqLl2f8VtkWoijvXRaQ9BJDqJlqDKXJ1UHvDDFXov4JKo7kDP/3G2YMZr
vZieuaS9xxfZ/CL/1FhtC8TwggQ3tueMRLAaGuU3ToJ3iy3VDv6FYi9wPzUj1xsUhrqBcyJWABjd
qKpgiYwWhFT0kkTRFdCJzUwSIe9PEjYCdeyMHOplqk2nuBNqnEPWZmXrlkrFnjjXHciR6EThmN4g
QNSpoCk9PtCKJbPPW6O/LDM6nvM5ObVQazv7v5tDbc6xJwCD0kYtaVOralZrpMUeQqevRDr0/BSF
keJVYmuhIPF1vxyH3agsR+IuItZFmPUUqMBcg45lUHG0vpv0RytqboluwACWta2K4wzsLpr3Kuf8
Glzlboo2ockk5YkLR5wpYqw57v3YPkdjUo6jyb5xPw7PPtsNIPskWJ29hBrZZYiURgTRpIv1i9Qv
8CrgAf46UzfyR+XdwxoOSvrCmpo5lOCwMmZ64bDahOElscciGB+juuyrmRAym+sjes2gcrM2Voaz
UgCDNe1z+EtYHKlZV7IFm3CFsboM8h0E96CF8reOU8aEiQhKNYBYntiob5sKZ3TnjjcO+37DhZOT
y9qSGCtM8HMj/AhBnZLVgXRNRTbYVSuiOcUX6032igxup4oJDKD6Gh6rbQf5jEcHrWOBd4AHjmSm
gdFbYymAeGnimvvc1il9H5u5M9+teCru8Uzl0jAZO9j5fzrxXBHf34407yTlyOJQVLrQcLA4MEfR
5O7FERenJ8UXaPpfG2HQqBmMHMm3qvDnzN1Hnn0vlazWFFRW7SLv6USR4QPT5RGDqTBJgXrN0Mqw
gpYCyljkVyeNUjeyQZMut2K3bIhcoX9S2qUPkPY5T/IJMxHpdZmBwF52QA25ROR0906QxUdP3ktH
oDqMR0emDxYa67o3gbuxcz9GsydUAS7dZQUD/KdOK3QmMi4JFhSi8/Zi2ZJCAk7fYXt8oNWnWGyz
etrw0ieS8Hwc75HiHrnP810icL5d2i0A5p5rGL3H4tWU2FqC5R8oYc1DG2Lg2iOyN+MYgThXYUVx
CY3t42SwP6GB2Zs4DB27NFOdy/bUHB5/7UmnP9hOMi/S8YMOvIyq0vbj0BV1QJGwyPnq/ciqtPCM
keivVMlkupx807HYgCgCl+RfubZWQQKEnOb4ZtTk+FwEPOXMcwLc/5z34GqBgBMd7MYQO2VXLzgG
R3STDjzvwDyzWu1AnpsJsDPFyczZp8eLokXkRRuA1bbngbF8i/vjjOAVJwY2KmxBElC9Ei9ssC7S
BLZ8ahbLinjtKw0V1wfol0uDe0ZvZ7XxCf+B3AU0/DyFhJLwMC60EmLo9Tz+NRJUCyA3KEvicFq7
tfkaJZp04tRpWZyCU5ne4MFU67OhDKmCo8vBgfsNJoDZNcuZOci9Xs3CpOisyncYMvqVrszTJlMu
KVegCSnvXF5/BD8HclksYURItZO6loBBhyUMDczrNQ45wzKjfnRJ4lzf0rQQAyfg3ro6frsMEAYF
mDBzX3sJDUzyVDTGaInr/mjOfPkrscfAUdrIoBOpImgVJ6wHJ+Bnk63UUOy1KsbFfV7yy9xeL3Xx
hd34nz2XxLget2ogKVjIxeNCY0Hp48ugKuCA8Jx2in0NUHlj5n9u368+kARo/ZkV24OZUEfU54wR
Qki6OtH+M5nZwZdb2BlCm++XHQa+fNxGm+c2F4XiCyypI9FTLeEISL7UJ58bYBBKXnjtgG34SgGD
eUCfVQ+Pkbl69vmTZdCaZ6TvFub3bhUy3dNuD0utnopbPjrTuyDlqMykbVqksztzyREZFFN7a5wh
qgOV8rS7tKjiYi+L4M85xr0YAIesn85I4zoUNaeCOwg2+2lgiG+p54GZzYvm+6uVpARS+9J2Tjaw
ow/d3z5CSXrH/ezCwmpxs9I+ajhCyRnyA+iX5HxFiqA0vrmiCZPvai6qsi06bwS6DMsBGTFNHoeA
eTcUnXAMNNBniD6rELYpKsoKyvitj0qvqW9svc/Lx79GMuVoHVrO/AF85UkZz7A0GR3LGbSxBF2O
5dchaUoYNj1Adt5ui9yWuea5EGIeenbpONVLA+VPgksgZvrqWU3C0Mj7yEfH13zmQG/g0MFzjO9q
unW6+GoDNQbHHTFk9bFP1hM5yxUEb1erQU40EL8fwsnh5wKQ/klEELKPPmAgfPmG3Yu8plbzeD/N
38ETOnC8ece/VFmzUdpe4M3tInmoTbwByJ48VKbj2j5GZ3L3BumBj5kMIE9wsTvGTELkdaHrjZqH
i9OW+3H/lG+rjQYLdjwaQDP9aXEJuie2Jk3HUIV7Bfrbk2bWyXw4DOVPL17PlZVE6LYkk6GaIy55
SsC8aJ9K15p1Kct1umOiceCp+hZrzAmjCVqUiwiLr9NFGE7aw3VKHXi/SW6dl7gFDIh4Nuk1j5UD
sHCNfQPTmWfGPp9yBSlAXzfzJ0/xrL5oKPPLJ+cK9vUxdqfB/pjuef4YWDIvSrgfYH7KAVPxC0aK
VKjCdgf56A5qUBsKvlM8utr8CQklpsA0k6q+Hf+EE8ffc11uUNmRXVEshNc41nMwIFr3VEm2br3M
Pd8n2lq+dosg2YGizBGhue0oaAFk01T2bISJquPZTkB6vuVYS+KsP+4nu7Ii5LiMBQNQ8+MxcfD0
SWG29sOz82QHARBKABCrdOdB2mqaqMTVQocjW8anH0Ukdn/5pwBhG2qfXBL1UdTo3im0f0LZ5cbN
VafIOJfccpCif/Yoj5Ym9kQX9UO5uZ8K30BuAOCdGxJW1YsVToBvUt529p8voKeqkP94LBWjHKhC
O2sVwirDeV+eaN/UO8gFh+xfyr/XJH+1GI5gZ6rgjSee+m8tJvx4edJXFlsbNG5/UolBLWC09SQ/
iIlnlyh0b/DvKK0him3wbUJ6s9wgkErW1ZJ/gY8fNXhZfEVx8eH9tgiX1p2usb19V/z69MFY1d2n
ZNHTXusBxG+Bj92S0C0L1ryj0o8VVggPq0NwDSoSaKbtxtki3Z3g244aZaGfMLpsknmmjSG5buCL
sSEPDOZLJ9CfrTVU1WZiFEJ8DE0xR849pzEjVebCtZ2ZUTFJNJQ/Lzfp3QRGC1+q0h/ki51CeSHV
gx56yRCTSN+jF6ozvCXOwedjyNRH6esh1RBctqDpApa+d5nOHVE/mhw6B3ebw37XTXX+IyxKeKJ2
rTpBeMgUcTcBGVYrVPW9A+3uRMIVuUI55iqBXhNGVMNBHTs5g0FVZhDwrG2QR4nGVjTDNttHGMzS
9QAXKX3ej9x8si32WJtNtzeQBSCX2wUXppmP8RcvqV/SV2qsx2nRqMZwofAgd0nZ9yhLivmZ3Rqn
2wSaAJd0wjQBW8uDFOJxQFZLkOzVA5GplcGc0/ja1WszC6x2EWUq8lPq7z1oN6z1PZXJAht4+UY6
zdNqpWKoQZxlXkIRSk1S8tlGBrWSxYdDt6wcunnstATLGkT5858QUfp+Y5pgR4pAoWEJ06aUKcwg
qBIMS/LFEcUaNIrrP60+90YrC+q33zd3FgqIzPt6fUPSWYP//ddVyeZ+P2EF/4XodrWM1pSjVXV2
RwUbMpSWuE3/RCG/uQv5A9tal+9+i637Puzgjxgw3pF4WrIIOIMKgLlBtdWpzp+DL9OJtqXRhYYh
VR28Mtu7HpNlAk8J5k2xTtrXHweiQyAOCozFDWwPdx4P9BHy6+RXPKIC26EOAouOdLWC8dWWMOwZ
Z6UKTXh2vZrdkZxlFx9dviQ+pmeZuSKlTewMVyz8t0rIK3wWmeh4TnlHCHfC3oA/G1HAgA8vfiCC
ZN04VKI3WiDOl2N19+ElvzAn0F9UdGUBunFvGnjtmywhL0ptv46uJJxeZ+VoQtbZJrABP/jVX9lw
2zlU9s7WS0ekOk+vZnyk9r0NVYUEdShbreXuc9ulqpBlJJAffjCwQAR44vBY3ju63Ydcl8xOEtWZ
e0tzdIaiEWznKFzIONP46LERqoziIEVPVMAqYm/5q20WrtUhJR1BzFHYalIefl7FJTgrfevr3IH5
fSfYJBYKaqDzFVyy+DXBvyTC0uTibR61ipw/OCsiPDwthT+SVAbKrpqL3RKa9USwmpp+rB2B4siA
kVg+ZelhuUXMvg7YBoWjDaYJoDCK4LTVwXRal84gxl0k8wuS+aPSckQLRBOLzm9RnBou9GpjcgWs
sfT0jKuj1D7vtdwwWCn9dM2kji+5Xf/km1OyPS+iU7SFI40P6BKtIVFM/SgIZ3Ivmb/fV8wGlvfy
stN9BmOgsT7H4GCqKCUPM3hxCgk3CLdUtDK9BouuS/9w1LMqwyON2qwMG+pxiDdVdlwK+09irF8f
QYFS6aoAXbPtNbGOm85kt9h/xUOv209/0IuQimrp8RQ/YdFMWGTZqhXSIsdk9bsvBL4dslucVSTU
pOeUprWBxtSKdSVDFYyWJqDgqFRdnwNtgSjHRGUYH7bu7JZV/B6fgRzisk8tQdFugaD4//XX+VkL
UIOkyrwdFY+697EIc3kiXf/yERpmZvm7pvH3zBHP2Jndbo5n6m6P/sKCecIKLwd7RFLHAPHwyNp3
0vTRLzitwbXBQXwTHOjEEKlKKrF5K4N5A0TlJMWlWzraTf10bD8gbfSMACWPm5LKfSq0YuRCwxBC
iBvlXmY3hhjf/7Asgf3tJgQScb43tJWZ4A+JgPef2fnN/XjPN/kBZvbXSZJgAXVE/5g+gXQjmgxc
zpJrliTnk383g40TIDwe26YY6bUEAKRSLuzQwBDPHQ54ikl54xDe7kEs+QAFLVd+r2L9+MIx65PO
lhB4jFwpyJSlmnpdRTW2U8evil6zLyObCQF6s+7Dcqq4MLmN1FSlttJos5RJlJM815Np8SrZH4Me
JGeyD7BgDHXFLQjmMGg5UCUOgVSO64LaheRpKnkFVBmIRo4UThnmt5D2JRSf4quW8SX63pypd9V2
vkMXr+6/U2ogZV7oeOszh737XSk15exYqOnXdaOfj2fGMc5/JfPqx3ZTsfi3sVv3+pYWqe2XCmHt
td5/Dj/FPcC3BpRlixYggivCU1TIZE0mRr21nDTa0+GjiLx7U8AbixyNTjrRLbW4QsAqNSLiELD/
xKVclH8FbjHooPUAf8U/4FDoLNmWfyDJGErIbI3zVqoKrbRWwpF7TDD0FGJZxDL8sDihfP8LB9Ds
l6be/u6CMWNAya3BH0qUTllS6metzdTNWIu2M5GEEhqmLTpPlWrWX87OYg1bfycmM22tN/7gQtvA
mBQXepf0JRkoaKBA8dn9HVsJBztDhNpyn6RhvPZMuZESaROd6q+cEfLb4oYVUw0tQM2KSFANyqPW
V0iIInh6ryGGmByHOng/k1xyvAkfeMNG47kJIVbs0ws868OkCzRikzQV968DFu0RLbWdcb8k4ojf
Cpx9/iL1m+7RM9IHx9XzyTDbl57Au4whFfKF8f/fTB1jVUQY8woAGgkNNyQThGLp8qTRtP2TH8wF
0PAuXxWgUgH4ylrKxreaREncVODADMZTCkLEx/mnuW1hh0UBoYuOLRbqe/rOx0pWBtN+NL80OwHO
gqKmMp0+X5zxu/y0PuAdClykUMQqXT9Or17qaC/4T4oXGQoqGCBo+Po1qBY6tOJzYZpFZL93k8ap
HZWo9Dd4hb5p/+aQ6PJDnG9diXyo1Pw23i1XsiRTsmzEICFKKKQiwAhdtx0qHENolDrto/O+aPbO
mJAtOa1KSxX6R0oN6bhYD3V88gUidkeP3Q1B06eQUC888uLTVir2es7ijUf1WC7gJhHot9WoyY5c
7atHLEtGvYaVfjHmVrBbdoP9EKeO2Fby9itx9yy6OSffEDTD8ClX7QkDjyXbm/Qvr32j5mZJBca9
SH/vWnUTXhbktREwTMmmf0ZtKbBDayI5VIq0VC8INFG2+pArlgpPGdCOMqJH4AzzAJykeM/WFuVJ
aP64c1Frit9dqsLXdDQi3VW9s8KtRRAIZ0Hl02cgpR+uwuKmElZFkDJipnGivIXfpFhaIt03nbDh
NJIn2wbVjAn499gYBDmHhUcPrZ9DMgkHUK0Pi+ugFM6I/p40PZkNu7jS6G2rkpPio2smKmHYxB5L
x1FGo/5oM05aXlz/Hb0gwRXk91nrGRaIM9W/SIZzLjCimc+PyKdEJxJRSuL6G97mJtkeF4vxuRvg
AHEXhmMu0s3Vm3pNs/R+zyp3z3cyGr02TeBbCaUj3j2nGW+IX8oouua4LAEfBYyAlnlqE3uklInj
94PsVP3EhLIH5KbCx71iKLZIqegOxncoCCUsFxi/iCtBHJx/9fx5Sh5AY9C4NaCJFsEJWjkdmISs
ls+1V/D2MSfmpbp9HHbk+VHY6sF9SaT3lOZRFdAKMV9ajt2QmWNj5PqzemW8Bf+2e7QXPlvE/u7h
8FC2PA71pdaZgSwfwWdYToVu0hDVWFX6gs+RpbcFVUI3K09hxGiL3M1vz1OoQ1WXi2G0KXOpMQYm
r7Srh9wLll1fj5pe+5jXgy+PjyZdiB4IJB/tcqm1vjYEn14ffcXMkskFz/0WcnwBVCXX1j8u+1yI
8rd56TsOVc2zAv5ES579F0KrAtj/boYsvNWomrgQuwTSBT4cERLdgH3b/g3EOHGkTfrYlNhwdggj
p4kniuk+VHEoiPgWiOl2fS8PSEE1KjSgAo2nDrHgDxKwAnQDfBRyHo1uobuk5ljAvtsAcpKgZxaX
hCJ4qDIYysnJ6dA+2VOnivRXjyUyOfGIW/ll/To6mGLJcrFawywxkak4qPNODbJdBYffn305qvi+
d1GB41KRcA+x2jje/Hkk8Wb/vasL6tUUMxqO8Btn6IZziUBBTI/ALyKe+U65++VmDbNfYNCA3AUE
OQzjAOGee8u2Pdv14l1rizBtCn1U1FiB/7NzsNAfU83UMhVVZxLJEfiHqgZ2wfCHlP4GNGE9bQsJ
LDOYZUhhg22aIJKjUtRCdNPeoVHm2r9seZG7CnyQ9XBXolD378cBYn2WMl4UTuhWyF7vyMcvzuq8
pa/iDetZ8DqVit9RNzcDk4NESTzqqCQarsEaPznRMFD5HcS05o1zb61WSxbSvWEgP018Nmis8tuY
bZmA0O3/HJnzUJnw9vvXI6t0aEoi8NnD+IwCJ5YynFjQPv3AGrooIE0MGLybNWm4C/VcS4tlxONg
UP4rWVQaChoUUZ7k3/9aFYq+7XpcdaZGgqGwQFT+AqE9j0Sqa3AGVcY5r1D1b8BnboIVZeLSUsvP
4QfvADypCFg1zSoam1iUK3ZN1RMZRci7rwZCvpdU4OGRXbjqalGDz11hDgMClHczweC2g+y51F66
fdvAU+w/T/nXjql6n/U1oBA0YikBvoBqjeQYbZL+f3ox7FYT+4t4fJ7r2Vr6fw4f3vdRInKbWu7J
VjwKzj0DmJcly+x9F1hn+i/9i324jWJvfsxYib8gfzwUUChTHxH0DgBa3FvMmvNiM/rUSsFKHPy/
jo31NXXETspx3tSTA5aRhTnruoXB0ukRD7fKoOAyt0EvemVkmwsWpzCW1HfKyaa1VDvLobBjYMcW
zNlbd90ggfx1pdhcbBlQys5IAx2f0vMDD6BlcqRDkbFoOExUKCCbyKh5pSE5JK/c9b0zPe7Evvu2
CCmPOH9YLC7uP7DoY/tekuDnbCTD8wfw3YiciAuZyEY08AT82Lzur1zcbrDdTSvFaJF34fHW6TYn
++vrPcMV+es/rkX0WgFBhhnvV4yCMYchsTh2HcJi41kOrcjApRbDEyxQBCvXX9QxBNk2IyiiY7bw
KmF7cnHpNoIdd5WVqHSCkptGu576vrfmIzv6gS/a5+MGmy0tQQCs/XFnia73FC0Y6mFhzVVVIqVx
g3aUycZ+Zc47c9/uyR5mldOC3D/ODHR1I/k+0dRXnpVYlRmUBzcNqgR+ibUotBYvdIKCTjfM5YMd
K3WcybZWck0AWWk+1VcVCgTfIZobawiTW8F9uZV4FthdvSMgXGys1LatBfzCB0yh5016DIG4hbRv
4xpvGhNIjxoAEb62nomaBNGCFSLbWdWrVZZ12O17ST0/0x6Edevh0jVp75chIp7RUmvoQV3WrQpP
IOqotFDYRhvEZ1AIYZ0JqUTLejg+JZXGY80khZBkGRI5ouaEr7IwWf8CZXuG/KBXqC9PewVj5cdH
q9V1aLszIdGli+jH1G1A7xDy4n3GBM18mczjf9biiA6/Obo3KFe2J5z0/qSjdySjcwHOVIHpFtd3
Q98tv3Ra/oD9rh9Fdb03/K+9ALnlXR0mrVo4A5hDrabfxGfM8wp9pxwmlJ9hSrUaBcfFQtm01DyJ
NZ4IJZeH6v5P81P+Caqh+kRHyNzJU62X6N2yqblqW5dSwHBogSMbPj+oaa8AWiglJK2+yDEjmWIG
rHG/M0bCOTmOT87UoOnkDhOcqjHl+AeXzHJk+tvzWkFPlXICedfWkJ4ShJXv1q7o9Z+NvZvKZLz0
R1yPSt48UVusbaGp+FeowUJeWZLCIkzMbtwC4tNMzAwIRJIgdc7MFRL0aBNeKn8LPw2GYx8jf2DG
XN27Mdf3xWeM696lNlAm8IX72aRQWlOpD/KX6cG2yEqQnr0H0aA2elTkY9rPVgw4QvB1sjYX3TIG
3eBkO+7pLExrI5/F6obR5RYoEheUuJgDoZQqJBnVlEjdTOe4f69vMwhWDoaUSsyKFWbb7w8oHobI
Tcyj0rSmmbSxPrKVWzcxULbR2hwQnHRxYY5WnC/bvi2E1GV/BFPJtK4JnmuYaEZzxEqJ/3z/HPbk
LQzy08OgQSSzC4PmGS9aJH1hbKAx8Ynoi/G4837Rf8qnXxdSxi9qICtgsaXB/k0ncmiLWj6EdUJQ
nA7+E06ClNoUmFG2ZW2OurDdRKIuZ0AKN9suAZoeA0FIFXGyrAE3E11a/u45VixJqArZdVVX+Opt
anxF2HdZWSN/dtbLfcglqQEigZDKCAS7vtfLmGcTIYUigqWNawzLq0FtRJHY7hswEDgjOBkoYdbk
Y3LM5elm4uQf0k0cmD4O+z7dOb6Iil/CXCd274Fzp35vo3QJUxPBZKPkiOPFpeQfyvgZErhcO1U4
KnhwttiAOb2C5hUJzM8Enhigo/bB/hb5unXuc1sLGMz5ryNDvc25AiDnsGKoao6TScRPfcWzplsV
hp8Ff5jmhGm7pfNw05wJMZbB91DmSFl68IEpl22NS1x7Lu0gPQJMN53cPN7v0Vb33AqhzlaV68qU
ZS1SiKYc44p03iufT7Fdr/tvWP7zIZnEiy/jKeCaXiFzCC4LzeKgAuoH+houDxA8dD5RSaCe2vSY
DPep5yFUR/lhO6Q+wZkHlTRSdHhEpHMyHgeQQyRIztthzOcgAwgUVNl1/gNG6D6xnDjCbl8KsZIs
TdcCECyBOI99udCYcMp6dteXlhJ1QdX3xlQZTDWu/ZEurpSCqXKZ4ELVilHKUCq0dnJ9/ZlT7S8p
a7XNHXTjjzFBsBDVU6R+yaHryLuR6xYcKgouYFttoPjq5Eo8wGSrj4CGXF/yBxAkrNSGnZm86DkB
neHiMQ6SIJupeqt29g7WPq9vax0GRgFqfdCFe3X4R6Fyb3USF8qBx0cyGWnqTjAZXwWJpit/Szmu
HcS6jiM/reVpnpHVGO7PTqx/KOHZ7pwcs91JMgso45fEK8szltfgC+L+qyZmTPp73Scc3h25PKEr
M9n/orMruOxfyzz+u+MASUnw7KKdTm7w3mGVxDnTpbK7w630rzD9A2pb6mWS+wC7BEd5ZL3gv948
/NzPpjmDLTTUFcBkewXeH/67hgVjpJES5oami7mIjG5uzogb1+tSzD5+jz5g+erbakzPAWXd5oQh
gfIRRan55dT1WTWhX378hxwlbEYxgEhv4DgWry2TmKpkp4kqbvAeMqwWg0vHdrPY5Bc2X344WFmt
fqOdEh5Ra/QYA4Fy96ErKOFCUzdMvpbhF/psmpYUtGCh+Kx5baP6d422KijvdWfFrXr256YpAIe2
rqCxJHNLr6AZMAEQ5shWrmEA74gepoJCak6xtGzkv7jItJZEWrUeD5cdhHb4NiKbOg0fPhx6IzaP
OtkEHn68Q3drjtPS/O8I1oqtF/AoyaSyIJt1d9Y6U5L+eo6agbPI2McFh/QKcftow8SLAgAB5QIS
Zi19NTbI5QmQFMWSmtRUfNBiU+Oh9xCIDJMBA4Jq4Wp+XFgRPoHPypkjGqIpOll7QOPxE7QNd1tI
+eGwBdAJgpHt5tMRXGAQ2wVcHyZ68h+CFoU25YzZY7J4K2x8xJDFzSDbncw1m2O3C2omWlUWuwXV
p9Coao6sZcF+33GQCLRdNtvSrkxucEcBklgB135t5OZB+xzqBsJV0N+QWTWW5gk4D/nKv50AlPHX
GxitSZHFyiFVIWWdMFBIPDc87GrOriVW8zt1C43/jdlBfYo0uwvPjX6ae02qvy82fqb+ik2HkcKP
R7Zqiws9L1YQGhXrE3/qccLvh0sj64TvXZTTrtk+BbaHSVlk2200Jl3uYC7G5HtVwHLApc/XIaR2
pEi27oyklwEqYTIKSQ5FMdVKtrXIQknv/gCj8Dt/KQcLrSc2SL5pKokRGD5gZLkTexaccgExBuW5
YX2BLmOrpuc5gaRxZ1zQRL/pnzcRGwkp14GZ4zKnosrbHO2lzN3Pq7UFsJmy3B1+TFBAYRo5l2SG
4VTiMbBeDWbkKYyDfGI0buy4iEbHshPP8M8Uhw73FLzCxuAKHsUjfK0AdcGjk/GYniBECK/huFlp
H6WWXlrv0TmqYWpcNxT4FMfYI0E5KMshvAmgL8DyN7kRQTdOVH4buLJpPnre9M1N5a79HTqmKjE3
7bHx9iLH1VzwZrpy6/U0H9Hhcp+kJY+OI3+sX3YdK3PgZ8QPmzELf0zvAMVUUkq7oFKZFrFWJDq9
0SZv9w6H9WGYj8a6A7Het2rgJVf+jM/5/QRc/V/V5ITDn+9uB3c3CJboWDMtQ3YtoU27C7D+KhWf
frPWErL9JktsA8oiYhvtJUPpzwy1ehVOXT3Gzg0Z1Oehq3P0XeDz+h4ea5Rnp6xNAjOQKOcnaaHy
kzxxc84sMK+L83uVdPweV+Ky5oi7o+fKCjNnjTCfgVaA9Pd1NwpElA/ZZ2k1LpHL9gLXGRN9SdA1
MBMqfk2ONd+wOmSLFPB4ZCNECjYbS9T02aLURDW8FYBwSIzU6oMi3udc0L2uPkUn8dnAqv32R1cL
bD27JzcrmDbSrauysvLMkOb4GTsFlc9PU8mA89nd4Ay9r1P4U+1rSNwtF+3RbpNLreZLjTrxvpUr
odU5AALDiQvaEbqZxRc0IXVbDYfefJDBvQxBCjV6D4DPswz6Och7dGeEcV3ePCTq3i9bGYLDx/Yg
0BOPOA4LNllnPtMOZgKStukA6IPWPivL4VF+1xpXWOCbGt7UAHtOLH0piLr9VIuOC4b7V2YH8J44
A9Vqc1rJYr75E6hGe46TGhUPb6f1P1L8lopWKWJiBLzIe6M8LqcEih2mMb1gTxa/1AIvd31lO4tt
84g5KQ7t849L0peh4T1vpnlzz0b5hGcFR2ms3wP3JSsUo0oqZLHGBHNlUE0ckRQKLIVk1iN3CaY5
ecr4PPM6mQXPFTpuzVCuhyCi/LxEJnXl1g6CUTtyftFt7A1exrcgzq5Jo/B+erFCWl7gp8cNetzR
2xjorbQ/+/9FKMJyFbzkjYtm3xE1/OwWpZQefkC3/e+LxBJ7tRqrztSXUezuvXtQND8U6tpGaO6Z
jzSX/g/VkcG+95zYIvj9WPR2YnvujMY84yGNIDj9XPmQlsklc4WQwsaIAYK1bCv+XCP24nzxbYkW
gqK6JNnQmm8ZrroOmlK+qTfhI1qK14VMwlCmPqL84FUQpHLQ2u2tDRme3JuSsVPxx4gRfytrgeAV
lbSU5fBzz6Wumhhl6UtGwwDNhcRtXk5PyG0C1iePD5U/ngwit6MC58xP52FtMqxNrZs6+67+lDEI
T6ZyyhJv2vcoZ7cA2pdm8dZvV2VeKnQhmILDs59DDBxU8i9zeDatR+UtLVa3r9qyvtNzkSbp0JUs
OVc9bKDS9BsPNay/23YinZy3BH10hnRvzkKxdXogcIN6rJdVq3Z1T4vcc4SrJUgSMFg482Va95b8
x1PZL6CkbwywA/bng2S7P5MYeDemJ5A5bQQzkhDPAMHj1TUudSo00XZkuTtabrN4eA9vhIoXJAlF
2Oz9w/pIAberXwKCit8mzcKk9IxOl2lfSaX9KpF94M/0uQzCZxuI8O/atKjR6cLJj310JKuV+Jbe
fyFTskc7PyDQ2gM6PoQkSEDovy4S1k2hDKY7haXC7Mv9UhRlSIgq9IoMqOjb+xIv2lYB+AlrFaqK
ntHNDttPYMLW7iVt4B5lcLVjki5JJ+Hq6mD/NFucasNsikvS/OMeswNz9v/FcQJ4NlBTt6J+HJ1h
eICTkWmw1B39uZxV45aczYUVh0BmkYyjJpyV2WIwpVAij0A9IbQdCsSUS52mZ4GDJ2iMmsBBpGRx
lwEm8BUov0tElyC9E6DnNvUB+EKPvdzA5TtY/5zCbcdNXniLyij/1AE8aqiuDRjHO1X5rMRcb5lc
um31PgcdTOJO0D0xHXSK26I1WOErydCJQiX1DQV9bPNc/DVnXqdIXCVQhk71ZfNxB5ZHt1c6of1q
XBRkyWKCGNFBkp2J0gAtiB4or/m2kxDV1/c8LHGeYgd71EFjwfR/5w2rq1ghOBZ74m1Kwi04vJy6
rgQnlVPe+ecFJJA746SMYRYxXyRJrCUHRzWlpNp8Kygqo/1tPHADqCsmZveMTcmeYisYs3Yjbve1
uoD7XwlJH5/jNpXiv5Vr1yGCcaEaRPxZmX/17xock0quhZrPob0sPEATznGF6UBJnZWcgQDC1II8
/ILg6Wp6sizUkCiBTJQIvSEXcTfzQokoqTj0H6zVQHHOXvuC2FjePobiFx6jiCOFaanuyVYGPhmN
5rc3TiD2tPIq8C2vGj9jEwf6w3FubFO+AJV5qzi2U3oC+hze5DOy6FSYLj1aL0Bb6bvzY0omIBik
cz64gSCWJ5wcxg4gy6pYaXjf9BmqJb70GV97Hf6y48KUN7Rz/7ex/frVZeXzpmja9qk6DfGWkHKe
9C4Bal75gdo2ftB3qIB4qv8BZCHSkk2ZCw2spJXLtuCR4JpeC5SoLVCFMRee+QoUIQiOv7wUIiYR
SpyKJ95ExvzLe+5Y3ysPGONLw4iOYmksYrD7FOhPg6OSu8s0CYO0HbBlyQbQgLUmUl3s+L/ypTmZ
+SZLH6sYelaK4BnoPymNLt61F/JsjmDDOrKqWYx/YgRGzzA81GCBgzGbMowBEp09r7i0J9Mk4M0n
FaoqmSXF8WQv/JsHsSXxXr1STL8gJmZaVs5Nt/2irA0oivl7xq7Q5d+mS1dgZaVry0pfT0i8YuE/
b3RDRTKv6n+c3PDOIXUVIpPhiyh8Omd+Jhnd79vKzOhepBElU0E+XkLwOwzhhIYGr5ZRqqyZXGoj
+1pstTOCFOVL2pYXWqOoZbtfhw2k3ol/G8O1YX3mAiY/o46j7rCXivW6oQ3yjTrRKh+GJnL132b8
CFWV1QrK67i52Dw8meDFZCYmgffEucoyec6sKARPagP9d2znhN1dKwN97eD6lN78a0OpN3RZ6z+a
Sb77+KRDAIV2IDa81wQHK54h5sQhgk9EhYCrY99ZP022khUsjN3HRwF84U2rs1imrqgWp13FKJaw
lmxxOwtpsCMm5Y9Z5Jz/jAkTQU6TIn/VKo+0pV5i6WNX+bqjsLdp2tmZyM2P8H/V3BlKDWEXX5hy
BAFvJFJUrVuzQOF23s2sq/r6fNRygwDuKa+QYvLataozNkBN290J0LQ7XpRNvUr6SMlNxrL36piQ
Ms/oz7kyPFfN9z+HgigxekTlFsjxicJbU8nTtBudqvnTT58++Rvy9dZSUno/X6b7GNok0itt9iB9
KyLBz0mLYtdBDYL6foHy1gpJPE9s0KtDpFr76gfIrbSB6VQQENlZpw4too6w4xqCPh4KaIMlZnfs
iaHMEK6RvjaUQv4RRBPK8R0z9wqdkXogphQCaXu9z/h/WZK4bYhdUymDPW1a00HxnbdTGpWaVx6m
Mbx0Te0WQ/xNidy6ZhlEngPgn9f/p+xVYOsU13IvxT8Md9hYHthGn6BBlCCwjzJi8iF73iERW4Tn
Wo4vLuAdwLqayLaEbeYpjn1YsSfE7p9mMteWPBQ9VGfY9qJXIQumxS/5gQGlh1hfmOWxl8gQYtWw
ofW2EjLIKkhZmc0qd9QeBAOtQUPtkE88N0LA4HrvL1fiR5B+EgtVDQniUw05NNK1Ubv7rVqt7Cei
J1pSTXQZaCHojINmraLgDKxnUcHa6vMa0WKTW5ZoEHp706t3869D3PgIYlb41TTAHZh5tpomjXdk
EPuCSvbcVp4NOtMSLiBAjwLC8wCHuaEUcUF9bWpWeGoTW96EnaErNw7Q8HD/k/bHbyokq+bivpmD
FweX0n/h3TmtKUhzanIIxdE46v86uHflPZjyhFjbd6EuyusVj3d3pX1KN7TovKVdH1rwYi2x1gHP
/7rdZKWZMZGX97XnXdc8CZOF3Brlb7HRv3TvHJQVJM1bMXz9xC9sVjnRPZsP2yT7Pl4mIaAZ/tRH
SOC8hUYRqL/A0K9DBhG2aQdjmz0EIViblXibNtuFG4z9sxOLU3ibwoB9YK1jbUVkb4QwIWdKTj/H
M5z8OyHuXDIIDWbwLwBFFHcFIwjBhq6RfOmGlyHhV6QUN30CFKFfTOkxw4BhIKUnVJDqaguGWMkk
cW7Hx/Fx76+tUewh/YHfhpCnhGKr9bLaJxKbJiTsvGK6Yy4OoTKyIetXUaMtwSEz0z7fGC4pCNVz
CHwdLgvavt6dxsvKiAmQN8zjI5nD30dq8J1bxOZxOFVv6lU+OyjZWA5WK5thBoXb6dwPio4lwh5c
EkBAoyVW/95WNQUElatAw3EktGDUbaUqB58qvdHkWeAnyLAAnvbdOHtV7R/jwy2N4y3ncAJLEtwP
+CIhem8gjdVirJBGLHMv5iL+20D6AtZ8VuwN99DD+UpM86GTJ+lNrfF/OYNegY7IOXyxBda05l4C
U5vdug9wUBMRv/J+G6dz9Ec7qpwltpuZZW5ECqOR594yj9y7ocG4iiiKSyJRXgAzv90NQaqnxYXq
4efOhqTh9Xdl3pPC+eBPeuFiLTLr3Fn7jvZZv+bWTqeY7+1xadBE5DCMANm3OYP0OW45Jzis6kR9
WljAIvcM+xKBdIfCjbRKkrTsYl2+820vDrGmQjzU/5MzUgcAC9+oR+MY+FkBUvCnDRExChfqNsO9
UNFjbYfndDKzaKKBsS+mNbyssiI2sb8M9hgtUnQtBOMQIgI9Li1zMnwCbkgiZEn+GPPwz4q3pq48
L8FRLmtSJ41Vlsbc/snzVKNQAcXFh/j7/4BPAsv/aQ0vTSLCDalaJk6GY21RxRN9Midfw/4z08BL
NG3HeNA1syYRJqwklnXWsVxgmU9HyNwj/ORwj3+XuYywTQhjVMGsQD18sxj1UJO/8i7bt/glG3Lb
3VsG1ZAKldgA2fG4J75nleftjrexeuc+1GAMSZYP+aOlcYTPE6T4u8hlEusWhUj1u6H3AbsZY9qw
U7P+UUvy1LHBFeZ7YU9Wgj4sHGOvEGNMZJDKruB9AI1Rz+//+Tf2kL8IWzcOy8D+MDZEWh4JrmNx
rkPzudNffb2KCzrxdwzakULFWapNGE1c+7ezTMPK+d822whpYUn5ZVxHiHXKkaR7nK/RMPiTkTUo
4jeP7U90An72SZgM4HHPJkyxiBZhI0pMoORuCM5RfoTAif65H8QkJ04wGgEg4gtj6+tRG9eyOb+m
nOgxCBrGvxFWkOAggYI+yHWdiMHfpkAuV4RAeNJzD16H4ECmOB1rYr5KuvhMobgOg8iWBDGsKAbu
dyWDYdMpGWMp1UPdJBT1fH+zC39z13ULmy2e9aJlZOslzzcZpI377rgM8oWe4Jt/TuX4rQI70sHQ
Y3x+yJNUXidgw0FIeE4pM1ivXTe0yxh7N44fFAxfGjcbLrIRWBSfC9T/Ljh5OLnHOb/SRUHbrMIi
tP78++nIvtLUWTf4XSVO6Iu8J8DewYk1xWCZaaLePpS/0v9Sgow55oXk/9i3jrfBFwHPdn1X+GVW
3GODZ5pKoreyJAoVqa+mGwR+Ey0wVsJoBAK3/VhSntlQgv5CcaVYlXxAqZ8iEcnBp2sM/MahtVJx
pu3yJVMBH4E4PNdlQhUOhOSt+ltkkySsh5arQZtvAwmrDDFyhI2uqvqiEB+lEKPA1eS9loR3x5U6
lMx7q0Akf6yn+UJ2BfYOGfbYD0l99PlrTplMNgOqfw0ZLESdTAFkNrtBxk05Mb7YmBHwPF9wZbAT
t92s0N1/qBu9md18jz5TO6bXKK+88Ves17EHNh0ePRDvRhLpTUAELAuqqw8w319yNSNHZ4hfyxrG
YRTy7M+9tOQnplMTTOxEUaVyoLVF/CifflBWEyaMbGCeOGOEcQnHuHwGESgKv96yEHMjprbWM6Bi
XDftRZfUho/yzhpx5ZmhtZsHVLVZD7hH5Ufg/NcEIF1HR5Gk1IxfIqcoy4t1ny1amVKosWX6NEP2
xwTHroGHFZqfZdKqSoYckuy8w37CPdc1Q/JCUydXag/Lm6Wa4mofe2N4IeFeytfw6NibDq3dACdW
7puD9y1xW7FAWLJvkyUkXd/v9csoljhjGI88pVUTCxJeN0F0xjMnaa6YTqVqUpHmLx6c5F9NEgE8
VznaQtQ3Qwf3D/4OZaWKUBciITJuTA6YP7y8pp8VmUIQsTSHqLnWgqQdZMLV4k8bx2K4OnFB4pKR
fPrW4yrl2qjAiebX/mjBQ1yLpQkyDvrxKfeUVnlW+EJwRCXR+8pW+0+E2kWDZrmqpTO4ZT8n5x4a
2y/8crfWfMmLysqytZfKzS1+Gql6Bvh0FuwWMRvDdsHDSlY6rcKICpL0t5YtC0ttLzRf3/IY+QBw
ct/31tw+5qn1YEosyPuWVPk4Rgb3jG1Js6ZKmK2E3W9jqnDzVxtcgrShXsMsvAF/eNXQEWFyBaKi
nSKiOfNoGda3EZWuDMnRLFmENVeyCR+Ir6wG4ry5+orxaFBWo31+BZRdYKMB+dQBLTWX3ojgfRyi
BU6H0lwm89tcqIqbkJsxV61cJpGG/CTQUIbIac4Zhwo+utpR7ZcqHqdcLpgr49NFc3RBYe1kF7+7
FHeN1+iLuR8gCpuvIjr3PeahtcmMXf37sXXXDguQ0Df1CJmgAarEyaeEsPmtPkTmMVov6MXnQL3a
w0QPtaETkDL06cCH1ywr2dFINa2+9H2UAbXZvLr5AMvocs+qmToR+qp1H9VSRItPwhokyBIcbwio
E/jG8+P9IRNmbxAa79Eu/zguLa1fQkSUsop54gU77uD3yHcCSInf0fNO+r/ckLZy7rQmwPhVCUdp
+hys+RULpsTcUspqjEMIjwAPeCO00evmVoXkLYVBdg5Izkuqf6Ygmna4KWx/CvjXOnzedwNb4hwq
gj2ljt8Kx0pgtJIJzv7OplD4yzl8VjmppdFoXMtHD9Ob+os1wrnW4NkVogg0ukTS59fGN5Afz/bS
wX7/kBg6uq6zq3z48/lmuefDpjKFWDULpl+rCfULYA5kfAdOLk0wvqbxJ8NiGVkLmL+1MRH8QmVf
XYeIx4HmKDtIsm7SW8NPCdNaGj7v8vhwOB0N1zAf1jlXNnYSPcT2VZdL18dB8F1xNwKbiafpNgUd
nRkr5GunebUrO4L3THlSllicF/fqAmjForSLKEv5zUvrBjHn2CRukNrI1SBLPvf+QEpNhHgEX1qv
utl/PmRy218dYR9eenjNqLwLyb9qascWMbmzsaeIK3SEmbAxsGM3GYXgpz4W9KSz+qq71dj6HJdD
8VJsjbcZIa2K/HGs3Fpdp1wVF/dDxOVMg2Gw8Xq5KWtcuAbpLmEudBJ/EjQhFFDxzJtkQ0ITOaK5
rw2jgwrpS8FSqLA1BJeDyg0oNTjruoxiIP10X7FFy4rBpv4QIvXOZqt7u29+Az2uFk37RG0KXUVl
VSNEfUZ5TagHTarupaxvnCzUKNKdOOLfr7z9tIitvJ3C2zp1I1KRI9XaD506CNDVHVX1oEXvsiZW
o4IxTAxdbcdd1Y/05wpwgFrdr1TXFs8GcrWJ33+XtoCg7lVYIghH5L2zmraP0L5/XusFxYHs+Jg1
5bIe6RzNLxFvrZC6+eoEwfN4slLl1r/B353lALUdRfaSX/02EGBWcz+/TnTSJnuJYR+HduZdmdlW
auVP86QC+H8YflIm4yjNtuxz6zZdGDF3YgZpa/VxCMSdaG5fDFfXkFenx3XEp2lxMVRsilit4DyB
67Vc+9uzySDFam2nzpslclRTWxjbXB0Cgn7RrXyc39TlKT8Ww8UuZXNGDUNPWfOdusvUg7eT4x8F
B2cSarFRT5zmdb8TddMBJVIt5wuKRrlzrAfPPzum39fAOLyb+U4eh9/gd3Pk8CG9mUkhgIdPsjKv
DihxTciQfinWxzvmpyaqjUBrosUd2MMQHIo+pXk9vNNILgNJgy7szBKBNrlBS/qlxYi56GIsdd1/
ubv78waN4ZcSe14Mu3GtwrvdyFtEi/vsb3g712YdigYIRLpsauLJVLf1Hg8fCkv7PEJOtrF3AMMy
rJlk73kp6uKPkq4vag5GJL2Az3LcL1J4L/mABHu0n90MRAhNZxDUzaSF7iqZoXGEpyh/0mIJvX/j
scbHp9edvYeX0I1ZQAO65EJ/G8nD59gaKvApGVZdCYpk3KDKLSPvxDkiiAUphNHoVcVF4Uk8M/bQ
oI5cKaU/ffKmfi+XkKC4s+k1POXU97TGY/+TMUNIxran4PLrr8qOhXVBgxEXhB/8IxjS6K/d5Znx
fp9ug1igyUN3H9pFxt1KNFvxknXzhhzC1mGP48elUks/yEk5xbc3EFEZ8MqKp/Y0lRgYkt0GKTWc
RF6A+uRqoisU5dQ8frO/l5Fpk8JDmKOW+YIisUFzLsgRJyzZlICuBQTRn4AlWAO/bsHQby6RKK0K
rIs9SghZeyKHJcuIiaOntTXpivrTaGA9juKH1qB6qwrXh7mBpxFghV122uSKwXnpf7AJywx8kojW
7HTwfaTZ9FT6BJPemyKw3gHLtqgFuA0NUjaXYha/PPLQYzEwEvaYSFPrel9l3VQutMXKCHK2/6dQ
ClOa/GE4JEHTTHCuLjB8H8aR5mdrga1sgUEXjbFZJEmf45EvH3dv+wNXiF9zkKSPnG3Bc4DNyvKN
a6PRgBtLA5U9SqOyM4+bVXbJYXJarYZPuh7s0Dlck8wvxzC48oXwYC09X9CmjjFe0+txyUULN1G/
O4751B9bBFhxEIPzy3PCt6KRvK0dUfHgIz2AjqOBK0Nbjd9BV8vLDHYhzWQmz3FBF+EEEXik7aZ4
lmvASaKvxYqTpXCjj8wZKP0BfVLoFHhgaUX+Vdhzy5w51s75EF9vkaSQY4v3zfuOiKL5Tv1vUQo4
+440Xzs5r8oURvTFe7DbP4+S0wmpHQmhIA06bVMKw3adoIJoJp9CBfIifUe0xTImVgREnePfQ/uP
CSefQmFSfWXf29j0avy4lJkR1TM4IGAvSW8InK7Z3Q8kgRPIuNaMUObRFWF51TIjq9ppUm/d/43c
SHR2YyQW5yS1uzY47XA/xS2vBLExY2XXmZBuEkmzkMsgqqDuhG65PxwOozKV/h78CSvTtw14oWFK
Z9BhTCaqhNMlr1QczMvwp945blCAf7CpxRtsIfVQ+f5km/nazYF7M+RcQtrqM818z57JQKxEzLfc
ldU9k84ytVcsvdHepryqSMbCGwiqV3m48Qb4z/qzSigZZiN+6od6YvJMAN/aZ0OOtx9Nlna10Cqw
eYJbtRM0SCn3e7/UnYOKa58Woby9QI5B75vj+OKiRfjF+JUJCjnsp6CcRItYsFCzYRra+YFOYX2R
oh0Au8n1KOm8RnXj2t42jfbbGCGsBbUyw4HTjYcMy0anezX92F4iyaAKNpyVovGOfNGRM4wk9Axp
76+TFciUCt1sHRf3FBuldu0Jq0N9KYHNJPT4Kn2OcufxAngq+KIK95mg7cy2Fyi7mBcbGNZigQn5
6mdfZ2rNj+ax86VyurWpx488mUoJNReNOty5ZK7EA/WRzd88XlMeHKdbyQtyjBVEI3wxfQxdNQ77
Pid3gjN0l7XjjygZYTXIKBCa+OZerwLY5oGySKcvlFUSPHbXeukQ95aRBTK6wpdgrX5unVO/qy8v
gLJuB/Td6m0QAFwOFfQofTI/bAV1/pCaRD7Glw+uXfhLASvV4qPER89fpIAEzMIyOzrJ6babQ2ic
xd3Zbe00uQQEL4kl8T/7G/YBSLhjy4vE3wr38sHW8b/OO8eejt3jo5HK6j3if/coyQIjuYn2c0ld
hEJ+YGtGO0ZTdrYT2cZ8ZGaXKR9WDgaMCwjbediQ8X47yrxyBclQNxqFhPvFQk7wD887XKg80a1U
Xd7ajqyDySqZsOJtKQYyx5gY/xeBhoXyGSozGeWh4mr1wHq60SWmludlc0nD9u9lnie/VJ8bS9eF
Pc4w/T7Mr3Lh1mtk8PYSNPjbD4TJAH47GraOmA2gQuGfQRtbUYy/JnNc6hJMSKAL4FGVswub38kW
cmFEXkrMHBHO6XEGkE4KM+wJdkqDK6IIJnYSb/vSDJswWa2hKUzP3TtBUrzx4ezCcmb2K+Dr606d
DFXQsSBTtmysR2FFO3jTV+FMnntRwRI1R+vCclwEEPWptNGSqDAGo6pDGFGkBUwFp80q8l9Swvjl
PIx3NYJYcFzQVnFX5SX2KdnnAprTtuDtqF9CNCimM5P7QTzlEFgUelVIzYekyDJmaILW+3WMS9Ir
UjfZ2td2GaElgX34vVCy08qUFqY+ejncsPyyNcfbaNe6Gx0gAcnu0cmgCiErgExk/+wCDGG91G6o
601vXD3qeH6t10kyo/s6OoXP645KFPDyl/Kb4gEhSkLAqbUS1aO1MWub7zs3PZVnbWh4fze1l6Kh
TtNtpFnhZUchbcdkJXXmFtIYdB82pPPss5s67lji3e8efx9sxfz1cd9p8RNRu6irbJDlG6G+abPG
gTQgyfV3pLrpc6rPReGNIeaxXm+x7nlo9SJcRLpkOKv4RynXH5RDYMlsgy2naliBnfg7a7BcfzzD
RwzvzkoXxT9NuH25BiAKS6beXbdfPh9MxGshqav+8Gr+RIn3VZPvrEo6hFTVTcZOQgW7R64VF6gp
GJRWPOFJXOKbMZsjtBf8I64BWskL2aikv+mXNHUzP/i6g74Vy+dgnKHZbnT+5awOckcF7p2697ze
QfdnpXXPI5QFgEVMKZQHcjWKMxhJ6J8LqqgtnCoJcY+G1Lvv87m+vZuvHg7D/iyPCvswrIHYiTBA
Q0K/u71vFZAoDBwhuODcpc8Qb1k/JRKazFugJ+XqqolMhu4OuwUbTpbljQ28domr0KowXK04v3U9
VWsuWzEoErf/RjeiqJFAv/RaeEPkq7mjf8bi4B+BcCgcs5ZzhMMpQ15wRBNnWjXzWEjK+9LTbwDS
YrW+H2wMfPyGQo9ePP4fR2Y89euMVpSLlAfNv2JIE6i7uR4e4Usy/ZqAut1HG3dgAw3xAIVjxDZT
uHWVo1madpmlUzNPc6qVecROW/sF3Y8Pszh3CoFgCSVX6suVJriZCZxQvtU/1XmnFL6j7WsaHU2H
QnhhP6KljPPjWDtGyCyOOkaMW0R6fa4A3m/XJes83N0/VLiWMUQCNC+DEG6X9qNfHMPyWVdBPkHQ
Q6LSTlF8KznLhN7EhXxSTPKhhItT7a4BjcX8K9cYEc8tE7s/i/myc+H/5Kn1u0Fvtff1sxIRXkkM
Gv4jkziU5wbwbXJJONwWnhkoZQXZny/rgP90Q88FzO1NYG1QXG1dqpW+c0ed+HxHISvll3ul5yJ9
FyfbxpGQjuBx21Ymyr13zzdrwFXEpon5kmc0lBR0lru4PfBdEcNcsND2DOoRHa5Khe+VPwjzFMds
fZT+5pwrHxrV14FF3jPrTUo/UcIRv+ZQiNVzrLMP+INZ4CkLcoq1dfF7fvsUfkl+MFdiZrw9y0ZC
v8k26yeA7fZuGfXJ5bR8YQNnVzcFAKxaBKlmtLKQ4XU5RBwGyTcb/OOtyotrhKaz4UMyY1XCO7xM
bCLY7UL4rFQEgX37yto/Ica1YZ7qp5MM/FDXsoJGvJtpgAI2Gd/dJLGHZ9HAlWuJgUEjfX7GBVX7
LJ/uGxltm+DIPrcCM922faY0ESt7zlVfb4eKLa1K/clsR72p+Yw6OLBf7IVWSqxqxEJbcBdMV05N
qFmZzpR1yIPgSyxZqcChHwsVqoxRxwMhV/J3UvIArN9toVu9O9PaF+87/o+RcJemiz5HvQnGmyVv
GNk429hGTdcKKTfUnSPfDLwcH6DEVE6cv1FH+5NQ4+Y9DWUiUBwM+AMepnvDJ+oPZukMTDfJsOih
lW0j3JDPonAG0xPkCSTxvKOUqwJpEBmty0vfg0HobstkoTsYMh8ysGipumiVPYVuF/NJQW/rIm46
ZSOJ3711hXNEN8wotpqOU4drP2VfOmPFzdljtMuoWxB0xigLS376bxVuECTTY0XPjxLGx8Dryzxd
lwdelIJvPJkzgKECSVkLq0IB5rEx22GTGeXpvOfoIiBy+UCESm6qzAcP6Zw/C7KX2ZqQedH2hBRr
ya9eZCQ79fLUjh18fFCmHRG/n/QMJYsbrcBoWNrGUlSXpnSc/9k/FpoB+SFFgG+um7TrQMZn8l2e
/tdaFKtgAYbgwuMRAfuzJ0Egj74DRxxJbTsv5cmfQZeGnP0MXzdzPhtFKnIs3Hw5vWVu7Bv31bii
5LhtxKbvL6CnxfWWo1FWp23VBUjzfE1KPxA1P4HGIvfW4Mc3w5dhWbWLO1ctc3OXbhLqxAS0nU6X
AiQKdLoqL8/uqiy7hIIIaFI8J+mGK9Gv6Y0pTrPETlPXfjsT/kiIK+Q49dAogHH4v5KH11i2USIK
3pMe0aTfwzm1/NyApKzQtKVxzDWTPGwA0gJ+j34lXRgGmKE0MaTdCtqvW2OALqHAxLvec4tTJ24q
Jmjy/qTsz1UY2THJ5iLZq51R38oMx2nN6qTrPvpgSXC6EVflkKwIRNzYfEkfkSXpvBVWcxHy3SfV
kF5dr2ckg1AJVfnP85g4e5iyHn1jDmKL0rUFqDxzzhIFZvdDF4pdd5NdWlFepP3+vtqvehIsmPJN
yhbNhQuzvrNSM0pglt4IB7IfxMUK6niPpznr6NbZm6gWiRXXyvfqAdBhoW5pwrQTjgJqD/biTcqz
UFTvYd+lZPbgCIcgAfefjmaV3WlUxDzR9XbAK48WeodcEYSMxHfjbBoIwSixmFIRm9ADqar5gtU5
wTFdUFaZKmTq37cbvLXF1uZS7BuLwAcZj6NBwSBHuz5iyRBwkWkeoOcoPGdYUU1eUzq+hNKy/Rk5
lbiOBIkLR0SuQyW6aKUpAcz101kQ3r3hgCWYH89j5y+8Tdg5GNVX/7VFtK1180LQZClzwRraln5B
ilUfVY2y0AGFUy6KiOkSk57L/ZXnpIIECWlWONv6kTppIGd3SJhPqzrmk1iLEnQ3TZ4dRuUwyspZ
aPuznWRc5RkzKRZaSaicTPfyJ2Ml9RwHcd5+MBDzDvn/Gi52PsGtIIF3F3gPSoH9qFGAMDzuvRFT
TL1piHvYUt9veH7HqZ9hlHZZ4+6/xKWvicFZlZzcP1qLD6ugFlV2n6gMfcmU7iSGOFY0DC4srIS0
DDv7qYJPw9p8k82dOtEOJrjVtS5w6v04zjXtE0Oi6B+M0ueHHUSi6Jlqx7titwl2n0zg501nlPst
qUKEfY6SKYQDZ4XI5gi8eXAQzgNnzUbVJ/nnQM2WHRXLk+I6QZoo9xtcURUnHYIIz9vDZ5ZQBZGl
o226R+OyXPcqjfYWWAopkIfm/Arbm6AFSsbr/iLx2+9+cBwDl4NiwY1pxP07hfeflSMujsRgHa65
WeIqV1Ra0xawr5Xq5PRGoDteajLu+95ud5kAQUnp87DDNz8jT+9eMiM6sMa/4kifYRxWpESloYNW
tlVApGHSPwy11g2i/Rj8cafM8qot39T6p0G0PHRsV9pwj2wFKAvW0RWffU0dZIsT35t8YxcuvNvw
vfi5YxoOz3RLijEqF1cuaDDBhU0uEqi2X6w71NV2DKFSi/rituVmLB2qgBp8YSi97lOCLzF0ND5Z
SU3ST4cqe/oVtalvnHc2jWL2jgmSoku70amO5bMSEDRRkoLGQrkH/C5n1PC3SJhvFkpU7D7L6IdP
7gxRfFNglYiLdjtKfMDKhBUpsbZ8vhSl1QlXiYYHeYlkd6h5fIsntKtJ9+lac0g0ioDytcuX6khp
Rf/9j17m1jSfV+vspNynnqbldoLCGauCe73p6z0Bi3gixJD7wvclgm3yGrjhJhd+sj0GnFCjkPZ9
l9/yQ1iJazJn8JdQl65ISxSDK0GCbL4iho6bFZTQfrwVCRAXDGX6+LWLJfq3PNhwetpZRo2nBx83
BpBJxJrIH4TQU7O02PmzLT7zpjg6U+fM0GPLy8B7iu3THMUGhc69YvRfcvFNxwR7lRKbmMiCZD/e
dToroJOhaFEquiZ9c5eR0p5/Y7aQBRoVqf49zCCTFUhz3krJSwxa9DpcNF7G5otfxySIY9+kd1Xy
KoQ2SY+vLmUVj5R1TqGI49ZUEN9ZIAOUDQ9p3YnzvN8Zk5zyZSNZP/qgydg1YSMRQs0RgEgyI8OO
nSt0xwKUrdHwnDbQQx4Nu+bBrxmjHqEkBRbV81r0XytZMZYvj/doT0TE+/VrRYkieX36L/JIBCNG
ScEzklVUckuW1Q9KLS2Ar2aT+vXow/rqG2F0F6f5xpi3yjYQRZT2nAuH02FaWMdH1bPNFDJKfJA1
qW2ZQ/G+MDNPsuWuZuRQu3y4yzb93nt4yx4Z0siqFCh52sjMdmjkjVWrx2zCRrhBce9ufXOhqVSQ
MlR0Hmn1IFgsXhQwR5F3mEPsj5kgjbsFpuMKmZykxLsq2tO4TXd76F3XCjZx0FgZN+CFuEbl8RAH
Ur9LgAIQvDNeK0KvmtHWcI32zKcETP24W1bhHZ0twcsq+OTXV5s1Wkby0vva29aQ2MAZskshgAnY
g/phoscPUcn69I9BVjNRcY2TBIi8U55Z77zEZlk+mVk8KwoWUslkfZ8W371yHm6mOSMU9HxPeePd
Qpq9CCPe3dtfJkl+itxuR8IBnzdo+HQ/ei4ZZJvLdyI2EAC6XLlZKCbc/3C6bVv2DJRmKhCxqBi4
CXSlCPGboBq4zhfJzjxbXMXOVjkCn+Vw4CI1vE5SOTrIA8vcdMriCKsVZkQjoMbDhAePzlaumr7X
3kGAPzbf3rigBYPgCWLy0cRVXx2/0E2D2unfUcmFG6dTdHvxCk1FnURe2pQ67KH2La0eV2gBWNgk
l2Qw7TeM4hM/hjOlaSz8gkXiL2+pAkxrZODXMX25Vk1kk1OEmnVDVmXVSVq4bzl2TX1wq6b/fUvK
fA+CwiqKebKQfl45THs/f8aN4DnJbJ9ZgvYoY5Lu7R8wBk8LvUnkw+Ubxz9v8s6PPhDRpD1hznmO
C+YBDtA7ciI+tyfxApza899zgX3KofKTyCnxFAzs1x4TXR0u+sYDID4K7Oks6XhtFkr1tO3L2ece
2uezvRFTFmwwbT6MpLoZsLQuFUZgghSDLNq7sLsQs60Mt4dM/H1bBYReqPs2xVKpVbjuS1Ov7/kh
DEkpdw4UpvrrTRSu9pA/yQkCZvwDOtCHY1qCIGBcpRH2/O5QgD1k0gi1ukYJL1Ifp0J4K+4v+6wa
pYJVgwm4a81VcL26r+VqLdvE97F8VIoKicdpaDro5ZQ6LsUB3nImn3JP8EcqqpULMjWFAbaY+6ZH
RXdw5DdEYa4k7G2uANzBjOfLBrHkG+mJiaSUTdngh9+Rid3VofEQoIgjI3NxGHei9DHo+8sktb5C
XuXbGWbLcUlX4Cg5ugL+wS6hAj0bcuB0G4XR4dA9uS+OcJoeu7EsZtrstU6nLCsRCdKUR0yXkCQS
hJZeL9sKVVYLrZ3NZNuP9jgqgyWgVmnbw5PBEmZ6Zldr6iNg2gAGwlsKxLf8F+lReFq7q9DETuyQ
vJ+p7vOEtSj7wcifcJdR2EmW+4z6N0czDUHZ847vRNj08wldvBtbea81sctj/VcnSn4sUgBrxuBW
oazgKncOXJSKHb51chhBrrMocpoSZFEhU628kDmHv8rCILXTN52LG9Rw74zbsbjZIYgVCWXVGw0Q
4kjjDkhuG24udyANA9fNaq5xaJLcKdlZa/5XZv0fidxt0SLdDy9e7nlorxw/Hq0yBKQbjtLfJJ0F
vDXdbbwKHGH/ZMqe7EGf1A9/85RxO3FEDhZxgeXb4UOrb0yhfzzwvCnHC9pnyTyv3RxmRyr6IOm3
MGPJntV1QoWJDbdKaSe1vz8CilxDoWdbTRbyvDHHhxiV6fZrkmbnPcpyB7w6eTRq3NK5Gw+TgRck
bWGww3qax4ZNL+PcN3Kf7VaDkDAi0jRP7Yo8gh1hrHYTjad7kGgUPT4loAraH00zU1NjpDac+OJt
gbdQlPqlgIQpEjJsOKlaaThCm/uTdjwrI4bpKTT9dNDDuI5h/kW7gS8Q+/Viu8wlqOHI6xLuutsl
ehRCgYDYj4QkhOrd3DLvEqdgdYw83SqscitApAKC+irBXwD6lJltvfYRQmU6DjtgWHmSqDJGfBfr
YNYSlf+clTsXFdTADM5Rl4qF5xBGBCFErCsLDBjJ7K1FMxZWZKfgzpMFLxVQ5qCWus5aFWWyxcxo
Hg3el2CgaAaef4ETlUcbzOrvc9yT89v/Fy+GiVzA7kza7DvdxyW4WnYPaWD9QbtwAUPsjYlWA9ZT
Si0tEijBkHH1LjgcIdnsWCPJkwcKiKgO+9VmhxL4zfbImcplit3lOJ+0Yn7h30aatqx8+oAKYnaH
leC/9vUOPZmq7Xc2b3Sd2ew/nVFddTnvn4xUMLTDhoFt0gB5QYfGKaxOnablSTuMRIXLbr6iAQTK
LOyBny7HeYpp0mRtnihp09TOCmbWjCp5oJhvUBgnONW2crrTYLLDEKX3TeWwL305Is4tg+IXGxot
zvSx1y+Mfagj4W36WqyIkN/t2nEStjyYJajsNjwOzV0In9lXMPl1sWxryKkh0MbNAgXS8bWE6ACC
z/P4MHKhrjUy4fiXvTQ0D2jquTQf2mCeGTTxHT2q5aWc7taefjzk5VFLIIso6wCpWOAa2XW8kYkt
FzkazAi9p9dqpENYBgdhDqWIR5udLR7dDrjaQy5sRcVa8RhPewcBhYi5QNiBRtBgfCWN6ph8DBCd
oDWLYSBqXyeFziC2ncLbMAilUbroVr7qXk9d3gtm6E6EkLWOIEMzQHevXqwK3fyhmpgHH7XCPBrY
VoSZpKP1hnA0T/j4qwEvQBhhhTt/4ZEOplcf/gRsJ9cQ0WtR7iYjPn8fSRnJbKX7q4265wEWz69+
0yQnaWou8jn9Wh4cZx128nSo1if+Zi6E4mubbhyAfSVmNwgFnwW+tbjJokmmC7T8q6RIi75nIG6e
SA64LIVtOYN/5SJxO489ABH61hEt9ZFwcV0Bh25ysdBM+NdQpVhBaRR7mDgo5mjJsKXFrTM606/K
LlRz0UKVTPihmxja92joOY1lbBV3x3o/upAE/wMKXRHrhgPttzYAYPj4bFv9O+zLpoEQBzxMrtrx
mPPxcVI23UtFFr+2D7mAbXMkvCRpdznBPVhSmQP+8mtREnZDB7Sxvg85nFvtTt4X81cbs+aHvihY
krJB6WP8BjsouxCQ6fUL1G5f8u7dSEgSXK2CQlWsn+S9nfQXBAAYPI/nmg2re2HpQ9YYbvCITZom
mao2pQzAaqBHceugsU9uVZv6wq+YE9EM0MHgRB8qP13OjATQ8B6gv7eSfGguDfiWZNAbvoDc30m2
SsvSl5i4CuEuYvMLAfFs2TXQ3SdnQXLl0CKyLFrzQZEzpbjwuSFhCtHxfG6DrMkbUpSFewRUWcxF
YeoT/QDyzKfyths3OXqufhjs51dPgyntTHx+83SKbAkd0Pj1ojMz1SSgqZvAtCmncSfrUQlZhZTP
0KpAmAjOh+5i3o/5fLqf+9+siuFeAC3N7dDjsC1RA3VEyw8Ys1ie5nH8Ru4OhLE3/ZH9RG0EbE5G
70Qj2K34jBSbHb9ym0Sau2aUS3+X2oflo8nHZI6dkR4AUA0Oex/AvFZcSXOqF0k9p/Wl/skfzaZh
DiNzLRnuC4ol8rMr15O6/eYlXmskWfpl50zYX5T/BtVSbnrllCYayIK9qf9XC9gA5uvN91B/MsKr
uoAWRSsbxCaqLbh0DExOZGdcjv8ZvHVBYj3U9xsEqyGFD7qLB0EAS6ljhG6rpdiUqVS64rwT9Zv6
xKJKrypk3jZhlHvAQJeUhexMVu85iKAtfOXRixcWMYEEsWlbmolwNQ5cCKpbaYymv85a2AGAOGlz
LooCEbiRFLp0iW9wpNC7Xs3MbuHNPp93xxywePUDAm+1ixELcENgDyMo6q6ZCExaKmqc94lF2esV
ltVLBp5MwajkuAJDBWAJTHDXDFMqRw0dEzxYnMkgni88CFCLZT7lZ1RcGv3Ab9apL0sB5KHU1tbx
FQrvvmz1RNQds4SkCSOUBITvCIXS/RLBE5wZnArUJPqBfeVqX0SLin7XPt3fHnzP9uNrrQl5Cn8A
UYhI3S5Swmuh0EMMVCzzvAS28XmWTlsNqwU19DlJqMqhVX9bp5Ah76nLA4kVtIVRc4n9YeEhmfhD
+4Ao4mxnGzpyrQnRaOkf1yqnwLQ7yjD72m9K8vUttWpH/Qme0v3+MRAJXt6BHSrFV/0cJr5uHe2g
oPp7WIUYSc3aK/mCm2HsthVhqYo6zHZC7gxCsxZbhGHNmIdIWg7nHNVoB10KIGuG3fhNlzlB8XV1
zcZM3maXy4b6GUBt6ZcxjdE3EVcfUDbOqonXljvKrsXfyIrWqw/0d/CjpTEASr8yJFoNrG1R0cVw
6TKIMWfbhGXGXvkZNQvTzmsj1rQHhoZK3JR9COkXtufaNqPDdYiNekzaUfmAcu6msSCspXyD76us
NEEke/IofvYizbSHJ9NFYYVKfZBVcWBCh2z4s7cwH9xRZMy9gRdA9YD+H8Il66LbnlGC4ThcYVLp
/pNW9NRXjfUxoWIJkMQVlqmZVJxO620SLO9vITQ5/TsE0UXSDmo6nd+MupvSNtHiPWmaxE/QSILE
3StSuW4cKBxbbURBbqiYPjv6H0WtEAkM+QyFCg0+awDVgYmQJokg7JXHCUY5zy2bE4q1kHupCWjw
Y8TrNra6bSOMHnZSdgtr+k+PBzs0RN4YsKqYZCXj5x/G4La2HiIVjCZywToXP9yUpDopbc3vlo+S
NTHhs3eXdV3gDJYqXleIuMV8l8qLg7ZqjiS/LAS1+dLiBoZ8fsoId2w0CnrQ1iwJQUIYi2TA515C
yII5dDvpu9NpEPYmLQ6Dve2krN2bGx8YMOF7uh3E30ubrGig2/LVuvPauOVbByzkjXWGO9r9IHeA
6tKEIM5RCfGM0VoqJYz0YQNI+hvXGuPmD9BqV50Sn6BnhZ57vO2tgvLbGPkZx5biJ9E0/1pR+94n
seDFOfyjAmXP14a1oPu5WPRoReKPaYG3lYqEvCzk4KNar+dX9hQIKZS6o8Bc6wx0vrbvI3PyLd5I
YAIDGdKI+AD2iYqtFh+/l8UUjmvK+MQCpTcgb+zzemMx7jYRXtIxRInfabe8arBHtMhYksWIwG6s
AQqXojy4B/sD8WNAEpT4OrReMyRT6fyUb55KW1K6TiQEbc6pC7QJxrYWo6cuCvg9zpAd1ZTpa4RI
ZWwgqSCrIJqFBcwLZVw2Zp4DYjDtfVOUDH2z2b01OkkN9iEwSTxBOzxJhP114E9hdNCl7Go7w86D
yFvmExPmmmniX2aUtY8XYD6ZEt29JJXn+qOprMgDaO7NHZW3hPHEDSN4+haq02/i6ZhBndXM3LIg
0Zl85idW1e6qLPvMlPrhyX6GZuvhSW9KkT38GloJGAYYVhd8z3o4/sCr5xWOw7MWqKUGdJYYfyNv
S+Z0htV90ZC9Uj/XJKkzKi3kn4D+EXkPplNV1Wn67nfK7NE8GrbHXI3c7PdKZ+txjfeOCgEZDP/H
rKz0r8KO/On39PTEP692L5KKb1sWSMp2To+KiBfECSn1VbtG0sg3IXH5MbFPNf84JTzS/zH227s7
PCr/o/27651xesIzxIHkH1amXbsnhGEuXyZ7PRN1NqLRhSHYMU2jfTGHPnxOoDcLgZTS/wyQrLdc
xQkePZvuk/0oyb7q05GzdaVCNFlmlMnhje2EJX3G1RHLKFyOVPdlUHtgB59HnX/hAPUuy28K1esp
/pPwpU625/MW3Pl6krGRLw6cC914aM9cDW5yyhcp8qi5gRPK7TdNF3halkQeIaOezDkJJnVxvU/c
jnAbEQK9bROPn1dXIRwamXGSOilNlEicaJvip4fyZ3LY8Z60rLiMLMqi2kilp9WVD8xoUvC3Rngh
eAFqOPw9LRr35u7mRnGfEmw0M1NyE4uer02zJofUT7eMG1e5Z2s6JrcKDao05WPjCGBrq7yEMtOM
oRVmGPEdKyq11+iRHs7y0w2IMVYGbA50nMtNB1vxMRvLnY2je9TbwMH1m+BN0P1vhiECTw8NlAmi
Q6+oohEf4bz/oAHD69D6ofmEM7BblzoOQtNc1Dj+VT4TXM4gA6+UFPKe2SdQZ/KetbtaCxe8AB6f
ty2tp/HWa3kc//jrTxRoQoXiz38pW/mXaVtUc/rjlG/Y0lKpbLd5Gx/n3hr/DmDk+iP5vSPI5p7V
pHZSFfMb+jFxqxMQP1GInvHgqif8e4FHjUK5eUaOEdkPMW88eZujLBuVvhcQRXS6Qx3H2Px6SS94
ZiDVQo2pnIsrhj96jyGqs2KfP9Mzq45+VZMlkEs50bAtzFSm6qWiZNkW0PV78qanUXCWQHUJB/gz
SEn0xAfHSICIKbN/bpT+Haz+uIsAtQ8sq9W2oscpolZ+gDW9wzv4fHVb2Q2YmRcMBN+Zovb5MDpq
PqBxxoqjWSTReWSZHHZ+cegLowGIxxbKyXbYufAbkOJwP+/N2VE+/CwmzOqsrbeeCeD34mFdwJ/C
G812naKY5aCulEaY0NwKi+COaWc40dihKqDBantAnlhbAFUR78/LbOJ6pntFH2TiFRQOzs9jc86A
ptG/w9AA5U/Vtu2WgiMditMICYOnPxfYMo2rOUvxFPmGrhW8D66FP8Hqgv7kfzUd2ERaSoWQily6
wWIBLKz5IJQUt6GILnU5GqOhvt+JlkGbSz2zuC+P4Y90QCnUZWxsCnzPLo0o3+q7h89mh08ZV64x
A8MViBVKMc+TCFbBcVbqd+xLNI6cZKmrtyNKCuIrjqPMGb8fgJuNf5LIOJyXrezPK6T5ViKWbtEv
+N2T1hCIZU/Jewlm2q7J/Q/moGGHopL2ROSuCyGMXK9vVoqya0MHv8jU1DwDx7Nl2uMk5nTQ3Wwa
218adizCFJEqxPydRHL6FOOOgoJT/PaJ5J+QrhG/dtiSmjCudl4PcG8RInxe2ChhV0+ciRVzyVec
5T8ll8hNJQM/gzCRokFoeUtHjM37TSjWlJ+mz3BluDjKABQ0y98vhP6dZtdUVhXrM7KMITaKgRz7
uyCyzLaYpn0SXSsaSnS3PMYxaiybevgeqWGvDAvtPw+vjlnhB6uqmJlpqVn+asNnamCFnUq78N2s
sJoy5ZoTsET7xbJPeannpfUwjKWr6eqVZanpFDtNbPg0lU0hnWm5/qw1xnaX3ltn34pzh14KqglB
San0fRIgMNbPmbAk+/lHQcC/cAl4z2fH48AR+LvD0IdB/6yR7jeCpYt2XeGHF6GI934z83KK//mK
w0M9ABUTABAQb+IwBN4OJ+vSUo2Xi5qNkYZcVE8AlzqpEK5FWkjmRM0/aSAzQ/zxSLty8Id8MubB
qmit/bOZftiH87Z0Ir04aA2LjSrwMyeRn5t30JxtDDhJcBHBRDXYX0aF1/lgqgCMm03vNQZ6KJBc
rHNWMMoe/0v3FsIvPiMDHJwX3XGcpkhgp7TLEnQw9wpblJ+xW4wxVM0TA24vR4FWHDEFiednVEke
AGL94pge/NpSmdg5azGIGgjs9+lcmSyAfQoxQeGOwIMoe5aukLbXCE6P5B60iZIWgVKwtDwRY4Zq
wk0uNRilDrMVRcySMHTDWwLyZPaceY00a0LTrK0HhSxe+txLTDqc1gn4Djg2ZWnO41BaeYw8RsyQ
iOKyPAqdlcEZG5/ApDlKDsSP3zgYuA95AaVWUvSP3U1xJpVESfvcDXcFDadrf9S7D/K7pJSL8qmZ
8v9UHw5F19F4s2bh/DXsEi8QAyAz41kPPdCffAFCEmdU0wHVjkunFRiUOa7MlKwz/fWUVxStkX4p
uQHaJeo9DaeZ/sWiBRt0VRtR+CnQ9QOumgVEp9iMCdaYUiPSnEwsUs+tTsy6VJNOPU69sIBubKEP
huMazGrrRGkeA30LnAKc4NccwWv7Lr0RIwz3pq64ImzwL5xF/A0NJ+DI/JdiouX3cLgHzHITleOU
rEAOZD8d/cwXzav4RWU6B7UNz0zuYmrWfnuaiS0hFw6bgmc/V0+xJ0kC2CoJloQCir5U8+TQRSOS
ltNdviXxIFsnbdwcsEYCOJmzL68pBaUbxOe71YohNesCQPfUz1hIurqjlNow1MFneBKg+nmNrdwX
V2gqN76bBZxfcCanzmgRF8qSMvt0dZ7uyVFJ8xoUVRxQEdfVQyTbSSEdc+oZvLqRiijNk1JhF8Ym
qHa9ZUwTOyrzBOsR6cwa1GaooFCbXCr5IPUNcxFzr6R+lJba0zLnzc/UnKqE8HUmn99uEcM7lmfe
PnjNBKo3FQSYVT4tyADONKr1dpPuSYVn6vAAyZZy2UY0eROpF7vAzHVkahK62aiGOp0QyoPggzyV
gFwaweJK9n3Q+/smt1vr7duL49jHnSmVSH70914lmNo3bIjynXoxbemUM4ynzjn/TvaMKZqX17ow
pwlk1JzPcqr8r+q0r2HeUkE8SHUjBJM/aef/hxRvQMWNATb3ulkmM0ls8xtLVYd93A6dqDwVU7nC
MlL2iACbZxMdEG4RG6lZXxFb9mwUU0wxlG/nOE0i/z3X1h4uU/gu4NQkgEbBECnByLLvCqkFNl9H
MtPB5BU6cev6/xoZnNZk3ygfb9UXNO6BGm++QFwbZMFev0EFIBPpQjkRPndtT3VvB21ocNTksE9f
Lm24KlfVnI2oTj51CI9egTQoabWPmQh17c6QQ6bjgXLCQ8kuwfIa7PO3daZayJ4MYG034mTotNYZ
ByRB3viCRkoQ78Y/7CMBeVLQD7HHyMSEKEhcWKCWLrWFsrcPbfMnCuDi+/Ze1HnVmVJl6uAstGis
7vB9foBY2m/mQfCy51SeQ1UR88rB/9N7+Oti9R9lgEK9IgarPtHiDyecWchBJ++Gf8VL3GzvONbU
8tBSQ906z58D1Ki0lBV91xvYV5FOK/e+35lcRBgBcCWtXrHhb9VZN3M1k7bbSrxzuRwwI/R49Olz
R6PZJEvd5klusL1CqKBI3npvohS/K8hRDdtHmKhsYuslhjNwhEavzSjYLNsBeFtMgjNXP2vvovcD
+Cmjh7T/y3lVjQXH7WM+bew2HNeq0RBlXWtjsaAqdxMYJGuY52JE+ulZF7EKhv4o4U3fOh7jOopu
z7ur8LKb1LRomvd0zcddh6fzO7Idbb4ixrklpgVWybdHidxCWzmZEZoBVI59UPZ5U7cOqVObU1yS
ZD3sExRPdTJ/WyTG4Ep7eZ1wPnUFhFkTqiT6WFevcDK9LgpqqqSh1azaFw6ucjslINp/D1RI/5CF
z5ELn+u5qwlNOgi3zzCan2NZV0YvijgXPyigvTW9oQPLrUb6ekiSU3zOHfZrg3Fj7yzGfrmoBIAO
r9g/c7qluN3TD5JqrF2kGETmMHwQJXIbuPI/pcJPJh3iYzXXKH0Yy1vDdrn/E3lYfEB/0xcpzxik
F67lne3rKMbjkf44z6dfDaVF8enbLlwhH/DK1uBnarJOwTVIiuUoY1Jm8JfE497Q3sCkOfbT0GP3
Mu7iCpwhxi/yt1DiIBwC8JY91KjXCybIQpUSS9Ljwg2nD1Dj3n/n2pm1dSOLIjhRUpu5yEe5q/gs
8wbLWoZwgcvq31sPTB4Inre8dFl/OC/QF1kDKuWpjqxj6kTBeBTil1tn0I7uL5cjrNTsA+Bd7Xg8
aW1EAdAK7gRsebq4X8j7X5aS9bwTcsJlAHdB7jqM9FyuIrQ5OZrLNAehhyZSK1aHhW813AtrzbTf
kbt06g8XDKNz1FwUpsZYXic3UUYxktpAj4/DDGqfWzF3g9qDzLTbEkvgM1LPTbCuNaZB2E8Rpb7Z
arococWmJm63N+BS2SRKcCy3e06P4Z7EmG9vGlnAzE23Qc85T38bAiDERMS06V9zuVL879cdoaR8
/7Pb32eY5/LvBLxgKtFVIuZfkM+Wtxgzj9Ayr27li0IGev7+pvyag7xc3TopDrAUBkW5R95USsud
9fNgNmOYlh4PGEZGktMAA9ZL4+B8iYUXP0f6zVJmjkXP/gP5ejM52Nb7krFNuMzGtXcibRvWnA1d
RnEue1A/xCjvUg9vW/c84weeAKMIGTmif+R2Zi4+QRmg0J7r2GPPlU5TOf3Fxq1cdThJTIatA/I3
Kg2JKI2uK33J1wzsVCdbHe0In9YlNMUKtSazIqQ4b5ynL8rxA69u/s+dh30DF5HtNzyEyWo8F5+S
9c0eX/q8nwn1GbbHvsCueVwGGHeK5hX1KX98W0ENgrdTLtWAhrH4piZoney5HK0tjuH9+lbXPTAT
Bi2WfT6k4RATQx3iINgn0rHv8MfkYYCKkupoXshLMZigzYW2LGVJFXeKCcxhgrsRdAdPv8VLtdDy
iU5Mlk2HPCD3spWT2RO206mTDmEHCbXUXTYp8DlzlKZ4Nqj2v7Pw+DejuRvrh9mnu+SSHxHuHf/+
/d9MXyyzpquW1cQSGEv1W781YvE7VpwXomB3uVV/AUz0VO62pwE4C0UW+Tc1hbmv2uz8srhl2QdE
1vp+3CoHRUownv8qqbelFrj01oi9VQMH6P7RJH7bMZJTLrU8BN+lvZHWPYRGk4ZH/KOwUXMuLSgV
kgKUGAtt7kY87ACM0WUOom09EAD1tC6BfcjPLq5B4hS5chfUYyq8d/5ObNuBKY/LZUoo0uHISQFh
H9YCfUUiTQIBuAEiSoZLsBBJOvuJ73D+R0a7c8oLtL4M0kRfJAo+crxGZqIpblVXs2YLg660u2pk
Z5yiXC9Wc2F8X9GCVNmWt1a41zfMJemuuBU7/nlcOaae9BEbvHL7NgbfY5v5TKs3P2tttYR+aXjB
dv7nBECOmAoNy1x99p7r/KOVe8bHzqfXWIC1rdFlKKTvTy6PoLhGBPtFWsEi3+L5IoD4ngYnNtfN
2qhbaTz7byTl+GM45ODGOurE6ko1rv8tDysaMLisLbj8l1dEacokFK9G3Iz7i+g2JXQBwGNkrZVt
FaNTKC/lDBkSxoxs5KPBHTLKVpeIxgZ0J3hNAvZu2k9ADmbnxFQOW+MDd7WZpv7O7cDaI3o0XIFh
8NeOhytIKjYH1FfaPdAyMyy7LwJMlYHkUMGQOOFrlbWsII+YfKPqCNzB6Um10WFNdE5t3iyXa+EQ
BM2xmDFWTl9tC4Iynk5g2lHDWZtGITJf+M+PGu2Sz08Aw+3j4m8HvPJKxh+kl6UDUTDYhXVd3Gtj
5Ibyoy2mYdHquUUwPmc6lA3MkQTKU7wawkJRUaoefZPTtJ6BiZ5CyMZMK3SfGlru6/3BZXREHAgI
ATO1m289siAZZX1iwe3xuaJJm0N9igZYAlDQWzjT4gReRcCaJiXYoHylnHJXbKRYy/8ikaVRVX8v
++5HCrBj6mDn8CAvlY/zcGusat+drWu/MBUg5je+iwfzrEGANlx9eq/B90FD7s5qWu+iFNUQo2s0
pi0dR2euEZhsbYdbOqLOjEJA+bkRqYFOTysgMkInFvQ5A69lUSSxJaBkrq5Ub0SN3UQVrX2o62dR
PMVR6tz2IngbRCLJkB8WBek0iZ9kkIipcgRjfHIPhG6yOwk2NLjw/hTn0/QQx1Bg0W86xCfp8nn8
mWAE/oUQIHwgmuXgH5Efu9xKRtb2hnK3LIP5u4hIUs92SPzJZHRTFRuTPkGU3NbI8s0a5XFO8dnM
uR56trrJ6vm2Zd7FzxCRiHQPJ7jdsK/8cWHESsmCv2P9DzkQjrM25+i1n7cFQBGtyLuGWWb1foAB
N1f0yOl+F8Q/JFTcZTt2WHsIelKCVatSDBusPz4zMI7CKJSg4IX82NwN76g9UJ5wGqSozfgWO6b1
xHtB6dbVv19/NJ1VKe4bWWoJXhP9qu33/KL67PhCR5Jz/J/zKZLUOugY9sC0NxXKSC9OPTqixWOq
/OWpOb8koxD7PJobml7eOxd1xE21KXZljkF6a6Y7v6sR8FRMQv7eKyrRsfu462pO9gyOALJtR1UH
K2G7umHdWs3McpwIHNq2knCKIhGyGH8L+4jMVbdGYnxlkDn+DPNKWWK4uHandbcY+2bHeG6SPf9w
MhjmXTtw8PeMF6mQLkkCxsp+tCE5vKd5JKwCsvUBZ7BnckkNceK6x3VePuMJUPTlgpuJwdJ5dgzZ
MEg0Nhf/j/UrTWlI9O4eBnhTAxtDhuyfjfK1ehL2kNMOwqzzs/o+lYz8N6ohJnWKkHLz1okJRbKG
peewmbFkD8C45p6fv0PVsaB9q6TVbciB89nTFErIVFChC7qcAtEXjX13TK8XvP6WpkIcBUechcNq
yTWvvZmIED6gc4iQ+h+6zV9CF+6tsmbzazD8n1Q5MWE5XZkTAPZEkE3qiRrmu1xPZyWszqeUi6RQ
YGP39sxyH5CQvNWlM2jKizJBp3OS6fIyqvf1MQttMU4dBoU5aaXJh6dPzPiF5e0JTWGbaJ5KQYO9
aVVBD2uJ7NQDw9HQRPP2CPs/ONRHAgzFxRjAwv0S2gkiqXsFj3ss6EfWXwGroHMWYgrz0saGMzQT
GvAUkt/RNxgsh/zLIx8x5de3pq2+ssUzCYuou+ALvbKp+09xXjm5C+FYFT0NrScJ3VlSGz2Og5iP
g/dWrKyGQPLxbqwNuDMx99sr4nUcEoEQcE0e6Az1/w+VbgSXTvgafb5rxBvL8XkY+Pi2Y+af+Z1q
cSSV+Mva9TUPeJ5MLuMoZIL0el07+RLe1Mf8y+jhbhhQvEHySR3OHaR9hgze76JkA5xDKVm8Ubfs
AiQYezJUNZESNvWRSrnrRpV61q6Zi2Z5acuhbcm9byl9isTbTKnLxSRRq/YlxpQu/gJtMFO6xS+j
b28XJZ2w57s45oxHFzN3+AE3mWKqwNcrNCK2vMHnCMooznfNPW5UwZX+ZxMAUMVj5BR7apm3mfYs
W0oO0bGbiyDs+8ZajKojUNpD49qlc3lF0KYXLm0Sbllb7N8xJmyzqS22OegswFKAP3oF/Bh7TK2c
vXkbRWNpFZxYQWRj6co1HlbOL4yfAdHS3Zyi2UApBizuyFrLaAwy8nwnbih8G15QoqmZUWUA/urP
vYmc1IB3MurWIJggdr4PXDOHeGjhIIouN4VmnFDNjRlnH6JXLdGqUGdJbA7kFfFYvCV6IgFsuqQz
b6/3dacur4F5aJkP/jKxeEpIYK2f8wEiz4TyYb/kiWu7gMPc4ndfqSNCQ0cRUKBOH0gGSQ0GKUqv
LCZxM+rNuz2Q7R6pTL3iuCS8MjY0SCKyzpi6aXLEAeuxTjdWW5tI6oUsQveHL8dpIHWsh6JbW27E
WlofTz/3WVmAnY2zaS+RnwsWt7g6wHMYVOXXCyfbeYnHWZ/82AOwk2wy1saiCCaX2j5CnsEpt3q4
i05bSQsDKBq6986w/6GmxrqZHszSLdF9X+VB8ycSzKdVaHjANW+1s3/0kJTOlpTO72JoWkvIOyQs
Nam8pX9iobrqdWUm/ERlhnb3gwqv+34f8H0smV5uirL07tIKnuMp8J1MriAKiZUqJ+Fu+Dh2s+U4
b4PRHSIfhUgNjRe7zac14VMa463Q4AZZNtL+KfQfUBaB2ybE7g0x5ruvUPi9sXQKhhBQAVma1NZb
vBAglcjoMx6b4NhAyOuZ/luvSM2HJGFZeUNBVrW8A3TLvAIukyJdH7AMNuL9i2GZ8N/5HCqJ1+2b
Vd4G8L64rwKnxKqWon8SytJdAG+gvVnNsIbI6sPK9fUHZjRPAdsaipL8kUyicrkGunJ0yEn6bmy5
yRElLA/Qw0AHrd0JoPuqffvmD0RyzKsLUf0hFx1hHv701vMiVvF5ilYSYoiiYiDnMCz+/Wn86eJa
hrxppfOJNj0EO+aOoP4KcakrOU/sTgoTtXlfb4+jw+ZqSDOrUtf06Y0ix/AsbeuZwMOCydUl0IqA
IoX+lpEk+BXo42c4y0BKQ+QZ1NxfSLgDdqqkXq+1n5c+hQnEEwuTq8e1lwOEyYMrvHS6Vp0lzNBQ
8xt71xHUjIVW2kkQXt7WATk0JoWUPo5D6lrytljZdE/YAUbDUCIE8L6NV0CdEr1uEmZbosBJ4GQZ
UGMzqf1mdgpSThmqWbMlcwOiNyVUZDm0FWfQwoAQXg8PHTO73Srte4Ka0GG57Mw2jhDkzdPK0AV/
VvnC2go1wWUjHfsdc81uBl0xVVVcnlJE8oGU3Vw6sY4XSResWb5buutO7uDtyFv5RZNPq10RsVji
i5NQNFaSM4Xb+tQ0trY3364f7yki1NR9yUgcCrjuRXE5pBllK8TDbudpq70gt79fMI3VJSPU5y36
WXa5e11maUnR6aJZOcytzBVoP/V/g+ACYTrIOQnicXi8eRDaZA8Uie3Cm6UgYkJELDflbYJH8TtZ
0sHv2ONo9N9iNJfwzrUniX28mD8WptnimeDnEcGHvtV3JVHZokb4ZOmu21CgfNlYHjuEpA1c8jcb
Xjbp63zEB8C3v/di3S0kgXwy1WkC5LFg+m2QOKOazsa4sNC3XmxdflHItJmW7vdKUPI7g2ozRT7p
ZFYmGKw1bV2hJLfnUjI+jAgoMagMlllkUtvE7xawMQXOzZTMQPXuuS4YqmYDz9nM4j2gYR0D3ADd
gSrxSSRnoO04jCPG5NZiVrhKZN8jXmTdaxybQrBzY+IOszti2FvpSB4CVybpDpEkxNC4xTkjXJ14
ZhJU4uKv5QHXNOh6IUvw9iSrdboOHKh0q2ORyYtn9spjsePQZgcvdZrL6BPSCRfxj9TKp2ThDukm
ZZCjUyVziH188GTtOSqrc70dog8Emd+oR+tMlKZOydCfOoL/dY0NdvX98DQzOS0PMxvIh2Q7Xn6e
i+UUgyBj0Sk4r1rpBBjGByE92Nj2ZwHKihMhMEHnKoR8HKDiPOTedBgz041EPBDE4hed7XjBQFhW
JzRBqKCOdMls5GVknjCrxrr9KPTvkdV0YfA45IK5h4TH44rB1eSNfuQK3O5nkif9nKT0eyXSFvB2
QH7Rnbott4SawXNfLPRaKh7U2gRRwYSpHmWTlTXAAd6YyT2XLdCROsXEnkLf2ApPfqgNTgQyOmLE
JnvI9Ei6DJNcWUqf/pk6oIiyayqmoicLYjJrVkRNCMtVfk/lcYbPHL6kl/8GtU+sv3dT/sevHurd
nvsrdkR6QnjwZik4QuKWtUkMROiCZa416UkYky1JQHL+kSCB9WAW4YfVd48CwQeT/xitLMozfcAj
QlefqF8dsSt+8yAbc2h/rGEKDpya1dcxSW70BwYNg8XnnUI1HOBMkKnEUU2osuJG09Y8uDHQ5MME
YGLALz/ontVvCyFY1iXd4TNtH0OpKFD4D33+SvdRtKMViO8OOK9bwjF4pbXMpes7jxqY9XJDqMP5
FELOUTvLylqoFcxnXOSpixi/M5Zrg9h1N12UoohYC6BMytIL1Xk3jhcHsWk+aYablzpOdOEwwYuX
Psld0N7YvUzDOuqkxJ+shLVqSGE9b+8gJaSUJjQ2NktoF2a9MDzXNjiNmC1PVDGLdY1VQvVwLveH
MR0c619mkQTGmFJy8Ow3k4AnMWPE8Iz+1fqKJBrU0RzdBRAZJSoDxCMdcgPXwbi/ANwtOJtetBZt
GBxOUHgR9QzZiv/WkL1IFlYt+AzzKAqCLx5jFr/7Tc1viSv1GWvuXp8Cki1Nt5TQdJpU/ofYiVBd
bRTejY8ksDWDnZ4xjUUasCXC1lcd3PYMdxAGt9P1M95aS/yO6/Y2RzVbKPJIdcxveDJBb8m0BJZX
82HXavmtK5l56AEFZjR8TYJKMFjsgwLR8ZYRE8vnAJrZ6JBFJxUEgsi4lj0hCnebdy1/9XMxe02R
N7I7afyaTJgOzh9G72TsZvQDHmmoIhDI1soF96zsiWW/G/Ck3znm4BBUWOWQzQhgpizA0YzZaiFu
vVTzqpeIScJErYQOtCCj0h8LgoD2dL3gcbd5H2VxBrXatGfwCOKv2ZjGh7qSQwUeY/OVQKtRZKj6
wdP5RNINPM/jb8zWPXiATSCS4T75XhUTXyzgPajJstAYlC5eGjhGiPSjmVY8LpEv5bV+fiZlkEUH
SqjfpAcBsJpHUt7pYlQliNHgshZoHxy3vSceGoFvIKbHVSwTQ0h61sE6CT6rCZK2PBgbWGfkhdFX
3CW9Q4adR6XIooGAnHGNcuW5gOe9BHAhli3FUwMP4aSnWKeGnxnExJFCdXsvIEcroCHvwxLKH9Wj
lW8sIi86l3rj50443jPIUmgDHO95R6hCkpaZAacNu5QFxxkDbJqX4iJbf5fansH3zh93oZ+oRbke
25CaZ2Nbj5b5RlWn4vKiBhi9usXCGU34LCEFjEkwzaCfrydEyXHSM2P4fxY2UywycT2q1hz+Fvl4
jA2djjsVa84ojie6lCdt0b926Uu9NAGBZODVX5yHyufXwsBRmeZHNfioqjme4sjYGwv8wrq4QSok
53qa94c7CU1mcP+a7vpFC6Re7GSPN3COeYF2D/pv7mLVZzkcuCAQs5IXBvbtrqBgZcc/DiRwyfxJ
ZxsJkTzFC/leSGyVeXt7WIjtGLB9EWS8tLshwTKwNysFhTa4Yqv57zn1LDM18JxM0CosEVfQ09ZI
3kHeTFPuvsjJivG8KpSiP1NfGYAousVQ8r8vuoc6XE0m0d1i/CR/mKERAu4Xe+mxaEKbCAZcyHKW
/b3IDxOSnPjeFbQWF5+Gks3sLVnUljzSnnBjnNwW9xdCawkGgNqVJ6lhTRJwQVJj0O66fcJQlX+c
S5b/xY7lVXzQbXkUGqINCrofEm6f+PBhVrRf3zsND5O5YcFw+k7MrtExzE+MlVMnaLlYPG/FPZgu
mV6lSyLBz/oPIg4Iw/f41ZF3PRdVZlCc3HwyPiLJ7mh0U1oHlenXpviVLuc/bBPaNkblf5QQJgGi
1W18MFjMW47zp77w19WKx9LbYQAe+ggWIqSFlen4ZmRb72qFXzSH18uMIJZMagObHCxVbarsGNkL
bnLg3ShnC5Fb/LzjwPBobH6vs9ogIlZiSzHPtSIoozuTzy3SiidwXpqcP+L6Hxai0fhQY5vUrXrH
Scu+oK4RGtN6PLq+OEOACkKQfhrLKtoCud62/gJ8yQudnghs8Q5Yaf+na7O4wr1ZIdq232+H/x0L
9HMetghsnv+iypuPBFVAcbskhDBlrSPh16T0Ue3wFPMxQYbL6THF20u58qnZE08D0cIAnIiN3xW6
pnBUszzTrUVxAAmaJlcSfptF7LWkS29gAlor+p9zSxWCLgMdA7aBuzThBkF7WUhwlLfDvRaEKj+e
IkqAwnUrMT3KxHeAa28lmKQS3U8+g0C65FvOkEfPmC821JsmqJswzKnmVpL0YMzJrk58+CsQ66CD
yrnaXQOk0x6IQKd9Of/kkUOxhOY3bN2rb8iqRBeouhpjdWJqtg+Sj4y+8cBkqYyecrWaxq8wXKQE
oTyBmzUAGezAVrg/SiaKKYyMASW150ZDqWYu/9eptMbGvct7CwCWs6OfxZA0EhianhAJA7SePT7K
7ip8otk2g9sT+ykWtiv5/SCb8agugfO4Z/RfjgXV2pL9/6oV8mzQPDZ+p+Si79ji4f/5MgzMrfci
HkqPwrKxaoadwwpmZ/vrj328Xe0t+YfIJqidF/6HPvfA+AJY8/gvPniOh3vg19TYKsyrlI0rMqS7
H/bn1PG1deBEaL2nt/b3mc/8YQZLmXtkFyB/p1zdcNPl7EXfciNfLyNJbrPSKj7hIE1RKGVzgIPx
KezA8Lccl4gsUKAl0u4IdjrTt1uxAjgNmnTUA0Rv2B6A5ve8VjDDaKx2I+z3FmpX84beWQFecg0D
5Fiahd5wZSY9Ax6u66gXoczkj+yCCOlE6he3txQvNltPJkvW3YRWqy/Hwt7EijAIwHLruUWiUWql
BMcTr5KkZxh/cS2OA+5OMU/rwi217ZHlxyLl7CbAS47uioVV5aqMYJe0lEpeSqpFo6Vn9bygTDuo
vG59ioOKo/NzVKoFkdClh+XCHpwkGp4S735Bz4FGOhItcGwZhSRu+15sUjHQL4P/hkqKewAkGKPw
+QxBbhFvKXqak1uoENt30LLeMagjrSkjNVb0y+2QLWSbw7JR8drvkU082clXEYIdNMJ1BiBp+e5r
xzCBx8i8XuKRZh9/9ZaBm5v5lW57Ag83tCTIaPl7zcXG4FDS0arZTVLbhNnfrv6tEs1vGLSdF7z/
Xr72+gu22avKQc3ZxMtxQYt/z/qOEqGqAm3OcOnQqbaRo/5nm13crtJrEEx9DBMIJyGK59W9hJue
hJ2btnVXRLzHuNsA3p6iyopZO4ogl3mu5UjNgRIYT2Jwcuks7iS4hAU4OfaLo2VZytVgC1T++/GU
wzeghmzL18CpGbySp8VNeotyXdP4uvUlfyJo1gyOUCExsiN1llMXGLguOtrHc0AjIVQP3oUFyiUY
G+kjhwhnUSf4xLSxrr/+CIWPBOPtkMo8Qv2v/hXYo5ItI9G+AACF7YBNyXYjyStrQGoWKBHa8hbN
0FvLDxq6uVydSyN/PHYeAkr5Lo95InERAzPVypRobq/IgcipruFTiZqkFzcr0zuXraGb/Szy6lbc
cP25hKsUK5cS0vnH6tPrfxP0/bm8OlJzmWbaHFA78SxWk9trMIfufoqEiuu6zZTcGxXraPYkPm5y
h9T37xTIdovk5ZH7JqTr5+gK1oSrtRCr57FxtmjqMqcbzp5okBmzsDnCaVt8RDw/srea2xgLNn4b
HSNCMQWIIs1s6zLjIbJNBrA6eJazc1ww2BrfO9L/WRfjR9TtwdFtaOGdViQCTcMrqVHSldGOKvJ6
TQxCWtdzl9B4W6MgR0BFVCSRbUNniGCSytYAeGxclSc1Yum4nw5UM7NQzEGyFLefHnGdz0TC6XrR
Pqk+ReFKAo+CdjP/C3IDb76hIMO3DQuf7HPo9JnXxLwWP6wlpyT0WMKNKCQPJCkeXy8EP7yYpysU
pukknpmC43gASczx7OY0KOhPIXRoXIYfBkbSoSgvw30uBVAiXF093vM0hfHxnUTKRImsYPkiauTU
cBTLvfRPakoBWX4BMGS3EfvWU4Jj26PkbSzAGXKzIXHgQSqovUpnWByXPfI+UlcQUmzPyFWEohK3
wv2ZUT9kmr8bj+8RvdVGY1d04xHSe2A9+c4lx/CyeIxdmZYkSrGeXsM1Pl6rL/XDyN8ad2cavC3x
3k7Amr6RtFmX5FsIz/W/jNhT5kHsRDOCSI+TNlHejpMYN0zrvjcEko9H1uNARImw7hiVNr2RnW7i
G/MUohvlnmYEVQxNJFo4rgkx8usOM+fdFYJ2uZ0Wgh6teqBod/B8D/Znaek/5EAvq/jtfHQRdc48
eeANPPKhwQAG/iNS14YOsxFP5tfOuQtantPPtMzVJUXW2aOfXZzbMbu/Rzud+8ItvAQ3K/rJbrb5
uH1X4OE0Bc7OwxIKbkcgkHBkw29HxYqHT7bm+RwRjkLattYDQBRXRHBZfsnXlwUlDDzPh+JobTvI
IAjgPwnyTcul1LAxqZomnaIDMjlc3rxhkS+5Ny+vadd3yKsqlJ9clg1YfZkxy2LrWX8zFNasbNpx
L49FLU6snv8rU30NkNqPJ7SjHlVf/bcqsbeMtt+ksKW87Qf+2jQ9MnuvFELDmlD6lGA0NndBujEY
s6VLpdT214xIs/tGkW6N1YlvqJwKCcyvGd9tz7rJv40Gcwr9lsT95VYDOFjcTaUs65EvkwU/SkRe
MiZy/1++s2u3B+rntUNek93Xqmw1mQVgC7s9/FHXHooS2kohFzLrJGN5XLFg/hUmplOF0zrIxLmX
8CheMXtrOXWYEBwNTvu7CRrVin2N+CDBZCb9s7tmqag2chjCUqrOkVzJKeoH5puIcLOd9mVEQ+Jg
wnl8Etdv3rMFFB0ZZVVx7mGo9US/bg5vCVHL1Y2j5Qt9WCjViPJgm5Pxw6rhWHWhqqo+5s79x3/N
LN8uXIpv+lhn1yX6/Q1ayAA46OrVg7kou1ORFQT5too5fYqzxS+YuZ+y9zAjWktf/1xWyHh8Ngfs
xo87bVUh2JoUFO2SMDcnd6YqwjkoTL1qjPviqzhTxnUKA86xoqXGPZwX5l+HqEgWBmaq7lYmA83R
WrrV1t+PbrGuhozpcRmp2xqpMrcjDtHRjwJu1dpYAkbdNjlyBZvlaWRu0W96bB87cEaDlyWv6FVZ
fZOTCUxzjAFsBHMtkIPsjN5I8o7Nm6P+YypGRADhHLxwA+PZ6b9u7SN7jtgjIScya7VXfOaldCUW
g6hXAXLIYCfwjot7BmWiCPybFHId60PRWZYX7pf0crmEw5WK7xphPJCs6Q/FwPzKlPyxfpsj5meS
UnwzGmPcW/0YuixPrqa614x91HLXyvBeDmwb565r6JT0+19GmBrZCMfKKDb9zw0DqdIxypxQOyVf
7BG+hw2BiJJ3cN2lF9nFO3LoejEaFgptXREycF8z/DybHzdCkTqUFQtUzlnph9Nb2Xf8B/m0JgwB
ox7EBQr5jiie3bRSo4fq07v3uWrf/JiPx1jBi2P7NAkdkLuywBsebumjREQY3Dn1nPHp7QGixvaU
4qnc0rxC5bXTonFmOgaxABqbvEnCECcffihgnkyompbjojz3BANawVt2gKIJDGbA6PcuX84GTtev
nck1BxkNRznAM/B5p+vdPIh8z5kQ/Md7FfcR+wxXe6bZIlJE8xlV7tCQJJeQcKjGvhUxdYkL/kNG
/3gsrpLR5ovxevJTQWKlOuLu2BoJaMk/HABbfWmCEoIlRhRg25TUnVFg5+szHsdXckt05rxKJWcV
odyU6iPGgbrkJKzUFtVnMj2Mb+szhG87QDvVZJP3FxdgJn1Ra7UlyaOpMpmL2v5WvS+BThR9T3FO
w7Ldx6F7AyEi2IABnuAGEMHo/jClnI/PvPS1OVgrm4CIjTk0v+onAZy6D6UtAmXj+DZAYWKofHC7
ezdfs5otVu7QVESpuRjltSVFe+uwcZ71KUEiVTZlcPZylOcNRjnP/UpOyzjsf67bohpZeoNFpt2m
WBbKlwNC+BJt3PV0BkJdcrU5ZXJARDEyzLIoWLJ4fTkX7olmYWZhJS4109wbNh1lcmeBUUtA00sS
DZx37VB2d0qPuAUDxS525g78q0ICFCTYolHY7GCWbvNW893iObTdIaCJqww3xJKWpc+C/pt03fK/
0vw4eBF8vhW5ZAvw77SbV3r2joiNxUfbGBRHp7D86lxYdw70zmhWbQBEQgon60uf3lhJ8bc4neTY
iQgpNDsGBEPVbpyHwsjtfIR7YyTh7M6Sx0OJ74hnOjF+LrshXyjgXSVptNSZkZ41kkkf3MNfmbwv
AOA9nVIe6Q9z59WHTOKca+F2MPPynTIzIHwDy8G6nWG1RuwGs8s92Y4Wc4Meki43HIemWopHxQUT
tNfinDS3zBM57j2EwOBZRW379WtWTGbFqedRYiIIG5tCIO/1RQWIlRxuTAMv9eRvUkAjK2r5BlT4
NncqR2bUi7B5yeNdH3/R8qdn0YQaRWMr+EYlr/bLZmTYBGVBIvMUsq/mz4aWXHIoauUECOBGeZdT
z0uTusmhnPxe182wTwJE2UmoCYlYx/zmTnXnoBaKG8+HjnVwunVafNjuYPjDTbfbOLA6utJj358i
i/AsS70Lx9wCKJssdZzLhwjbAzxJL8BvEeK1Svy8K54z+Nm99Hqfxt/0A4HtRiLx82NHFJvxw/sa
69m+UNVL7NGxiw0JDCTL2DjjAmXy8y+h7acQuOPZh0QBTOt1G1ix72GQG8/TC+yErnHGGpih0Chy
XLbeH3PmP5R+ewC8j+JxXAmzOM+Nft1SDi5PolRzToc8VeZriMHr6Q0uLA8+33VJWqJM7pWf4t60
hFaWICZ4S0nB3SayIqNXKqaom7gVpFX9qDGKcheCKkqYlC+LS2GWOtujDGwJGwjFjGG3Y49uTzxq
oxqUUv8+5i9Aya8LTSZinoYeBoMivbFHUTlCpwQvBJs1ojxv23IUAMVfvzhv/lsc6wCcL8hce0uy
96EfFbzgN1xYwtvdBZMDPtZIVgN9p5pfea/QoeL0wY1RcM5aBF3qQu3QQJBpy/Ldz4rQ4nuTf0Uq
wHTO4seSnVFb/DtB4/L66/mCAywpL7Ifgc1QB/OO9GofNhQicuNP0yMDdBeaEwO/9bhJiN1LQT/m
tqyheBVWrZwI3s1EAihnRqSPTRPsBTrlkOxMRgiLi0FLC36sYfceOAMNYcyn8DC4SeFnOoKF19/O
cOClodeA6WsqNSHinMC3yJgce7ezMp93xdHyU8/gDJqLks2rJH7ImIdHCgZjzSKd4kpR1A5BoeGM
1cPdRD4K1/OQt1Ah390Ch4sgAcPbLkKqHwVBm9s0gxOM+eYJp/y1nepZwGUfm8NFNxlsAENW5P+6
pmqGD4S8kHeQxmnuOrfrcoDWKoTYUEMQsUKxJfOYgOW3W1yeIGazQfp/uF7fw5BF6zqHkkMjkXfe
3ei0enD/0gydScIiFg5Mvqa9DP1xYJ6ez3oToz0g/Ft3DLMITLRt24aJh04RxLh1jnCp4mZf62Si
C99engIPAxYFAN4MPV0MTQ6VN7nwREAi/X08P8fqw1+oNAxLzYU2l72WjQ5P0q/WWgmM3WALJF5j
CuEq2ocKfGpYi77PzGARh+W66ChW7cJ11m+cz349Dru83TpbEpDfaToSHokaNRo4JCXYoBzSgcaO
1Tn4a7QYC8V5tSSNErV/6CGQylMGSYLX3gaRaR0Fe4qyltEyZNvU1qJp8r2ZA1K1LIPh+do4kRUe
LCseg8msAQjMWU9kcfJMMxW2Pc1dYp68KFrsv931NnI8fqdLRp126tFnsmJd7qClXj4PMVJ0mG2x
G8yuIiBKAni0rmNDpAuF0j/0lsZlXeblFwSjbKiErFbsjndu//zlWeGsogts5YUb5oMau4ToIMZS
/ACFDsnkrdTpalPt2iOcHxNT5k5hNMEJPjvvx1gunfay+9F/HgAisdplJLs4N+fyN329gB51c/oy
uLKJ6tlvdwnq6aqIgTpfqWh/YpIXsOAEji3gm1sQEpeB1qqyo5AINeLs90NsPfv80kdq3Yp5hcCE
7Obihso1+u7HJIK8S3eWV/UCcHLaxEXkJybzqbIP7eXpDxywzuFxCmlcyLzhbANSmYO2AfSZZnJt
4z15W6bkDegBJVucg4r3dKPjwG/8m5J2SGto3pgisO0I7dwS3Jl85GklWCw8G1ViHITaHivu452w
qsmOb5IYA1KEsuiOQnIbK81yBZbitFnR4QqT9MEDQzqqQxXvMXk8Lru52OtrlZ07naAPqdgVwhNF
Qh1RNpBAJGpxkObM4JKwv2pyZT3c7PfuiATuczA8YLA3xS7rPrgwDd3zVRQYkquK95RvrsPx/B/7
ww478DE2TYy0sNDDiGY8QdqD+GFeOff+rSKCCNG/JJF/1noj0au5XMa5R8no597tKpMZYLb/jv1b
m/bAYP15cRYZy91QMVBoGWepsItv9bB5wgEG9XusUxKmEuPJHlXrpm4wq3dfDRsDwyndpk39EWKn
kEpBwV6AI8x2LIc1mzBu4lfMsykvU86jXNwTiiCDMPfbXrNJOJeS3QaX/rFda1rhDMehhkozE4JJ
QIjGDeSM4FjZ4XzUDlxKOREfZLsCumocRkjSQR3QfOP3sqMw/xSP3tIMu0tBNPPcraTvipoNUM3K
TwWB0Fu7Jw2gEOIQZzIcGSz9izZuIbynb/tY+Nh9CyBGQ6HvvxKdQ8IHTnY9cqhOqJDFgm0zIJzy
0+ehx00OaclZhho24AlsAnSWi78rK0WRFj2/ZYl3IdyQsZNsid4NcTtG2yTbJW3y26UKwrY0CvKe
C97ba32sYdXv0cTOENvJyRk46ypbwGrWiB7n/mq+hVCcIpOFYbWRRpAVijwj/ncHtMdMXl4cvb7z
re16FZq2ELzfGD3+y37U1E1ygKAUjGaE1B7aQjnWKZHdBQjht3groZLUEGRAtWRUMECVuFC4pZzV
So/2mE2C3YNR9MDi5YsBW0ZtR0YEtM9bdrPA4ZNfhpGl9Ez/UJkBROpkk9wgr8h+Hy080lODZ2iG
rBC7XrH1fabnOjQzpuYvgF2ne0GAKCaXpSYj87ncZiXiOmmgRVRijfMSbV9fp3aCZDD20f1RJvtd
zna+UAbEfjIEZ75o2wyaFT4+MPwamt5cWnvFfMRKXtbgv8Vvx7H2mLh1xKzayBWRTEr5Zfrmd1UI
9PM1AV8o8bLeHPugbt15B/4xpZRjmQiND0Sf7S7xCNaz9CJhrH3SbU8wcHeafTDe9glbKYkZDNqU
OItOi9Y6DDaG4KN9vW5jMvSQG0f4afkri1YL+ktdNuKkty6JqfM3jVmw5+QOEsRQrb2nWZvLh84U
bPv/5opvQH3cENLSEjeWERiKBtkFl/56I6swt3GG8SSs7eEAvc0WXjJYZGz8S4ApraI6la/X6SmT
YYnWKJG0mWiTq2rwfD1yYOJho50TIGb1Q763ASAyHHjWwKEwmJLDCkbyP5d7Cx0VDBLuAYehHCCx
pSiWMm28Vk7gITC4nn2ggk5g8bsOZ9CbA7Ce2rJb4/ZfZhpkrrG7T0+SEcY6WDTCTtVpKbY/4wsi
prYlsDmtaKaLPJpT3L28wuBk8/UNci2dYbIQ9E32wJmaCb/ndxpwdlZyoRhkFNCiJd6TfAsYhwax
MJUteptwf5x8y3QOwZGK0vCA/VBqR/6b8jy3QdyO/aZBQ0fO0OULr/D/ksbsJj0mvOyMtnJ/9+X2
TO+Lv1j9WU+TBcJ2fv0wcIViGgsBGXTNRBXlTGHIwSSNBD+ItOAihTUabmn4YPMDWTqmXAh6mdBc
P+B393hi/LeZJzJip/+zAB5YUSmdPR20xLj3KPIwaNqU9fiS/X9dtAAoxsA1Qz7G6eTvTHS/fwUN
bJ9MwIigoSPjpj4JNDSxOQt80DBrk2PRbQTGIZsK01Wt0N/4ZuBZjgR3rKTtR7dCA3j0FnfQKOLJ
qtaHwFBZGO8UHnDUdGKzaJHnu3UqMyUuK8zgAeLf3lOlH6IgomQ564nyNPi/FsnEK91pIOmF1IEA
xboXKN1BnroVv7OSdK1lQNSfyzh6KbWS/LqH1CRFo+vkNuPbt3TkbEX6qIMOBweiUU0RdIMqLJP8
XRtkXTLcekF9x4ljrZ60mv6VQZTPqY8crqMNp1SKzv6v+5ONkacv6zvxr9jDBUDMTV5pvedB1ET6
XGMrp5vCYO31/mmnUspM+/k84HWqZRpw30B0w+/dyhq8vlMlN/b5WAcePG/2DMUWlbms/R+4UxIQ
hXrAx7yPnVIKLNiogM+a/ETldPJl+Ufjhlv9sbMhk+ILOyzVlzknbgnWx/ttrh/vMLMtGf0/L7Bt
sHpdxTMes+t/tvtWsRDflWzToZEgvYPUgqtB4GvIzGKBOjufW5+2tCq5ogP26jVeTaNDthgx5PvH
hw+4g7HDe2BVG+ZXSdc/4pLsYrngb0IOYmteHYFf6i5pu8RMvh6SDRrKz8yDRs1voe+oGIfOjZpS
k+IrteCQPZIP89A7/C4RHFpXpyyGu1/xukH1BtjAfF8pN1lgowBc0ir4R626cOtWXxcrayuBRyq9
GyEay8YVw2Mfn/thjgnROsyg2m1X89CuoTN5HUxXi1vk8qOxuslaCHlrjLnBEXfExWU7ItU+zMX8
l3US1sBXKSDQjfcq/wtfQrvR0jzUme50LWVuaxnGukKXvA/hX+VuD/mRg7iM+ankO6NPTQSV41uR
120eBhlboVl0p8AuG3/0TbTDI1w0HZy4W0XepDvRjQT2vY44NMtryLlOqyMc7u9VXYHc8McfAAsD
c6NXjflEzEgNE5sQobn8B1jbRPvc9lKYWjr8lzqkFovp69OyPpods8aPR896bnwPUnbWgLLJZr6K
z8ulLV8cwyR5NNrboEimjAvjYgvaFP0viKYtELXrDVtymplfBpZul42HgE27MEC/7+A6ACxs3w+7
7m8AwWaK9skXQuzjckwujoPckEWRVasVBDwAL/kmjx5l/OSH3WzTlU1S1c4JPx+F2UgNpVE4YWVy
FyQiSDdPRiAPXZ49iMck+PPieo4axI47zD0c16kH0R1pbyX0vk8k/+siZl9vkm8NIQSOIyRr7ndg
MC2ZNUzlL16vGsnJh+aMFCmvbPGYnHQwO+a8KgG9NB2LoMovdnLG+cVhQnMazgb7mWSVa9k01v/u
PhTsnula/tZl7jwjGS9Jq9HcLATkPs7TFH+LDGCU5OwcXpjQkPYgpj1gzZUEFdxcGFBfWqAil3lw
l0wHrJm64xmim9E3ZMGL6sAVGgzlo1kM3iet7TzfGRk1xPU4XmFuopJFMOyQurd0J9zu3dJCDSJ7
AIH1WCqi48p5/fNXid/cgP1fvkjO52h6ZWynaTm4jqKL2XZSMFVldpeBEwRvPDZHAYdujdO/BsPR
WH/ywWgNrKE5TO2Cc2SvMIet5LM+QS1kld/sEXHiouV7TrKLG/Z5N5ejM7a5vC1yNpv67psa4I+M
ddU2Jw6SAXysoK/DcnH4CgHPYLri7Ek/InfV5JbwjTpkPw1a/GHFdq51qmYFutw/9pfMCr60KK21
hLNhP+27/ZbFl8X6GlL1VnkDW/nGsZeT4kL04GYvXBiGVFO0OcftO7dKZox5IiR9+pipKRRF4SUk
On5o1381Hdd4XOgE7VeyH0FOx5m9kXu08ZvixSZNgUbG3+fX4Hef/5dmOllO34JkLMIPL4b42m4v
Hfi0b19xCBuv16rbs3ee3v7YvdILg/DqL/zYimxYabyDNrUEn1r0fDuOzAT6jwPKZDsS9kBrD9UQ
MCyvDwUIyFr7L9M24gLPiq3zFMlvM4gkixM2r1bKCLbg7//Iq24Gw7NT/3msaAmy/pJ4oDSab3hV
czYoc1GoL8VbULNQG25FqKsLfr+BkzUT+CfbTvZc3zBp1zFJpw4gKpodEwNy2SBCtXXU73576Dwb
xYG9VSUIGwKQml7/0ftlBq1CKbBK361Zwqyt+3JZZ2Nxvz0BkVO6+WCJNBeVWgrfzv0T2PG6Yh0V
Orm1o4veD4pc3DIIz9+joiGA1bA9IpHyKTCdQhC9r2EczfYFJ4bk+Ic/QuBt12/reE0HVeCLgHTY
pLQ9EKTcngxinqxAEiTjSR4BQbkBHuYkqWYFvLtSxvkRrEMqMcgk1xuybG6orgo+8IPSzfbsIug1
z2usdZI3dnC/962DYGz5Z32CUU2GZ7SLgHvvyLp0dlTVKPZgAkuvTQeJPOrws4+UwCweyVnHdJDq
vJL+HVdpRErZN2Fqx9k5ByYiIBy7pZMZYSoE7FzUtcRbSMoM+sXuLNLrIZbcxMsKz/K2ghnLVsal
WG2o7CkCZVm2B/fvOvKULDNXB56OKcvzn5YEHqf39qwHvWxM8nQnz6886KFIrZVHG32O36SHocjN
U6VaYW6V9n24hi8A1xw7Ugtgx2RQ71e2rGAQ5+B6i2CYwOVcvZLPutUBNCdQvj8wVp3mQ9DLLOlN
L9XSdfZ2bJByJK9gMvtTNFO/KUWrg95jdZb1Uz4p+AIq2DH8GGcO/oP0GJDXfboUwP2Kfvz/OXpp
DhvX8JvvaO77oCKpAWcl95hDm6pZ2UC+3cLV6rGD2vvXAaqtHoOoQ11Hz+MyOCe0pAEHaHSayeKI
BJqpHPaOT41Q585Nu7cfC6s5VfIvTonXAP3oA6nQ2oTfcH7AUIG/inqc1M0vCiojXUP/7N8PKXPq
VMY9cLHCM1oQqTI1t+hhnvn0GEYeu+bNUs1sYuLaZVky/pMGn5beCtcW72GNPweKEOWM8BHgpFnE
pXkzlvHxZa9r9o92O/ecLJ4dhe4FAA9xTifq3Gk63Z7Td2LySbG1EbazFRfAx1J6M7lQgwPP2+4X
cR4JMft50zvm2O8h6YFTVU8rw0fLCR7aHDAmed49qdQ4xTIUPw93hrE1SQh6xQlK+z6x8QoO6vBT
WVQqK2gKByxQl5h9hOiWDHt5Qb3dcpnuuHuGyAew+cbvkvtz3VNq3IU5KGJweunKidhcYCRb0NJF
sx3A67XmEdT0KUlMqnJ1+QIvcbqLi/uku93jfprRttwRS0W8fztpX4IrnkE/g2zjpf+dTx7tRAjk
PvB0kPZWKRr+JaxvNwnwWs/Z5fx7b/P0Bl/kwVvQ8lIGTWJXiWmxb/suxp3j3jRrhZuIWpqf5MHS
3rNtHGZd7JykC6VbBF3XVLWqXQD2c7dh+irILXe5X/02YxAzwhYkhi16gN1m+opM3+UyBSlnnvS9
QAECLoQKKvxLPRJiZT0JLnM6wolgAFn4R/31v/PuWdhVAEczE7OS/DnzEOXqW28/yI+kBf9Iz/2/
3Wj9PiQhJJkjzYhnWQLZw8o7/HG7GJEhtGwe/9e+ZUf/8fHMBb9CKahIOARLV1OxE7jfabnLbss6
3OA5E5bLcWtsFSodu8VvPTwDDV0GPNrFBytTNkV0dS5K2cLYMfQd97YJzgsN72JkXP/N5r9p6m6s
4ujlf//9vuNavQxXytj74xMx3TkrFIcUX21Q2GTiclpFhpiSgVfIaLV3XSP3FEN8j8o4QNxwPaGR
FJYZZebjpP+kuNs1ShL80IyOIp8U5d0CaP5NAfrlrIgg+PvDizGIz9DGtd+5sngFYArm7aP5lgzS
ma/55wVAbFZBnvgzbw/XvpoifNE5qtdFl2bBF9wXfBdELMkGTNS2QEefO4+GtbZBslahnIyePwpB
FIqwvIK3U4R1omZzCEr8bxhV7T62/C0sSSwCY41IYilCudXcQTHGADA7lJ28nzpNI87PKqFVTK1p
+BHTX3IUToecDsPI/tcNI00K4zSdeIbvm4k8+4vmJ+qMps8RS+H9EzlbLz6kAX+ey3r0tFEtqKEh
jFQyP6rrTTtCDY7ufb03wiZjq4c2ZaXxOtzDoYiAo7+5yVE23RFcmKqqUTwQdTG1UgsuKtCwigK9
d/n0TP//IiYL1pHznDfXy7xw79q4mNDxYHv7wQPKAsgirg/sXwWNJ5VJKSf7QieZF3rE27xj7XAx
p38UE5KUxqS0sherPJhL2KJqk11eYATIU/GZwIZUv5iR4O0Etji1dBu6Xz3O8o43mm6swNcXUGGD
+4jpZDfn6ZiJadXsQ7qWaLnwma6ZZvDWRg00jradCeZ/UKnoLRTaBHJ4whbUOG2eSOQpiWxIU/EY
v9iJs6roCVCR74JL2sALKEfeJQP5o+yfRzCbnl6yYtg8otTWJvUjCVTnyA++tpHkJH168o47FwBL
x42jJEzT+B8I5Zrk5vSYr/fpWHDOMRiA1c/nHAoTs0QwON7k+tGY9nObMqj/1GsefS8uoDOXQOPe
nYQGapBQi/zfVs1cUBSM7hTbpESXmHsV6Kj/7VVEwmryQcRtWqY/iiE9JhrSHlCzqWBWxT+l4tBs
9OLkSH3vQWHmzHUuBeocN23Z1BC9f6j+8a72ZLxLKRofDfZ488EQKL0hUE+n+phyuAVcgebvLsd0
gSH9ruKHWoQAA3B1XG2xVvg6Je6mAVLWyPWe5efK+VGezDMLEhPIgOT1iwttoXimIzCF5mPEsSMI
APVGMSb2KDv0tzj9AWlVfIVPy4NK/NhCCW7gNemsbXtr3KBdGe268ld15Ca83WdfFnRxNzNPjUW9
Os8lWVQSe92em0xI+g2jfWtyiQy2eMemiAlNbmVahcegak79306wa2812Z3su+UsfyUTQjJTQ/2K
SWf8yw6rIQHwCCajESTDHeBcJynPIlbDoGydbPfgMhvb0tiwDLWT5iKtPZACVgCqzOSIrVHVTRUW
SidDtWCM9Fr/ztkjr3w0dKwUeRZJPVH1RxGodvOvlLbeYMRBLdjDI4YcfrXejdbu/CTnM3pKpSH4
MhlpqxYKh5qwpnztc1lVfGhnjgEzu7SsqoGOC56j79KDoa8WcG8TNRC5PF2nhlf2QkA93PyZ2XSP
QK4/DssVyFrv0zFC+7e9XydwTUWQv6SkFmzeDfuRqImlhMFKeDniKtTO/zGYDptTTq++Qg3x2oCL
JK1wN2mqumA3ZUaHGsvoQtGrZ03Lixt3KQMVuiQlXiwheKV4lap+wLOiD2jtKpzNuzlwrIFewDIr
Cg4emBznD6ydBDsJsophobZHv7YrtnvlFsB4CWoPuVx1alKssY64yQZomJkGz2qCE9Cz3K04tkOA
6l1MqSU10InmdLZgNklOTCRhCcEaAk7M59hAQ+8KPr94kpg7bwbnTzPv2u4wS1lzbAZScA6ZteNX
20ec3WEE8AA+udSySR7q1tSMCtGaZbh+ZhsnSkfEAZHAuAhohdFrdY3AjSNn1iT5pGVUQYOyg1OR
VevuKEBWDHEFn9WVrzFktqMYvGOC47oYQz22v0iq9F5o/OJjQ/MbAcjgyS0eLBcRdBOkuB1iPbYQ
1kxPmWCepSBtC08Mq4Dq6Jk8F0ugYREtptFBykk1vdIJ7gxcbPjlRsCYSEsjYSW6kOcp7t+dJNp/
WgRTH78Q2q+OquqYtYurPn/IMrrYsMUtcqJ9tBj3rJaPIH7EhWqjkHbdy3EpaVlTH9wFUuO4KmsS
jjAory3lSggOSGlwxRxRgMSp8j46X6jOLmJykG3gQ+LGmrktIOQ+FvVTUSDpEP8MrIgYurh86ZH9
SUFyCaEtDLOYAytYAaoDemYV9CzPemDoP/MeXipcYtV8LnCJhRVwdAj3ceJMCgFJUc7qorhXsZB8
nEu5a2Hc7aTJFQsVTbcnu4p5KtCerxjWSswfERRrEaVnY8NjxguPBJ1LHtoN8rKlMtGVBjHzI0xm
OAN7/0tI93BzUtDgQbLfQhoUcVmBTIinT2cbJ6GeyrRqpUcaPoBbtZ/oVENS6ptfTDRCudHkL/bY
leU311ND8UVuJ7KT5hkBkw+sG2eq/n0cf6iRjCGQVMeVYtTzM46aUqhOzp+rEV1Qog0XoiEv24QV
gzN+KTaqe0Jh6FfBO7bJalbfZ0rZFkjOj5HACTyiiRKYiU+NJfNd1TTLHJbJIxSl6uQidFgcNFKA
EkWmeh+1MOBwzqezGoRDeldl+7s2In2S7HLfdDiG+oNCYyP4VIgNbh3bPBnE21VtdznjRbIZenon
hfmat23wE12o0ewBI/3gBAfQQrnoFzOSxmbg8nlpToVFnDBZRqVtE4MQpUOdrH/2jWbtog/ZzGp6
FwGbyIqQ0eetvs7uYDodoQC59AkXkgLJqWNwtTzPpBr1MRYEgKTsDG1qD7ganAfqF9YkyIY1yPj5
SrQj88FqtQERoQVJCftXSE/9PNeMyBiZ8X5CNr2vYqFN3I9gmcNpt6+AtgUXvin4ddy5dwUPF9zr
RKJllsu9CajlEU3wpJgvS4FCBuaQPybWrmkXZevz57ZOgSjZZifHMxTx5YBjKmis++PE3sbZmh+d
xmsKnXo2f2kEPCEMQUm44ZzB6KVxrD2uFawVEYiJM5kKhuP5GhRjV1WmiUFG8VrsPb6R2gi3Osx7
EngWqaaown2uJB6N+w68uQGEFN2QBAKFsXlxlpvLQxwGYvZ8T543kiPQyMZ4+cqL/elorBSjdgj6
rn9l17ai+Zn5YEEt76G/yfUT/wjmPZ4L14wpNTWOAC0FppIVhIV1qrjIwLg6pTtKJstlQMPs6zoC
RmAkdkq4aJer6Gr2SjfO5e9bKaYVC9vKZMmZjgbL6Lg+rpWCD3kg8jA7lM9PYafkCqdDGRqVal0V
ZpJUEsNwW6yuve/oVTUuG+5cfSr/Mo/y+vXSBV3OsoW/2+fj3iSt5inhhvkDa0CqwcGf4QLy+k40
LNY/+DLQHeDSxv9iUJVAUiVXar9fkd3WStEkVDCwRsl8CG01n66r8ORG2ivA6utmzpHd7oZzz0Hy
3sP8NlCPwHxS6RYbq5f0zemFKDRqjth7Bg6MSWbEu1CMfc0VYI9jIxAGDM+ofyGc+3xbD6VvKvtP
4E539SireQBU7Rhz7D96tIznp4UzmyauwvvnwAg5JWfe/EN6j4DxBcffYug4yV/yK22NHIbZLLjy
zSvPqDACQz5+zA73xXjuwcbTXH0jWFiO97iW7WdtNyot1nHcYvKPW/lZlJkHzs2/iqWfXLVe/J6H
ChdJDfiMw3FwJOMKqxLMQoRWOB0l2jlLdgEwVTkW+rcufJ7QbE5Ux6vt/bUQLmb4CBZS9wuDTZyu
/lGe3VIUtXJw4hAbBk+NDs/Qm3a7+YxK4hnvC36P8sQIPaHkxoE3m5Nj+sX8i5f8xo8odkamgJJc
uIvUmtx8I55tPLPtxisrX2VtR6rSjdTWxW4tRrid+8xEgSmmrtLaE+UdC1f+4QqGqBkJbHGQVLIB
J6lunCPnY1tuPVc4la3uH7JOqH7kO7XgbITPGXh9DuGtqN3gpV/FO62XzWcTDWlqnA0EXqYVLYLt
voWMf+KAXG8yEnLnyBv8xVGAQygU99IYg01lNJEFa6F8DuznmuQITItfBjC6WIyGlY96T3nY3xaH
9OSPD1TAaPP45MwOwvGhoeXy1VSmrWKyNxm7nMLT8KcKqKUveys7920waSqyhnp29peqRZHD37aL
ZOzhE+lyL4pfJgxCk9yGlM/cf8EnSdP0RnhvOxwSJfcfeBKfbwl5uGXjsrbMfYKiQHCxjL49jk6D
oFa+CsMUX+ZYPFvLi7mloN8tADrqnwQPjgPtb6SSnwf2MCEQ1000ceCc113qmCJQ56Npb00+Fp6h
ZLpzIjTgvNVr5ChiIQCOQN3UYQBqmacLcUysVfdmar1YVdzZwLfXcMOO9trzfZp6MK5TnWGjHCNY
HeQavAs0AZH/IGQLYM11Pc07wQH2LysTFxdzCb0MXO1Up7ygq+RCzrZquCQKgxAuYUymreoSR5LY
giWpABkpjA+gIsg0at0tOcx8iknz5SsBSPdxxUqgMyJhWQdSGuf9/644q6ndHyoPhf6/RW//FDlx
shpOjzVUwkkUR6INl4WEIRLKfE5tAEWI2ztgb/HJVMWpS6WSBI6sd0YIu6YwItR9UrqxDXHRaD7/
jZIkJD7mDyD4bIn8eVG/k1KByJzrpYc3Almd9lw1t7u1y1nZefhNw7qpDRvglmzDbI86Lobue5O+
I3x2qOqPLtEnFbJiYmKKWEvgb98dMXExYM0XG5WXP8wF1h2XAPqXndSc0sQdnNwH4NrSPxsoMnjM
YeOJwKIfD3mos72CYADCNebVLVBR2+9s+jeuo5mGoTN+ySZxmy/N2s8oM2lOyaI5LtGPuhGlEUog
dEZtL2EnmsrihDuX5x4t/KIOy56YvMfXO9RIk1/HuxihpKbOs4qf1mrqRoWTfkAr7tQWPYpGAlJd
VNuosHCpXFUKiPwuQomyEiqFhPuFbxqpkqyZ2bBEXVQpQ4KcKtkUWcSKTlZlmi98sGafrJFDPnag
0L+tDcelSoRF7IMvELColhE59vBl6mKkYJorw6PphR/nyrIy/zIhDrfr88V3IqjjINCGj0opGpDU
z5Xj7xkmoTC23ML/ofB4cUuZg6FHvMB8tzo8vImrRl4bT/uEQHw+dNQooKTbNjXXE0D5I5uvei5x
xeTQuWgvRT6Zi8FrSTASdmUBsquZwzP+1mf18bVHT63znKnGC/tMqkMPwsoAtRGKOfjWh4QoTOVu
zwkzbtVlRAfstRnvAwnimq/KuOr8hHNrUL3XnbKSp+qFrDebgIWAhPkrMx6BcqvWXQuWLFrBHvCj
L7AtakFW7Ggxbjn8uzEeHs6RV2P1QJIb8yfRAlZa9LjMAFpLah2kxJPNIKei55f4DupKZMfOeRnD
oN7YIqIve8mpeHdmawnsrsLIaTjSouigb2nqQinA3GpDJrtm/OPCzeBSYabwjpzyVbti5O+MqdL0
QWgYWb4Z75qpPXOoPDyVeWi3CmBpPfOuLVHNX7R2dEjmC98skVtMEVsOoQYxiTo5IWat0Tz7o8uK
FQumJvk/f5P/BJ9f9axSb6H1lwDaiHwq86Gg++EoThA0mfQTFlQANl4qTiVZbQ2PMoY0a9wkReM7
4cEqxWquOQLLtDhhT08r2+4s6U/K/2K5RsCjjSQcglMYAud3PELje193oReVil15Zl5SYN9tqkQK
3cssRFYH1wXqqMj9qBsl5iZ4fCFapGn2udMA+JZuYosFOX4I3sHnWiN08b9hcrEcy8aZWTpII8ul
FleC8fnzJ2oe9Ws+hISKNjonEjGs7H35VQK0WEAcVZE8UU8tFxKukwLCoDYWwFHpO7l4QTLczgLV
oM84mL4JwJLe0kEtVXTioi/rrj1GCORD/9gKh7j/dPQvPzdmWN4SehULPVdACuyOHWc2zeWHEhAw
e0rj2MfNevItFgM3cUzaacyvW3VRdmMD3nOaq021g+P0bnhcCnQum+4Y7VhqVui4HUBD75SIgqrN
PluZeP7COjmEQcwNCAV4ej8Udlf6nKFtzUo8ohRy1KZEGHXNFm1yXGLhM/TbLR/a/uM7lMLnuY6G
bmE045Sq/Igkvi1XdyVVWaY5+RHkWJtCPZUvjXU6P4tCUYGLxDrFnY2KxJLR/Z07WUzj+AA5kdJY
Df09SfjDLCnEgxJBFGPw4WBibFn7G63/EWC4Lz+s7WE6BTD1bgOB08pr2+j3cafdGECnrgLEYRcM
NHOvd8Jl3G6m0fmCXXXvQz6gVZvd7Ahu/R6+i52q1tnyRM5FOsiuKgDTh7HZWJwl1aLD706VSCue
9CA2U3ReKGmyQ+uon744sGv1RdJy3nijJgr4zYsuVYsg7PIPrZAJBG8dsxZ/YsjfCDDXHh3hXtKN
CYeCnGICkFYiOSPftIaaFO9eNRHQ63Oe2F0JnDDy2Ru3K0zzZnYIW5zIxCL/KEAY+XljE78qFz5Z
X8xPKq7CiUYJoyVwCXVCE4znoBxj9J2neuD19rONQ+AYKbw/GkOEm6vDvpLr0K6kFw6OX0d5mfOc
NWfmLVYQUzyat6eDyJsntz0AxCeb92IG60FtanGhc8q1aNH9W95TllzvaHCrZ02Bvv6nEOzToBjW
NsbdikCKCh8gBE3HolO8ZB2uL5jKSYNuYf9jIpaug40Kewun3Umr47ZNQlVo3EN/aWyUbUAnqnYj
+uusNhIaGdPaegyTwAv9Z1D+gnVarvyOPM8437b7oz2VrKtssXD0M5SF41G5YIPkBrUj1SN71DPt
VLhUJSv7F8DsjZzUAZRM09YDb0E58IQ4s6M9O+PCYFb5tQw6iEvC17dcwfMWxJ7nGgcDNHols/81
X9IcsFPyJ3g3NFCQbXGKnZdTik+THtGuKrc36jV68E65tRi+ntSYcWidAr46T3lGi53gnhmMji15
MeJHnDnPgKbt37oqredTGJgb69IxFA26lR7YQkwy+GEi3Ar2sN3MAOuf+T5mr6dEvo6wcTLiOa/O
scwq2xL2x7RCY/1aERNUT6K+a1BG9mHvUf4Oj/+CKFNqDSbEBYU1DN/4wlDN7rOYAX7vKhO+M6Rb
RdpwN3ho/6GrBXHEehD7UJ0VZc/p7y90BKSDS2zFPtqIstZgqrxjQfLiqKPMSa2LRMCqpiOV2WS9
Ew8LkxpYkOn4FKc4SZ1/Bavt4R0tNQ5UhTcQiZgVoSWh3QrNRBfnhLnL1Fih5/h/+36MHJL5uN+u
ZBODfYVBmdg7dBOOlQP0DTfzxR42CIWvx+d1MFqMhmSK7fSrULW4bvEzDBICk3bfwrOA/1A8l2vI
hXZF8auipUOM5wAe5+YGxpGo0R3myQ3OyMR4++aUCVwja9Hba5Vwv0NcnzSFx1v6zw1QTVW/3Ll+
CJEBf912AnEyvRaRm7LuWRiFMfAzhRxeBTnayneDCbQM04bGDZ1KS17HZghbMOx9TBU4wzneDdkh
3rf56Ram2NS/sV/iuumXj1k4nyf6IKZCp2o+U0T+Mw4jxCbo8XiHn7ldWqEACqbbAMTHqHGMiY7Z
kFwGCTtG5ExPe5A8P0KfOjpWEdKppZ9qHVKshrz0S87/t6xORZFsGqS0ZkUFCzEGVvkqDs1Kuox3
4gZ6cBeKcU3TmBRi4RCh+YoRIp9A+GFuxnuc6bvxqp3/uv4+6F/DUF8GsdrlKuO46JniCZRlQjPQ
MXlxABDW7Ks72Fqbr7QowKDjbhXKBX3avoUa++ilGWcJdecezLbb9x4COxIaE+jKH0ImxcKlAFI0
mNmEV/GlVjvWxILtcmKjo2O1Pgzip3xKpPCPdCP+4r9g4R4Z+cE9o2oqfrUrl9RSzBrGc704rs+H
NFdYM/IWLmBpng/iVAVGyoZs+B3Yjd0CB/7oBn8El3lrx9dfZ/jlDE3RznwLriFpqXs/DlVs470L
w5yO5eKMdiBdYw9g3urQL4+2MVICpk9c6Fi9/2CK8SmdC4zuiP0WXV5iXCX8ArSHOtNrBCIfB29I
SYLnxcm+qIDymNDqP4lZyDjKJKNGVAWSSsXS+Th6/cI5xb5DFxsLso9lghzcqeJZ8K/QqHs/VqD8
Xt9Bkx5bNXhspJXYDTu0mejZw4zOp9lXY1JwgNw7USZ6j8s4IR2cB2CpsFlxPg6jb5yd68cEVjmZ
U/nH6ZD0jj4pkTC2ysC4gBgyzKbu/wmTgtMnapS/NG12nsmCz7t4HyV7I/Vr7WP0LB5TeY2QW4Ha
6I5CZNqsk8Fh144tAvbIy6IQJJGzAR7JhMjPMWadUz0TFWOop1MR10f8sa9mxYOHdUluddOd+byF
w9kFagSrG5oelNSD31TYhmJp1Zwnj6I0uxaPjRb35y/qqliZBRJee7Rxa63PrQTgmP5uuNeFd1qI
M6uBYodoKobgUvJ6o5FhgDa9wREfYfnlSjDcbzkIfqTYpecM7rtX/Orq2j9b6u9e/GVjMMWZE5zX
lAzXc/QgsCtKvJmZKWGVOaIiuIRjWZwCZfOvRwI9rsFvLrnSy9NGoqCTjqXJ53hi/xy2ZKdMi7Po
wP+eBQuTjoyk7RuJFZcTJ5txE989A32rZywknd5J2WKcxm4YXfL7OZceaErmLKC1iIyZusklyR/r
HCt3X1t4bp5jey0KKQSsxoiBdB1jBYOgqrEfebFqfLGVYEvL6ICmflEK7tYtnQp/tbNk7nDsUckL
BcJRmR42fImYMnOrktUGkf2DBpTzQlLO3CpY6lD9PrzInTy1/2vVHNzEbXPAjm/CYnlNhn0txhE1
xPL/v7/X+oKRVzlmYDF8134FBR1PoHcmrbXkGoQgHuEtZv/Ac+SnZPEymcOLwnNOBh885UvmbSLC
gKWeAhTimEb7u0iFJ3HDUdF3MXyKdBkeqW+xseEIvr02EydJR0CBs3eCwHgeX3rmOAoaj5yyrh2o
5Zer0CWLoCDQULNx25VNHfFTBLZg6XKOvOGkrAKZZi7Ccy2+adTMXCkGmJleLmftx9eUvIyCMQdZ
7Ndjsg5EsE3PlBT5ID6qG71Rtid7HNpBCSw638z5NbMKEiCCxhtoi9lVd/cThk06KEPiCwqk/ygj
po0jbuP+qiQg5IAj2Tc8rwp1o2riydC9yWNAMIrYU5Q/ofa0YpJ3X+w5qEOr0J4k4pgY2j+x1fHW
frzz7vfVM+Uoi8mQkGil9gC6Ji+6ZLmzbKhKW8bKuI4tOICYDqoGD5UPoEI637FeqvO5RxJ3riez
WvPdwBCOt9j6KOmDM7yz/LKiW9VzeD2GvXKfib7EHQyobY4zxaIsOHI4kSrCCjnqy04TvsegAjDE
VIh1GczplqloBSD+/0MZ/xzNZUBhu6oM5aV5MQX+GC2jUoLTVUtzb0O3d98S655tFAK979E5dod6
hHEYDsoymvOE+VEq4M36ZA58+3ergYNcnzrdb/l87H5dj+AKJ+TND2FnglBYaUzkV/GyOGogedsv
oAvcg0INMZ8jkfcH2djW8fLY/ElXuUjAS2dnGn89a1PDpi0eHNDXy73feQXBfQ7RpCpitx17Ja6K
WNdSDMEJIGJQWa5G6K9EbXAb0MLStUdIT1JHvT3CFmdGbIzQTPw8lqauNa01cHDxhwp7y5oRfHi3
Wfz6envDi/qctX5hz2rN1FbxausCWCDJr7PnEOpUh0/7YKQvUGbv97t5h5fbCMDkPO4R8GAfeBuD
X0UVA2g67lwMd1YshP7HET3nqDVr/QMiZDW5h4Eabm5Uuzae0+DqZmt1k5Vp6KFDMjyWnZpvOznl
Zxb22SQ9S0cOXExknA0aprx6oxzlLlo3PzsVj0wfojSrhKNVFslpDxq1X1R7NPByNwwEFQOGG4FP
5z6aW7g0TJmv9tWepRNcqPzU5b312XdrOSYZy4goSyI4mPzXEOE1Q/dgSoU60G1AQLzxjduZ7HLW
/zC3qSK1pOFSALPj172f9dx8EowDz6cm8w3pBRXsbsC/liQfH4qaRo/N2DNw01PhMnvB0SiDompS
aou+4SFKhfTUgLdMGOdImlamFgVrv8G3b63vTlVnjdXwo5nzWYaBDbiiwxbXTyQbW/icbGzN/2+c
xbXtPaSSy0VjfHM1uswKEo7LkJgpyRdcw1d/QFIgfp3bcdJHkhI1uGgFX83mSJVVrkTSkQ9kHFjQ
vFPFQnPokfpHdRiQnbDVhtC2nVGErKqGG5/zatH2nLYU5dBDEapJBpPRrdFISA36+HUa15ROq2jH
/vmQH8GFyBU/A3Z6SCh5kBHFIl/o5uupG0xGqIHql/KiNxRfgeD43vxC609lTqdAYqecIo/gWkhA
ETGXB6d39jODXNZ4zjz5xUT+VIi1hxR4tOzJ19RbSZHY98HiaAf5Rei+KxMsht9v/6FL56x8OEII
FuzyJukQQNblps3iX6xMqgrPOn0FUJc0+xoNRjCw6fZUn/9lQ6HBW3OoCM/pmNufzLa4suDu6Bp7
/JQcHFVPsQ3NAQrupOuHDawQkjY/Pem4BJ2dPeJJOHGXcebuzpiaC9Ty7Lx8hcOYIxeW60QxdQvn
4bFmpl/JNHmVDMmP/Vb23ttrKliPY4Qgp9VBPU/DaI/6MBhyfwnoGZekIQzymqi0noDeP6cO6Lv/
MN4JflRnf20lzhFy7zNot50LBbpZR4BlMU7rwjlXB/+RJAfLSnQoktDdJIK6qypXyX4Iujia3v5b
6pIB1QOMMERMS0KcHODPnPbUHgIkdXC4f/EMgC46xkjrAiJnBKnaJylOLSlfZwE46bvs7fIHypX1
sF1/6Yl+l9onYVYpNkO2u+kJRy6wpVnykT61MYEvQ5K8AoSp5hM0llgQ/QQItwXr0B0HPbSi0MXM
/7EHeZM3d4K4q36aq+gEKDLGUHFjoNhzHUuqJzHXWFI9M9QGYEiinmmRT+wnJf6PM02q98x4biNL
q3CiialHPi36c3mFfRt/TheOSktNWDHnOdL4NSe/GHdpzp22+jzlgY1N2ObTBR8rXgTjvnmJyvlY
r5SQvJR+6op/VsaCjMcwCTvDk4VqU7gMUYEcULpsQCTf3eYF7EdtBI2j8Icld7KrzQf3I8p7WrFM
0Nv3eGRAwaPuWkKu21YZQ+k8lDNCvuIFAEKWjlaYSAZ+cTj405x2brppgcCT4W619ExwXJ4IhPcl
GR5SbqAsnjqN7MTYqejUuP9Zb04WVDganHIjkN46Rj5QKrqkSjE3D4urVTW1ovj3eibparkz7rCu
MDFlC4EVOPbYs9l0gxKILXtXDIyEUCXdSFDryJcGD1+tUL5ZT7NGdM5hp9X7YCGB8CVfGU+K256C
XDeq1LAoGwwjtgsnwu2TxhrZzOqlhi6yYh4dQktK6jHJpfBRZ1BpT6aafuF+IMpW8n/Znep3PrhG
zSHsYFCtmepB7OawD4vKnZaxYj2GYXTtMORRp042BuTyWxLSbXITXtma5nmylc9ab+sYK+jfTNjM
LMlFcRALrMxvoP+V1Mdy/sz8GKKqffBvo+rfmRTvh0I0mr5deF09VbpOXwfg90dJbRmD2QiPW0Yi
3ScVgiwHuIK4n8ZNsjIm0NurcciwHJOaW9utOQ9zePfSH2qbU6bqt+GTppSuz5uIXS02VjQxogVX
i2sBjvojJu8D/fLjyscufsyGu0FJf5moExHYrRLx9sobS1vpPFJGzlq3gmAjnfvNqL1uvKfVAM7g
Yv/su5VlUtS4N1O41t/KAyyJClIxWEyPjfxjrjLTPuHun1E9D9g+f2IfCKnqoOK0UuNGXUb1UN3d
eitMxMOhB719ExjBLCMbVwcaJRgaeypkPRKaSsVy9Kh2Y26NB0QXid4dHirjquNH6fbNlZLDBTUl
kBvHsxXKun+Nh7TdmhoOiUwYTRzHIk4Os5mf+PGZL/hGI6h9TGKbvvrKHydnuq4E7jyLQz6gYjP9
rIlXbK5NqulOe/oHHB4mknnV2iFqMYxdwGIt6Ae8T3GgPzHEKEPalWwgIPq8Izr9rRjedZKZYrVX
/g9ULD1ZBC+8EEIC8NJrAlmMaS6V4g298+mrrA9UKzZWact5kwT9Vn4q+O00XlRKRgG0Rtj5l+7d
Tkf5f9LYdZkBlZy1pAFIOmp2ofQkJIY3vPllZ7wf40SSTkhoxnvW+zYbeO1+n2/ilOcaM9CLNYIM
2HP/PbReTVflzDysRQZ3NN4kbs37Dc6KYPhTo2BA66IeVvfwiSsaOLkJCnNnJlnGLnQh1oY0bDiZ
osuA8tApGWr8KWVuooVOC6+0Jk7o6iThSraQQ6L0PPsIBD0UllIJSDUPHD7w0iP0iK97pyFdv8WF
L+Eh/tjTx8FQVQbOFxSHgWIGlbEOkz9U3dGGZpZeCcdsxuzKiNtgW0bMXic3n/CJJSchqhYU3tGd
kvtdtlNkJ3+B9elQraPBXM+mmb0M1H/fnspjtaUjQPkm6OEsj0f8OIJNG596KuGA5crj1eFdeY6u
/Q+sCN3xwJusfjwobC9osQYB22RKq/I+NmtN/7wrlvRAcfxgpAOB3ftSOqp+MSnxueTzwhjmwJ5h
9xjscfLx7uQsqg8yb4DkohKMYoDNXZ/W3J6bw3LphxKy+rj73m8xZqiwb+1pk+iwGgSgngdf/pgA
O5unkA94aq916st7ZA4JAy+dYR7yPG9f/9NVB6tAUQvCUN1STyurw42bIRk8euCuxOJNKCOr717i
GmEVGzEuqtwJXwem4mZLX/hMG5DtMn8zujDIhq33uulMPUSg4NiVHkyQQdyhWdTSb1/RfiHVGDLr
x2XX/y6PMpxXJdlK2gmFf30hDf2sfVohZLrHu38vntNHBQelGi4tWdIXl/k/WZSfwKZVboKcVx4b
OWDjGqaKS1NwpCKyDdQTiozrZzF2tt7Qeoom3leF2Q+I6GHxa8LirwTrIbt7AZ2v7vCiYyeDzyxO
SkL0MWJZy1j4ATWREFQW2uc+ArVkdr+CRoOjvf0wxGhWkVDQCB6DQxgO8xhdxTc4T+E9goio7xGD
tbTE5HNeDTu62VPMK+X5TMMakkGCNQ0JQAS+sRpcAsqwdMtClmN0wyZtx+hJnCIhwHaW2qXtLeSW
glMZo3M2kb65BI1rqACe+tnViEAkc7MvMpxOw+W+NeUV0Vgd/DhZd7KvH5fklCBTrloRfVtHRvmQ
MVGzTAyXOgZqADm0Qj95v0FEoROW8U+OkcF8VGrdBmjg/9UnLhK9mAxMuMuKIPnJNRteXthY94kJ
WTPbzYAmlhTedjDOOzeYgoBB0CsiE4GEOiwPhID5of4ciDeE1gkAflcAMXalh3O2wLkIYO7+0Xw5
tGmLUh5UQasMPYoU2ikXV3u/fOzhgM59qODJTheIYW70EVMDGIB/Ng8f+zhl7aciveabX/RE2oHN
4ZZrg+xFSdndxn3pRcM4JlyFwmSJyTHcdoyKPDoC0jJKX8vil1k0y+4+ioBpGlLCLkohHIgnY9Hk
P3OP51SjwVB6CPfPr2yYbgct9L02yt4Iy8MgYdWd/6qf3noMd0d3OhvGi+Iqj0XYOqhmktbQSPI8
OnTzmPOEIN8KuCRc3SzYTvqivZFuveW9RqueLVDAB6take7CuKyNk/wgVRD55eWBCcGMuwLZnT3q
zwXrI/9Z88q+HHhEw5ERM3B1N8HLZkEsJftyc8d9fB4YzgSaYKsBK1MQsmD+Ic9VFpHe6fn/I8KG
4b8H5DRVg83IdAKY19zmHn8ngTSD/kLE2xk+JkOTXMkQYPVZHPAcMXv2QFQTm/6uxf53VP9p/C8V
nlf4YFowtuXkLHdLKxaZQ80Hv7/5u494U1F+qHWdR3gUIEDRY1T4kAWqSFfgmnzIMIWL4tYadu8+
I8Z6uIUWKtaXk2ePU2X/7NlHUEHZD06eocZWJO3Wt6O+KcLueEhzodDha8PLfHMGSh0bFjXUSkBW
Pid4/LwjMiCTbRin2RnwQH8BX2bZsmTOORymzsoqhgLntu+PWwMsCSdOmECLdE371u67RNPKqv2/
okNMJPHLUnys0PIxG5TG6t0AmbOhINLOewV2ZRliovIdYuRVDESXRPbmBbsEWwWpwkEM+KAtubLj
MLx7mWueK25ZojUMKzbfyL5+dbyNlZpVdtqpSHrzb0N6mxUCNkyPSgACzdXYxQu48bPWYXWijdmp
yXPQY2nIWNzBZX+pOIGitdzDl+tSGhCMeBBbvJEbXYwV5H3UtV2qslYP2BKSvQIvQ1ZhL0hdrhMp
xJQUe3cEfuAgguyDLsu3zGx+0uPhxjhTtn7yM3ar2XXWxre2eYZVFe9skhY3mjFlxmgruIltt7qP
s7oYsSpnufls3aWVX5NhB3bFmneD/EIt8zsS8mn/8O+Fyqfc9pJThlSwlqeBy4QxBiElgb7GIsJE
8PlHDPdIwDHRytQdOniv9GHXryL1YQm0qEUX5SRa5XXHmRfFj2J8xOXEsdNprnTcqVyHLJxyUreV
TGV1efrZTuEwl/lqpewL81dIyLk/ZfWC//JXhmzv0SDswJotxaT+3fXcolKIKmSEC9TDqwi0pPZ4
TJWiry+C/aOoiYE3Km9V8PWZWvBHUelt8oK8Jn9w/mHyI7Qrnn8CS0dDvsc0IYy5qSVGBPL/AW2l
ek+1K76vdfjcz1CCkSZLhDHwyGpQilYQoZYUnYi1G4uducACIch49FGxHgn70xBsnuVnQljzYbOP
cbPCTNRi1Zq0DSQ9xdAMUkhcNUkQLjdFQDnM8BAH7P48vqodPzMBWUA1CbQnJRRBFnvONMVMRAXA
nqrjjYKNWzIYHeb6RgBKbisbDT1ihnsUxVNdRE4qnIqWH+lhX+mZyjNu9Di/kIYQob0XJdsv+d01
b7Cp+CYKWZgt35nvDy4ElEyRUnFz/TwoOeBOJdwmr+GyAwX4wS8GYT3eYaNwU3Zr2UQbOIvBcllj
HlcyC4VX6mZnVPQ4Ok/HHnwG2+wurf1dgP5yeaHnCD/9hmdfseupB45qKBVbbPdsl+Ht2OkeeBS3
4m01lr8MkUWI1Vvk3eLtHNZC5fB2K1y333UizHuIIqT3SPrhaiFxKLiCilNH4o9oCCWp+OZ7Xiiy
bIkzonpkktb/5NQa8cUzFjrsTpz6JMcMVSIjI6bteNhwkACQEsbYX1Ky2S7robZNF5xU4CtorcUK
iNvpMsXmoxHDJtAD+j3HP+0eeti2oKZ8d8rlW98RrQY/ancNFsJ1gLiOzC7mkQQRCF7JXOPMCaKT
sqzCpltHPmowdcBRkO8Nip6hZe9W/5hCHthjtG5zJ46rbtw6Naw9d3popCwxWJFmb1vnAqEqZLDm
wbM69+nI4rqttDglpxFDe9JsY40RfJy7tXVkTPFEcFofbjU02a88nXVVLb6wJrnDjciw4Rh++KRK
lAm9Sbjgme1DxKVUbWiwM6LZXGTtPGB49YGG0BhAlUwd/b5YuPc8NIu+uWjR0pQ8K+OULi4XHgbc
Ixq3e/tQSn6VJaL/dFSpi88oZOVrs7rE0A77NrneOHyPllgvUv9oriP2gIfMP8JA14d1ASj8RDGF
mGLqxt/9WbzFIOKbwaxqHt9I2IsA8kFZ+9CrGslBkpvfZ9Qk3pVJAHfxDriVAaowl/k1LPgv4538
AzWb3H8cGnjNzhoyLSkwdMubYiloezH+9zEA0oW8TSJkmGjvV4HNhFejgo2KpiVHO7VGRzF7b6Xq
UZBVMeIS1jL49BNsm4txlSlCwr8BjsN8Ss5FmuBUDA22TqM5gDvdSVtjKECop3QwN3JbTj8X1eoe
5ghPF6KAdPySeVv/58DfbFU/rqzSSAuzWWk5Lnv1fw+/jRMZ3fFTK9ZIbIfERiydZjOsRB+Ax87X
FiLEqKVMZKdjFpG9Akkcn6xno7Oo0wNfwScA4WRmZLcCohZ7uYeYGlMriwjA7kSeKh/eqCrbu+0p
Riya8r7XkG1UCRp1LitHx5h03opykU3a40qmgHBZVR67we1Rsd8S9Jq3+H1rYi9475crzptODuTn
MwWfh6Pq3MxY/e8Vd9kMhRUL48b3eEkmLcXCe86nT5FH3jDHIS27z6i+PH/gdBpSQPusazTvrkU7
SJZ8hBFsTEO45WRDYFfSOQJKxp4agqRim9JEL+pnrhHg9R2Ml+xtE2N2I9xSOEGB1inFH4mmrvl+
cKCMQCyQKByDhOeLyDZ/I159C2t+jm+JJeOvhh0x4MRB5560S+9T4did2O4BGX4f0gL5h6tQqvZ4
LYtnGfXomBVYT0Ycto7Yhi8EV25jBjCrCiPM5wEyawpJqeC+cLSzIQg1Z5Eh67Z19Bec8gZXSPkE
x29g/PON3yAPbVXBperw957DOvzWZDTNVumXYnkJy8tzI7xKZFzRMa4qqqKz0gynzZcqSe86L1JC
+lPM2033WIN+ijbuNb9JeV6tnxy7NCdBj6Qsf9mOhgi5DV1xpx1mSXzEHHvJ6VnhoRtH6e6q/46H
4WTwEu/lr/Ue6dA3UXMlQfJonbcLM7sRLH0X3utNBDlGKaQWuyApkAvePp0iyAD05LksmdaBJ/M1
sjMY1qp9RddYJmni9N+wMJwER27FhQ+EijSqaqt5kEBX1qnYgyOplXdB+upxMVBsmYFeeFw18xRo
twuYqFqdK4iEvNhRu1TE3mXTbKFidmeuAluaI6EqvSjOPrmgLVpCAqfqaeid51t6mZ8/jqEoNaju
iqLse4VQ5fPfANQ3SuEekcXxpiLEypioUTW9QJtYpB+JTgklfID0pXVindqDt+DLbovSCdZ/pGAj
TIRYZqQLyKCDEiPQ+ZY1civTfsEj7FlRl7Q6W3Ga7w8a4l2Q5DYdrFSixYTPTX0dlMrAz1VgQa/E
D2n6EiuXGwxbuzqsEO8z5l63H586moEBpKwsWxmKXXe+qlCBHLUaKKTC7UrQQr6e9J/K1IsnfLAo
ztT3KqZpbvXDhhq85ZYycbYknU4amu9a/YibT/yQzZ12eKFg2Yo5A0cMADMdUimmuRBWQE59mZwI
2mbUnz+mhkHbZgOHFGzSkef9SnHMjVOCkLW4WwX6bahC5eXAEfNhOhLxIErCiHhxmpl4lA2eVsmt
sPiXkr7SprwKSdejC9P5yObRmGP88ZRrG9BMN5Bzm+zqOViJ97Mb8optKA6L3wbwXRCgeh1WUfIr
DlQIUjbeb571SXmR1FKiMl7Nk0rZkykXRYrgcbaQ7kKwaE3Ty0+UglQxiV7lxBIPxwROILA1Q0TL
FQ4QBSL/rPP/ZqFqPoyFErpztcX+qdZC13aOVg0oo4fhiwjRwAnrMjEQ0RJLYfsbS4L7LBFufj62
jeB+5lrvkeBn3ijoE9xSb/+127DteHO9QXo1/QgrGsB8uepDMHB+p4qS8A5aqOjS0it9cYRa5Jwq
hsK5tzB8loTv5KCsRIzfh7x/Ywuop5EBVZRQX3iOL1qpTV739Ud85fG8RxmD6xM9vAXqhv+mbIn5
0N3VzkDZ/XOP7WEKhdwlurBFu9sdrQMIpQSxU4so0rXBxeY/S76zrgq4i3aT3cFNIhArTOM5HQg5
KI29mOMCpNf/QfWmnOljSOMK+x9KM/kh0cSx8FUxa7Nkaii4rVv7Dxlije3/m1tOpZ0w1CfDfptt
9QLkXCWCYUE9jc+XqV9GtW5Af1htM2qDDf02EOJ5PtRoAxlokJbDSuJVcldvgAU/HzMzq2wou6At
uqQjvW6Ywm5vNFeCdpHG4EoZDy6C5iz22spROhha5DOH1ms14ITqWnEK7rMCATaDkmWDdSsZBzLx
+Tfes++33Fn7Ud8cGj6QnL97sxAqUeq35E6XIYN67uHH3tWjvnfmstSsenfXW0F4LzTHgmiUyBM3
SmGOdWc2vQct3mvmqepHVuryJ8j0Or7OeLRZEe7b7kPWDrekFxWX/fR5NYmBLS094XNFDSVGYT7k
fAh1UjUvA4TAU+nmimCm8h+oeOchgnZRkzfHyC1BMDxLY8eetBUv7pKQZgzmusiSLxYNPreuU5iC
qsqSk7TmhK7lsvATbREk+iNbOT+DB43EfAhoL3jw2NqgDE8OF9zqYzf1Y60acooqyOc3/iYHEWhS
PUT7Uz4JaEe2QETIcUvda/6g07sost6TJ3ZCQzEWc1JNqdGEukgpPpUS5V53uLkCyk3hJbzdGDiG
omK4cXlsx9BaUUCVGiL9y0FiIYUR52+5hBHWUpc55ldKxaLh9VXB9USIlX3dvgfGtSOe9uKU1vTO
esxbqyI5gel2Ifi3yxEY5jgM0wQFq68K478P1G/4/xEenuJVkCVETQkjkExJSWcLPJlVg5oX/rpC
bZqCqsLzlXKXu2vZRUqfom1aj35/YpqnyiJ3b/J+5YWIrz59Wtox+V+b8ln7EWo21tn54dUAL8Pw
cxlfkj3aN810bgpFe8O017OrQo691AxxV8+9At9GHkmV9CKc5q0+rZ/CCuCh5/xsPQt/L++UUesX
2j+y8KODTEXl2cyP/iAarZW0qbLT8H5jMwGMvgGVnK1yAD/zPno75lATpWF0bDiRrPS5AJ0HiDqv
izPMQFXpds7y914QMTo0zreakalH1DXANZ9AdA2TXjBtW1du173eCluzGXRA1AYz0rQhtxB3+B17
cREQSXOIKk2SluqwrzXhGeaARTNrStHChNXeNl35oV0c5fXWdHCecDTZlz04h5lKdVMBDTyYNG5t
PBrqDLRiAAGteIVNavuNSgxFlkLkIUq2+oWJU+i/cx7JlF0/LV80sHUSS9AWEV7EWq9kRPpPJ16i
H/XVyCyF2XsN9FW2j7bkTOTK+aDvIf9TLRbmhKkFKZXm/jyZEwnV11zM5wF78XIzvfW1GkPqki9l
VXgOOJp5ibuUkX+b4HHllesQK2qiQsyJEuuCMhPXFDPDqVyOVHH3xzhS0Xd8LD8XVwh3ihhJz/An
8Frllk5CFot49B3Q6WYVgl+yA+Wf06RONEWnbWPYGZ5BIno+T4NamAC6V9xciNMbD8yG2G6+Xwmg
eFH7rgP1BOlryaDdhZlj4+NNdZDoFdi2JoIhCw6pOD6vcCtC+uftvpymi5etfcMBL1SypyO98aW1
OWyIkv0r1wiO5NJxYxWBa+yMDXTXpeQteDM/82ZLhWuZJfIYwE4Hni7xzpUjN20FGSC7zs9Rhvgg
HpgiQjstQe4yjX/HsrqWOixgiuG4OjZGo0AtJNEf9Kanx9/MjOtgUtkjAdz1GENElJmZ+C0WnaxK
aHTMscqcyhkqwhYvLCO5dzeBbHDSYkMpE7Orr8MxcOy/i51u+YD/yayura/f0FXfBbHiLIa/tHOM
vbvPYIEmLOiKszEdGpOjKwGZ7il3QIxzxZbrZncOix8JOk/TraglC85qhSzDVSN8hFfAFjTQTGuQ
WRvEe4WIKW4xncnMUyEOOF3EO8Ajlkcwg5jyPP3dEMgeH3pP1UsvTcv3v2GtK1L8enW26HCpenHp
ZSxQ4t0jDirb862kBzXqHP1PWAUA+X1GXtlyKPZp4j0TDu+YG4TQOTLP/IkSOq7VxRLrZJBNQAMV
iKUDStz09FoUlgTPGK17ptAgdpYDoPs8e4Vhkg+ngaYFQ06l5ZgwtQaYyYpuG/U/DuSWfyyE3nPC
sZ+mnwdxElianpKY2YpHQi7eur+WtRweNdJKocCs1JD5twgcrw7z3qAn307gp68xW3lsz/PGQrZo
6ORW7fHpGBHMy5/GT7mNaMHfKrrYMXohaOSlFABf6WLCvsgNEW0UCXMGPuhIxSvZlcTnsXW7x6ue
aJSZs32AKFfuCLZURcohPy4z58ihrKdmWPvt1UxP0rKHXymlvqzkzO83+Wi9ZSyN1TuaH5wCbcUX
bTYr1VC97t3dGj17A/Fm7PVNZIUbI5Fo2q1jRMjvvDApgKyy2Xo3aKo/MqsaCWNmfgn8/cfRh3N3
sfL0CWrakOnzCnvnr3mJCyg+KOvaDx7pxMtLYv9F9JfJpGqAeRsoK/P1D0KaPb5GR+vJ6Py/VnKN
Y2x7PR9H7sP8UhoHWKtHdjdGiUa9HovAUiK1Zn+m7JVhAGpofEsZB/rRGlMZ8UyLPYmt/UTfSi00
OYyo/OEhcIa0P4SxFpKQAYRXo0yL/T65zaK78Nj9CDstDBxcvTSP02JQiVT6Q3RfG/H43ogPru9H
9vecRRzI12OSqY+7T4N/vzt7gl3loQRhNSxT46CaTgxcWXp3+V0bElhElBU+L4EZVS4Rgn+uOypn
HMJJDv7BXtG43UqOJyHNnexO/o4wuaOFr8e9xMec9nQVEHvuwQ7w1cYO4NBiutnwIF2ApF9vQUP6
mDcUhw2uF31U/Dc2HDqNbxH5U1buwORNb84RGCAHf1dGUHKuyFzjLtezTyJIicHOEbRd/Dr1S0Xa
M6ass75Bndud+pMdDLdnqU3gf31Mak9HsqOjQkZTcbI/n/xn0s4XBDH3OjegbYkb1aETL4xjJ1Bv
nMPDAF+rIYeJrlTUIrKyKiw44iPELLp945S8UoTFtyTYGfeJeZF4jNUW2p7DJv2PrMiNPPa3coRf
4MdXczzFGv0ol2W60xzOXY6DDq7dtXxp/LuH0FaPVBN2DdW1LllJryj6/p0/oSRxyb2tDeTAesB9
HMXAlh5752YEo4XMEGM/0NNiBWs3ZE6bVgBDAWC5a1hbX1o4g5eRK3hZllDli8VTWmwIXY4zxPF1
EJmxDX+t6I470Ho/obibRfyrgc0ldZfAMRB7vXrQchgC70el41Pni/XDYZFm4w3sSTo3Gepmc7bd
XF1qlRcXgMIZqoOjI/VYrgTUi9/eBTmC71pcyVlFFlTzpsgEGhAGWk8wi0QrnqrtX88EC+kZ9imA
OtgR5/JBvU3nhAiNPo8QaQfdanAt9Vl3EABiXHyNhMC1x+Rqo47cuzEjiQNVIF9LzTZlvTmnLs15
Dgiw80ELOsAx/SCClpUwS/AOCAwYy0ZbOfVYIjF3PPfMMlTQGwjWwr4AspirPOiY0rIzCG0j9MPk
39kBt1WWExbrO3RAzZAS5PaXpbAWgaCFPVvyfb+Zinanst+TE2BHLezb0K3RtGWcllc6cIAaAh7s
HO9aDBbZCBqqBwKLpljl50QS9SiSirDiVTPOPgq2INmVK3JJ1whERtVKcHD2pXZVqVCj3lNqrjGn
aoXgF+zrhxATZK/LJT/8FhxKcRhFft8oWIUkcN+OtXQJ5C2USTnvu5Gmntdv/r0Y84ewt9cavBWG
DCIdIIPvVWnIEH/alq5GvBTqz2SoKR1g9mq2ZJvYx7DqvEJRUOj6lYNrWL+UEnNAwreKpGrZke1b
/aujdFqEIrbLVTjgThUBSeQDv8lC6Co8ouG+mqaEFNAzuaeYl6QMHOopOW3FrUfN5wcT3poEReDN
V+p8f1wL71/dlammJPRW6EdEj8h9rCdIfeFkfdIZ2IjDsuqzm0zwEeyut/Ajlqcaesnk2Bj/MisE
ZkQNKhtCZER6dhquy/0TOdXFnWcJvshw7H4uDjbiilosqo6F12yrDy5bGbf47BZUjYQwC42LPMio
WOGz9Z3XxcD18Q7dFrFG9Ft5CuJVHPMMK+c6Qy1ytd8mBwWjcIGUqm/YcRzkLodxEcAUIz1jxO9p
UrOXhu3bkq8rNuVLhrly5SgIg5ZH8tq4cLFSMjZ1IqBEvD+Yj6z5CI/p+d2MFqu5yrMCucQlaKX0
BJDUPDNDg4D9+5ku+gwxDCCP3xTU+u+sT9+L29dqggaGmFCTi05+DShbXmITsXoiewUwDR/tjJ/5
dlA/VZLgEQK6voU9qunqt8ds4NotwdG+KHXcJgeEzwxGTrDatx5sdkO0Nb1s3m00Xhn/LiWmcQM+
48BdvKvY14KSi8s5bNJl+h9S+675YnXcrOSMya9pKCN3nk2cjTkUPbwzqiT/jhG4wTnzdkyswmcp
xor4lZixGdkj6T6oSCmNs+ewEtckyNXy1w9zrjXSaDT4veyz5eyuZwlIoOMi8HCYLOpwMsfoV8Qk
wtc4RojdUmx9Dq1rYzyhpTQBHq+NGADoCsBS40YM7CYWPp+kBmKD1WJR2ORgqsSQAB1LR74+dwnj
znhWepZYObeMqT8rZPp7c1QQJiN6hJCMf1fov3hltUnVujQURrLxdHmfrtv1ue8IYVUv643O1LiA
PYa9Qxttb1mlPyVpkSxWkaQLQDOmWtQUD/ZlD5NoFjablB8Q2f0DaQ0eXHTRdSj/PLSu2UqXvHhR
KMC+tGSWNvg0Kgo0pCLsVb5d7zVWcmTUiULNpbS36mdEPRV1vn+pPhJ8p+zn8GgWE7ikYOwJ08cR
FbX0+xj9oqkQIcCyJxGT6OePKoozxo+T1GAaOL1ntLQZLmA9SrW8UzZj9vys3mIDSyBOyflZS2+Z
Ppg9PQi+7dbdIhFsLHP1ed/r4ZXaxpK6IrINlSLHFcr+Mtg9PVuixA7ecsqIfegbjsY3Z4/m96w6
PboPqag8VUP6W9BD2EEeEvalhBCHiLbxZLBTIi0WsZgrO1tCElntwUqruiRzQLgPvby24EYqEolR
74Hcjf7JTinVePW8w+sTjKEVtNM+vUUCQWSEEXsNLQZhjzQr9dXi1WmcCA3DVHLqQeSv0poA+Cac
J9XcuZb2iqUZQ8ixUBdiJra9ZAXpNqS+lR9FsJ4VuySAtMBEX7Gb4HYbET3v5StF4VEtPeIywbCT
U6F1Hni08Kea+6OuxVfbJxWShEyULr379qpVL4zQnCn9hmdP6ZLybH8wWWF5FKTvaM3qbQrepWhj
cYdQmjgjR7vFIU4CGGNdw8cicMqF06WHd7XwQQaVuidYHvBvoFgRuoi0XwsTvRG74Kw8IB979l52
decuH88Pez6bzEhP6pGGghZ9MPGoxqPYhxlq8/BMsRvFvlzUXs+4O6RK66/AqCU2trz4nGjh30iK
+rURb6O3ooFYG/OB/zRZSeP9D9MYqK7I6z1C0WaS4qUqc76KkCygFrhkyE6lvLcBjGBekhuUpAC3
jeEAtuXzhc92kjfK6QeSW0mFANJG/Ii4prfwFJdCbMkYHs+nZH9X/v+7X0fYhKQgruqFE6BC1eDs
Qyp5T6zpE7O7Sih53MS4gQA8bmcn2tzS3GyVZFvXuiLYol2uwY249s8oaVhfHxTdOvVTqI65fXvB
daFVEhkwDYYNopeki+rL7QRZ//ngkEs1uherGrhZrIBMU4sHO0nA34ZTV61ceySjElTRCEOIbC9J
64oiL96vsW1gtUGXUgJ2QL4qZeowD86cYEf5uDeYZRlfCWobTBSr6bYHnyE5gstU4bD2i4RjMWo3
jkvZ/gE8JyMjlKpNIygehRepo85P5ib8agL2N5doH3hi3ofhbBh8n8GItqToO0p/TwEFFP7Rbhxc
44Q9n98L1wxEui5sJILlknRjB9JEkd9ILrxIuCjwlKB9Hs0NvBMyNXasV+MuQpAiSiHod+O6DrCV
fX4Kep9yQwwkf2pXZ07/zO/KaisqtEti+JPIgD4/0m7SxZgT6CjAfX0mk5kao345thB6I+n5umN0
7dWHYzPtDi9ySZvoAiV6NPuF5L62hz/BLQCfJL7rh6/lBg/5BJhbwJ9YUzAMCqrTqiiH/fEZchfy
oeQmz4+dKXaRqwt55rRuypEW5oxVU7aYkXR9alkg9zLyGe2foeR/yzbaUyxEr5S+266XlKKX+9ID
R1B/vqu9c2l1Ba/6OBzDXaIQUt4bVfIWJgteTLk/ANuj70wk2mfFbh8RrxHkb1xWd5MDluKKRpm8
Uz3/UmAiQ3UebgvVb8+3ymZHSWb4OZFyxd518wVQaP4sDOh3uICV1nJlxb61X9R1t5nzbjn+TU9P
zC02feKvhR7j6TxSzqCqgwjSzW+Uc5Rhzijn+JLTbfwUGlWHwBZA8J5v5udO3CZNjojEkmU/0DY5
F6S1bAWYstvWUSlCAS5+2ARulFBcpuD97zK0FQ39bR2bKdDrCWyFY6JHlzdy1fkI6YRJ3RsJieDv
LkSjUKlW3yI3u3a50BalN9Org3+eT666wIcHFmNzj96G0QdLEayu3VLhG83XO9+X3PK4Ge/QohJQ
qft+FwHQxCvNIS8SJXkjNSgrI5tf3w4s+9FQyySQ1F3HMXrMN3Q+lTHaWutzyb142lXVWkVw6z1Y
YFFnBi3BByAT15tMuhpE/ghDJPMzZJqRPke7AgVYpl/O5/coU5CegcFzygfeLL3qV6U9AnDFZf98
kVlm7O/m43TBnreFQSpp+6vhOjZPMCJPxPFolF5dPwgoZSDndSBeUKRGErFDaSfeC4cxw35oV/pT
2/vpp14KCsDDXRTwHte+yfC0CITUJOuiRdhZXnj7fRN5w7oeyqbBNpF00zR+VGN5IZlb59wFUjYd
nZzuadK6cvbnP5sWWUyAXuu3X4kJP9DW4Q+OiiZ4w18YFVljSfDzHk7M6m+5hGMGbUare6PTs7yv
VrZSB2DJ5OzWASRVNlr6NXnkcV5TTe7qu+0AGzJYHAUPHSuReIWPAJxjzi5X/C88rxSycCmRaWul
dMm5xDTdO/3E3FwTL5+7auFDuJch7cyD8lC8vlH+n1XiaObsfw1e+0iBNVXrqXsrAMy482IQdn0h
6SK5ddW4wqQZhtYAQP76jRZywj42li5zRY+VV0HpUBNMWbmoCCbtv8T2a7Vu/4Luy73FVRO44XfY
TRYze64Sk69xwkEtpaq86PNtw4U6usttjcg6WbmUwrO5CryQYkFwexjg+cTzT7q+wBz+af6/xwlq
wX88HRYbSVl9rUsDprgozH4mbKstjMF2/BzdUGmaNEO10Mr3Z0QG6b9fa5avsfIuBW2lAWOePi45
LB2bTynnLl6rW6yNMB4NH80NaBH7wC5rxH7VDpq6fUSZETRyin0QDWz4/a3pxED/3MI7vuLHni/a
1JWW4JaBcADZ3uebEob8UKqVCXMU/5280uWzzTQRcMT0yFFMFkhIh7pmKHUi+k8+PFUdBr6PdlmY
LYT6s9pYEy3aOKPITtkeQSYSAzFR0bIi7Gwb6lFPNdGuBDBrjZeNF+2lAv/qOI2x1UFif/CqeG0J
O1vU0aZsj9H86P+esbyUdFwV1W8HpW1myxsyxoVrWqMck38RXVTgHYCIFtZJigAx+YY66bXA7/j7
cVGmSP4MTy7alaBF8x4alwY/JZR9EF0Z/mV4tBnZMyfA5YvF6xndc7uneFpXm6hX35LqLm3nVDvP
lf4IvglJa4q+v+wdqbNfnn7mowrG3E3bkRH5qzzePjA7LIscMGsyW+Da7zwQCTw5z/4QRP0vnqNq
7TcWbkBAzPhFcRmxu6bZU5vo07QfzhuZ2PusfFHuJOaLS2iGxRgVewFIgrmQ8Rswa7KKGJWLsGqz
gn40p9ovClhN1nGlbUbpUFFp0B+mhAlBPYDmbN3ucZBNWQre7DS7O0LA9GN+LbUAKEUEH68w8xoW
wXsKM9dvG5GjkN9TPp2vNk/HqkbnRUvDwQ9ChR07xdBjGkyULJzCIOtBFGKlZZzBIuJjCa1ntdYy
jzEKVfIatLYW7nTxzirR9QsiUoFD+ENNlfZo2C5KROvrxk/xENeq8JvFEgtuHheVNtV2gQJN3pDt
4ev1jgaQTuXj6pKWq57kQpN8bTFLIEyNo76+NhGALF3AS0peBJ8e76LScKNSpCgk6MJJ5lvqjMHo
JOOGYqb5gCPrj28V7h96M3GbLNXGY4JHul75iK67bZI5VnvNInmgx4SVpXnofKncuzIRVJP8+lvw
rdftIBku5faZiNmrrWxiNgIbBoXbfb8/XdU4l6r0nyRpr2BZJo8wURYhBNO8aBZZQgCzDgGrZi5o
V4rW7jWi41fHX8Qtbul9XLjqrwegwPbfomDXKNSuWcBHFVbuYZ2B2mS+/3T0qYlNQ2h1ie9XvOdi
OQ5Rm+LxNsBMRu8eMZ8Uo5MBO2ius1aQOQqh4Sc8k4Q5mnPAuf/gjFNFZ7DHqeT6kj+gti3Hljow
2mofMnNiHWqohyO/npY+GkpRMZoDixjQqrznlwL+X8uI3ggsK86F4vcfXdHNbdLloHfb6jNzuKip
0AMtd1BNpT4ywdpWzAteyCwLCq/jQvnrLb3MJ0XKgtZetxbTnoT+TLUu7p3lo1PjgvdAi55BEfgm
mOayuq2H2kdOr39pO6qr2DlsS7ZwrDepXsAFefCHMVAsYkZKZZ1Fa1nDr75QaLL0sOyBsEKYJ7zL
PcwH/3lPWtjBU+3w9u2pVUl10b42aFfIQurTIiqqrD8Ynk4VWCTP2Qxi5woBKrf7FEllUNr4jZ3E
ezpDQTKaXekw0qbattRhpS2EJTOFb3o4SbJQLjm1Mh5fShqbHGWNAwaTJUS7Ozw49Um3A4TwuU+W
z6NkWWTV3ARmFRQ2gM9A2+D+vi9U+hv6n4ut3Of499M88xq43veuIiwrNdN7iokeilECbDq5Vel+
NkAMk0Xc7ISq11JmNNQe11l+vzf+DnAtL1eZ9ixM3hTu0ZpF3oBNVOoY9ecZbC3EBkGoE/hMYOx3
9rF35kN06jwF2ONDIZXybXyv2Gjab8epKIxx7lGpN7cxWNpEQQEeCrll+i+1TM8QYL9QSeU4x/RQ
LcPf/6Q1/V8hhLzCFEeXJn/RBfYt41ltU0uSqRd48ylQTLO5DmvScaCrqHr93PUStPQzjDm/guBg
uUDnVuikrZJHN/XKsankgShDPMFQz6VUmtYz7QMoB87UU4kxsj9qoVOWPXBuzJdiZujLB1e/4mnf
faDASU3OUIQiZ+BN5VfAfw/XpHtfiluR2dJNQ151p5ClHqyKcpr0Gk6KntR/0G9bcLi6B/n7B40e
RxVBzx6rMRaRP6fFEgS0h4uvI4Y5jOah5bSg0bc0/MkajGOfzECwxlryenYakYI3dcS5nrB7/EyK
ZdF7EKsFJV62RwkZ6dp+YqVIqgcUS3u4n6lDahKBEWMUcairXpXgccmZVkC/RmOBJZYjc1pU08zK
qaNeuIb/Mzy3y6CdPnL0kgTe36XL/zqEjzhB2V2hsP4mdyCTi/sFSPWe9abcYTNcbIkcq7VXsjoJ
vEbr3z69iXZ/PpBokulkpcqzxzVLzzah5Dn+Z4sugrPiEe7S7w+o/13aJ4M4/KOFsUv7nRBDK/81
WyJRlqc7Siqg8d06uvdjPnxld2h+guZG8tqdwUYGOC8WaEwBKHtp5qYwagBbeOLfiszzXc52EV9b
6U6Gc2jsshaMDWl60I8/FYQoDyLB34bNQgCdBwh+UbEU2oblKEs8kIm/4HS777BgL3BPyT+bxkZx
IrQ9wF4kcI80u33Z0R4YAv2m5uJbPImuTBLFXA2Dtqi1SFtax8gWsyV8JXi736qSxngiRW88aKHe
6HLF+Rg0spe7QwekDRotpAf6z72TpfR/YuWGjqKkIsQariKmjBkr32/GtA0xWL6VRpwdsu4qS5KS
jQ4Gw79M7AyAk00AAV8cPZY2UneTFnNPE0bJFRcgSjCIJVKiU0aDV31GED3v5hx1I6bBt+NRsHgY
t9Rj5k+DEJu0HNL16h9q8NDs0FgXKFMB2wIF8wzyBucGmFkZ1pxiHoY1z485P3RqLsoxy/x7NJVE
5ehfNZKiEf6trQydzKiQ+PcRYbtUOK/IjYdIbHu+FtBGfQjfLJKOHwSvTg07SooBX14mSX9rOnwE
+raWhnGKLhN5nPXcL8KhALa/8tlfScuJw7R44e8gAZMuUgZ1W8kN8UbtyPwGkWRArkCMfSRMLOOr
Ytw35L2SwdO4fpc5N01T7qC+jxqa17mmSZoY1h3cC6obTbR7/cp04Bi5BbwuD1trr/ZSjaW5v3qD
BDXhX/62F42D51agNoIIkqjeh15sQ/YwEjTE2gXj7dtVRDgTFex2J+4I3NfJ0R2moSPRrhQ4G/FB
nRAbGNqHpPmG+ZD+E/mlrf0qOvoE6o5r8gpX1q6iRqb4MHJpe2HaW3nT6zHZOgHHbOG6IKsgtUmo
coBakSQHCetsotct7kQ4PrnMwIOFzwgWKdkR2kkZiZmwf1Pu98svVHgaEgXwLiWDlD0O+kTal9N4
Ypmi0ezngWagyAoysW2VSdro8i2V8d/gqsBTlzSzoIIrJ1zvWeY6/3oYgkAKFpNm6jLFhquyFgBR
eoFmfOJoh+gzZ3MYdWWnYbe2blJhbKrRLs0QaTZ0Xv5e3h6JWoSyrJmb0eNvXap/T61BODHTHDZ+
oGHS5ys30oA07+cQt0Gg8gd0uRy9Qv5dv2hlbO5tPq+K5R5zzakHSzXyL2zueBPR7D5YG2ROrrWm
yqEWUjSPv++Y1Oi3EGJTdhHxv5KcT4dyDWhGzrMYLuwmV4uWhUzkpKrigZ6kFsEAVQ5o/3tDYhUU
ZgHJWZyuf7gGfDV3QLNMAJr/rSFLi/FWM5CfppOCCBawuP0XnEV63+rk3ASiazCPnKPRk0BuK3RF
yomoX50aMuPyqZoVVM9VmGG3j8GicWIUxAAfPAma8peCBfzSm9vvPHCSTv5n8iuKfQsbx67nD4zs
W1ld+dOXbW20oyKUYnW5rnrD/M74TaHx/pwcMIYt7UTKAKCDXQZZJtTmw9E7k7TLL3D//QeqeK8m
SQdiipnmLmWDJhKyhpep4KMZyyk0Yy88Xw8XbezI8d1nIgx/qFBH8cvMD5nLUX8r9L1KeBYOyAUd
fo1WqO3GfZsqmI4h9P24/J9dEbTXCsp0tY1wOC9dJDiS7gHUcY8rs/RzcW0zY8+MhHXTv2DgfbNM
mqNwK0wnjVPMkZVIMjbWw7QYy3gvnic7g8ZMUsO7sOIIVe+D9Q6RfGBbdVaJC0CcwTTmGN1wzQhb
Ge+Eu9TWnqQgmMLkfAi4EcS4JdP8LD4mxlkTSqw2EqssJ3XhC+GIWrwCy3eVbRtc/aM3GqqID56e
AToJm3MPY4KxCDnyA3gpISkX97wE1rSvNO0HhQhVHzB5lgAGNv/qbEctiUnYXbAID8mqVxvapwER
9lt0I5Cnp/vzXuOdpUvdsmHpD2kvLSBl7YkXLB22XobT2wdmt+Wu8n6fl+1j1/iO7igz6rnKOGTN
3yuIE3W8h64w6uwtd97YGlpMXvsOQyi8iK2Z/K7dRtzf10eeuDylw2l8Ly8TMkDOSmr9RV2mt89k
rmqE/TADDUXCUqYv59rkF7mnq3KNA8mHwvJ3meiSxEkuRbP638OD8K+i7xsfTnwVbOXFeheSzyAM
Ri2t4hHg7kQPB3kQUoTPQGdFcySxOgRvLMkxtVA3V/n0RklbsV7sOUdkrxg6oBAooamoOPD5gdD9
8Bapb7MiokxgwffqCRfaawdEDlL8j0DoNbO+aiAWjppX0wtckUsJf/NpSbR+2rPYXpzydrJBeVYZ
ydw8gb/2H3yJDoeOLv4NhC7gmxhQm0Spb7GgMu4PIjTxLu3MWKMzmZSfOz3q3rsAuXFR4fw+Pah7
vOID43ITrrQUkhmieBCKE4MGLzMgnjxyhVXTI423hHSuwZiYckqntHKzIUT37rtOOQxk2976LOUo
Mky301Pod8lTqIQoG9gL/4y5LRc8s8Rqdart+ezwBsn7Slg9TUOLQr2TT7buWhKC4aGv3I2uxrYh
DV4Dj+jXYLa2JYywU25MgQZYA1iXXnOSjfrPJkfSwSL7D+VfyofbG5z3BhNloDO8qkoP0dKItPul
ujBtVDy6VXqsK9CvvdDSdyO3nab39pbBSFkvyn80+twu2b5lvH2N1MuH+RE9S+lWgTRdITzCtPF7
lShfOX3nilLpeoU75TIGN/JJ214SA6dT6J8AojodjAwiVvP/8O6G+1kaQIaPdfWOEv3cqvt3A8Ro
IGPMMday2N8ol4kZ/rgcHfwcn6qlbJNDo9d4D+6ROBulHILWMSLAcpTZVNOQWUJY57zNdKtujH50
uf+eN/riKQPelRph6PnmSA22eKJpNBQ0vmyGfT45a3hY2L5Uqd5xkSenSTvI53BrjRaV4qOZWZUw
rnCRX8gsmnNgNlObzLCGiagtTmbOdti5iZKALeStJtKVQulLnpS/rOvmI0Gepqh+Lbg6sKKrUIZ+
9O89+mWYLSLwWEHDfuhf+Adokyfw+326U7++gvkzewJRmzflTz3Ffpu0TC49M6IPBIn/IEo67u9O
Se7KrWBXSH0FHiAq5mIDWKsFhFeMC1DIqVdk5NC3hMR7D5QJU8BEtz+/h8oLsluxBzX/5UyE5Gps
3GZNJHgASgZIjce4c/8WroIx194jYf9eUOwjpijVYgSZ/9EYcaEMuf2mAOYGLo5a0VlznE5hgymb
rvlST0I8NZoYpJ1nGxUjdhKSoFaKw3FwervzlWk3Ef/IqaotoC3wkSP32W6ueQYV0TcSnq/UEzet
YvNMpqWLNVEDUI3MZsdHL/NYxCE+9OPH9s56WJFs+X2ALEWj8o+AukX7Oh2ffiu5/JNI0CZiKb3W
W6VGEpUEH1HbiUOqt2/Je/7ivsLDHoqWAmoLE/xBcYiXLRfDZK3i9x5bVJn4lWaYcwXDDs1PRM/F
X/Q07O7DQ9GLJHl9kERTPRFLkjXf6i6O32Qh4Nr67L/Ixa4xwonG/7x9fFmJwq3hZn8uJ9MLuJZL
5XeN8rSFnVq3gEfSbZTvPF0kGCtU0QE+NMzym+nWnFpK5NqXcfQ8IitwEm1PwSAzqzAkqNg9GfJB
Z4+PaXeQFGafG/sC1jXavmICv4h1EbCzpl2CX5Ahl5Xa3KQcaJyakEjTbrsdtBulokquhwR9vnuU
PFxdZV8BRAd7BFXpyNgvVFt82w/n/J1juharbVOVWCpuJuuRP7Ny7tqIWqD67ktgCIKbaHwR2oml
Mf9+nuvGgPsJpDcKYTZouPkOwbJ+g3uocXfpdAPsAayICtPAfu2mMfVDkl63yQQR8H1Fj33jYyWO
I7UFcSXEi8bFiXM5ddSFmJ9dtZFeC84SWdTWga6uFTSDs//o9MzNuBsSBtyeAfx9Ca6d5sO1v1/Z
EDZ0r452u6fc3moHEyyJ+15ntoDTZc7DDKU5HbA5DZPGfyeCb1bL864ZrXS2Vzt4HgNX4azttJf3
s+xnQzlcCDF34Ql/TwLJGMsr2P/b1CO3s+DuBUsl7Ajwv4ZJ1CxBZ7cIN7mKbcvex/6TgIZy2lK+
Yt7d47mxI4sbOhW8RN40smjUCh4OMLvuSkMilrlJEPqQLACVpR+ROPOKgqle45lZfA2J+BQB13mj
EgGIcol+FMsdLzP8IaVE+EapUmy7pYv5+R13x+qkoRcEpC7JTMbUDZYd042suMx5ad7iHvIyluXV
S8sIRUkZI+iwADA4N8O10U1oxHjpFtAl+8q5qpp2TVMoEamDgnKh8wy/7QzXLnMrMBk1aZJyfUe0
DaPCpJTmN9P2s8v5BxXvbcnywXlkQBdB2OXH4EtnhoMJNyi7NkX1FWaYIPikHAzE/UNiE7wA7LFt
Em8t9SB+YRcvWcNjKLeFAWapFmbzun7/0pHKhEGjGW4lZChH/plB7FESblH9+QMOj5X+HFNSocF2
JIoiI8bE1aKFwrFdP8v1WbGvIkYWumVKhErmuoJ1b9hiy8ukYpQdBn/DB9DvvQ1vFt3Xj89Fjh/6
Lj7R/QxKJDX9HoEIK0Fq3ADJxyA7Hj/J8Ws065sC9/fK34x+aX6hC55KQAwl3vZTVEcJjdRjl+vl
tR0m2kXbGO4qAuvyPa5pCorQUIszCEf785AQNL0bx313toGF4VIWD5cEH5Hj5z16eHxMa+GXfGdK
sodSNXWysm28OnUwEw5Vdrmh3LJIMicEFfjMmKRwRyMTnZC4kywmIfQoQszSMTO5L0W3Hg1yG/2x
1NbUY7wMUmEz7lBHxI7USNlrDn0aoC3G6h4X1TS6L+f8COD6WZGSb1uibiDGQ4JP9jNaMCJidiCs
Ft3mY2zOL6f4r0SeSQN/GunHsa02BHP1yQU0dwOj6G/kiO2pEuJjFCBk2xP0EyyfIyZiIhwYxE3g
gCTa0zjW8Y7C4OsYT0mkmBs84amTENfpssvG2XKcG87eoR+pXmVR2d9iO1B8QkLqXB3wID0JUSSP
PMXeeoDPUKg8fSEdX79527Q1ZVcXE3j+RwsxaBcKUxVuqIK/jY2Ms9i+zPfLPf+de1YjZXFkM02N
QDHJ0NhsjDqjmn7YZFLW+aI9y2BF19Wp8ITI1pKIv8YJlCOOaWJCjOIsWKLdYawec6SsiTQh/q+m
ZNavMIOXOc993OgRpk4qKrwX9eLLkiN/55nKFqblNRwcoYeOi+BA9be8iWHJZ+uEtlzyeeZDlBLv
o2DjMQpqUCyjAwnipxwLv5pheNrtitoGQamVKpBO3B36cZGSvNr/6Rjvd9i8bw1bpYz51EA1IVY8
txjXIY1iLnXOObUpvp3Zc3XemOkzAIlx7Xggg1lD7vfKhqHyaBc42+dkw/DBTl49N8Oh3PaIic8t
6TdJobeOJPFf8/P4bEkUxmwmtcieyJT35aHPrdal6KFMK/SpwNQcp0Fb35jjEpT3wyOfFl8z3OMR
8ZMg1nqMtdPvcLL4lZvWa3CtiaaKI6A0c5weh+DVIKdL81/AWFAcyWZbeiNWWOPFrsaPaWq1XT1A
kywA4Bhs6KXqWAv39JjCvfQKS9MxScyjNF4n9bPZ2VsIYwHMTQoGbVTGaFzkfiZ4Bg1Wn/zVEYx1
5er/6i/pw6o4wcdIBcna+W9O/FdyPiwyVOIJxXvKIGizvUQJsCcmGYce4s24UIzKFX2oyiA0ZNKY
6FFXvt4WBNRzMHf7mgMi9/UB574ODCeWTmuk1Y9/oaC3MP7UbdVNmGZFca3mm62kCSQ8XV7KPE+X
/UznLIkTT47QohZK39ltJaVtP9iQLhpXd8SdWg/Qnn+qyR5zjo8JXuEOcdyynoL/Kv7DF+dNXJhz
k7r2+4b3OA9H2GUIFv3F8R8vkr/Uj75rgXVzOJp9jtvebto5+BgATG+Tv9jW1zSgiFUFHf8Xgjau
Q2TkUMwYshcfRwtpP0C2RoAI5I8pn24R+ZZqtsgF3T3J9kS/e3S1EUDrQusFPzuAzw50y0RwO8c6
aFx5zIPHA5mKmsm2SJpx1lEuc1FlMHlPH2zOfz0p7/rbuwCYO9eyF0nwAdbx3IyDUFiQqrOETiU9
EkHhqwHxKJ5gRg6H6BgvrcRpOXiYYw9GHhoXuZT4KpZxYddFRivKTQl7pFa4BHERX/mRU3IueIP+
q0fyvRrTMTaMpSqEON2nxCSxwAs094jaw5xz+RLC7fmmCK2duD0hl4yCJlCu9L2zOgz4Cj4VQHVc
53GkRvif9OyrUObFIfz6jI4KqX7YgMHvfkIFgKI7ZeRvQnGvm1CObQb6XFCppwU42RoqGgEO4B34
C1XVA6KAfaKL0Za+iIY2CfKCLyIlAhphbG2+lN3k+yGii4qzurkhXYbWRfG9DrFWPVJU4g2DcWiu
zCX18qH7u67Cx+amjedCx7SqVSo3gunr0bknpaP4DVfCr1P6M6L2OmfY81Tul9G5Qwm3x5BhfsQM
p8FsszIM96Ptf3dK8EV/DCJ3j7axH0YL+yPvaIhpZDF2ywWXg0KOjEB6txL5LK1USMQdyXGatZ0A
41/CiKK/PDlrbevHhVcO7E2LlA+JHLzwd5FNRnWpXYhZoiOSZBlM+nEyvAQfJ1J6440D/B2W1BHL
2/zTYDBODiczxcHfp8ZNcBf+foECRGyppeGGC9uaFx0x2Viy7F5fXtK/SsW+UXkUc5gsw0yWP9Bp
SH/N0ICjGQWK1wbuApmd1VoNgD7FiGRXl9M5YLvq+BDuyW/hfB5y3vEN+ytAlJ/feld1cuZNIO8S
ezBEDMSXog5j+I5/dIxOAor0pnXAvkC3Q+TBwaYiCVFVHq+TpLFj2IIPYYzgJiiWX4zVg6U3XUnO
74mr+mzOX11E+Dl/PTSZV8U7GltOAAAyC4MI6VpFbuG+qEwBPEUH9nFpHg2p6QNX0zFH5E+2Ah8N
77N56UiAhkKTQBxnsJsRnAgYUY86BJ3t6mFJLXI5U+kOHeOAkn/336Un0f/v9rEShmwQ97TdJEls
pX7lwxyf1OI7totNlB8r9INWhy3DK3Q5F9xwjLf1aFzuxisRum9A26pgZwjkc9a6ACw92PNEk5Gy
BTDZwZRW+Tz4meH/K/AMD5v7Qi0dXRmMh2lYZ8m4cZhJPN8+4MoDnxLoPBu8sQMqVEuZHyz+ap9E
jk8gpkX8GNqjhKbaBSb3kLC3onmAcHnxWulVeuwtxGeooV04xe6F8TEeRS3L03i0kNz2C/B7jtWy
jbD4GKcYZMoa92MZksyHGC6PQjGqhDLBQHzRJF/PcBme/G4KZ49cicLTLNnRz+OP8oaAJONsX62U
jH6TURhccNb90LrDiag5sGt3Bg5E7xLC2FT89zDZrSIkW1p9z6MemP0yNhzNHQXoZyfn42eqh3vu
fhW/496uDZyfOPtIZbKkTSkgmG5LPOHLUqBHLFd/Rk/eRSliHEg/zk7f2Lkj0ojaFmi8lOANnqog
Ma2ikaefPW2zkZXby/5qfQrUurkMIbBDoaZaLn2zxMKu7BdYTDk6CurRndm+f9dOQMiwE+x3fTLz
6hhYB2WhgBmqb//clTQUI//E1LiB03x4b72yJHwmVYDmpP3ScOGrrHv10LOa/qiJs2QKLt/05FnD
WSfjsnDlnRb0Qh9MRwYvsgm8pWkon3DHyl4VDtIuGV9c1hjpr/1gBXO4osToPltXY2/SDgRDLnVN
Su4iivdMk+Ke6OsDpfYByHjImR0J96Uto49yeTkNVOfFxYH6aYZSgjzr4fH6xUz2QwCTVLAaGfIa
2SfOX2QcFdcPxwZumRPz/M9o8fDxEl+uRRpEITmEMznVZkYVvp7RJxWYS0kMlVLithRkGr0Ziex8
mS2VxM4UjNDsUS+lDZyNk3gWjHN2+OMV+gugEFieKYKbtXxgY7I7GjT7iwjMM/DX7Kz1kUoBTn5L
HTjaQNDu1btdqEyUI4emmhO8umGppOTQ3te/hQ1nQzfIwEEo0bU8p1B8bgZtqlY01tw4P2brlys1
3/Jrkg+rxPi33m9K5fNf0UWB3MidgbtNDKvsEE5bjxHdQZd6/XavW6je/6jliq729PY9aeZ6sKbN
0C542jJbwM3ujTVV9LwpiXyfBpS5E12Gsa8ik/1HIz93Z36r56rGyGhFp4Eee8Dgv14ZOP+u0KYT
QEDxAKHs6MW7obCGXzDVSFAW6MloUg/SkBr5BavhpwjO9p+uxrxm+MknTNvGa+UOQYmIF3b72RG1
32X/csnPhvH/+f4nMaj+N2t4ZOB6uqXb45ZkjUw4D1KchjkZmivBal23ZAtBM8ztQjLG18iSeLgU
EkQMxRiKW/uixOHM2gsvGq54A/+1LXfnoVw8+H7kvhcO+zbP5nONVWxO2YJ36+BPJfenZob5WgzV
eyw631b6ABrlcEqcwNeTcWb1JyJ4eza38YQ4vA1rrG7qHwApwq245wVbb1i8QnZPXYbdtb/WEa3s
d2xMoVU3ooBtRU8UuRpaooRZOVPC2vJQCZ+LSPlZuTOmbwlgTA9kk8q8Sw5OHsFqwsu6uivEqge9
vcjPGOdz7Uh5XlG1DMmHXy4+vyh28qynhXvQcsFF4GgwDMvl/rfBzIxMr1+IeJYLY38xyRAFbQI5
HWKQr6xoNdigG7PxXwvUQqjrw6kiYbRR9Zfe7tMb2LSrseJ7QJrk8AmZ/7qhXMBZA9m7JAqo5ovI
ICmI+nXnFK9iyhT6MTbXhuLuCrCBvEJGNNsuwstcYa7ehU1iQhafzvQCx9ykglMHh4U2CsW87gvD
CrYpp/GH4/lWleYAV0z/Zl3ScaIwUy6oLfUkZW6/KUthRr8dkjvuTwSQclf/MMlPPelRM93YnEWK
Tr1DLYjT++o6znLByay1JwdGWNE2Q6jUt2giSP3OpmauyTTfKLhtZoCWBSmcVgr96KKJXuoRqY+R
HT/1Qa9aT8FYobXcHJlRhGlUQbpM6dc8IcGDpJ5dERTc+QIyzPz7zG9nVOe0jlDSkeODSiD4qxbH
f6tUiicpxInJwnfXGayueB/BPdudohiMy2wT8Fl7Mionrs/RSLubMXK8215uQBbYNsUI7e4efLaj
bZWotdzAqj8ir+dSS+M7X8kjTAkd/mlUQ70XK3fYhkqEHY/rKVESYNQyAfE3qOR/ecqXgX9JSzFq
QPLjdIPPRe9TRek7FaWFlHbkNhqM3+HkXoXHKFDfD7G0cGZ3+O9zcw1g41ERSKnsJS8BtYNXgoEt
XD7/AzwJ3Z+WYyhqjAGOgUrGbJ8iZ0w9Rux8pnQN2pTp2YMXPZVSpAsC2m0JhdgfaSUEj7GrwpbO
7gOihYOIoKBelyIRnCaoGUD50nLJaAaXg54Lxl1oUJK9H6ZoHMlq4cVyItEhDI5kqPUBI8pVFjTK
kzb3JTNR3LbanwWqXcEP2orlNUnkQxKOx3IEJ2teyO2b9YCYTEdtgMpUqV4mHrHG4hwZMIC7385b
U6e7s+8s7FKqpoDONBUscfF/8An1BDe992uPd9+l3dupCaWH9AFFGi+Safzb2y+/hvZw8Bo40qPz
YV2nWnPxTSDuhZ/Mgd8unBSsnv2c5CfIKQyRVISKMjD2IqpoUGgTzc+B+N0zXwWv4so3+3m4armn
nNexwjRmVyB1ciUvtWa6+NibcaAvIEV2+sHuRkf4ZNew7uZOeGcj0CVBZpnQdWeYGHEJ28tj8+vr
29GiUZxRAYrkvto96fu7z86FsrQUnxVb8WXw79Mz4LcwN989fUHHF5Ilp1H5ddW8I/BsU87tzeYJ
7p8jGkk73ePJa/rNv4KkHIPGE4AIIml0TlcUgOlZ9eU0Jq3TYDvCCx1IgqoY7NZhrmj/zLGi0gbP
5FxcI14ngDVWlGq2D0RvcP9nI75VfwfkuqYgqjT68WimShRNXwOx2TsGjLSx/hEo8niz4bPizN1n
FyBt2WXM52oiOztpmL8mHOXcviM6ACy8Dly/6pH31udtUwrPC3V98aCOzxV8IambalBrVFOwoh+5
71luEkV9slU5GOl7guH5mt2qTe/rAY/5oRVf93OtuaSzasEMwYT4AmGoAvQ1sBiTelPOLp/2Hl3J
l/7L/qIOXdJEl/7yMir1WBlNBbn3GYHacXup9rmxDzGqpIp6/wa1tEzSZW2IWu2bD+7mrcj/B7bl
2iHyPGduYZViX4CjKMEfJ/afCmP5m7P/8YUyuGnANaTx1jKm8WSXKVwPRXwWYvJaex70djPeYFhH
uZRZZeB+G1bTfL4MnrUtg9uzpDQojoK2epmy555G31ZpyPk41Qba6aKz9sg4CSTP7kFYG7nZAzAY
7vslHJp1N4GJcJCBQ2DwW7SKID+4EuD8RMnhAyChzOnfWOPOAG58MzOppt4yXd0gWPiaDuowrrmu
60yhK1aQsV422ZECoZpJWMmu/w7papWzB0GJUZ40r420i7ogsIYFwbrbBBbfpjzvjXnTnF0vjUQq
Em0Cpfnnpff+cxkoBh3HJeBDfmih4hSMq6YOsnj5UhPIHoiGkSGWwKSbWz0xVC3t3ln0kqn/ATes
8xRvt4HVB/ctVIIZtkbCypSQ1VNY6gwKdxH29B65fYWCiqZVyS+t/TpI67aEJDu5qhyc/xxE/uUr
qJGKijVzXKYwhHvdQSdtYYsSg+oIWYJrJnN5KpyAzsewc35SQHMIbATz9k1UQtaJePNjH8DN9vwp
ERrWraVL2GowCpdTKjyaSM3OuN5evyzco1K8YbKhLTEjDtuNExY20I3Tz/dtYvUV/mMMFuReMNoF
AZ0i8rj7A30BGh6eVKa8MbJv00jU6T6PqMDUUKDgmTZ6dN6kjuqhPzN4ZxNMX7HW3cuVCP9+3LyH
sUr3n819wmIAYYkpP34P7uT77Ds9hUCFWtdyO+PyatW+qzsd6feD+hJRqAuvgLfP0nrwqUIzj80t
JZ/03yIUXw7wIjQSBrmAzj3WD2UO++sE06j7jeGjGIGdeVgErTmkNO/3AvSSxdAAbck0+TTA9A9h
c/wWCLQs34pAnZx1o+NTb4GJjgbHueWIS8GngjoMoBuo8OOHwFNxKtTLENRjuyJ6/iGZ0+YQs87r
76Nsac7RyJ2srFHDKjSviteFBZm5A4I3riMDKN8nYZC5DfEN2P/U+uQYj00oathbcGhQXIYhefpa
CR64UxYUh5MiyqrC1Fs0fwgvwTpHpm11z8u2DQsdGOXCN9pTvFbgDmq7vQlGBGZFrotd/1fpdsfJ
wdMel5FJTBTdzbsFJivKeySLCkuZmcYs4UxZoajaUYUykmnHdv4XOqemxF5orQcdU9feBYLaO9Mr
uDVAHYQ4cusddFnD1U9KhZjbReAPq5d4uiv0+oUw6Rocm6jDe/Qntk+yn7hPLljfyXNPao3qGJT9
IGJfBnHfJQtEC5GHUUm9e2s1QBOCwePg63fnm9Mj2RKNFbWRnaN6slP2k1EkWdHnclDXmScV8o00
8Zifki12t8f9ffSaYij/lEBAAlAN4ECpnSGjuaoZZzz2zp7sqKj7R1iOkMr1oNCPJ3nd+AdxiYcb
66aHnLs6/35VobwilwgVJSHXYSOiwLZ9sRBGcboVpZO8julhqnMf6lKvSyKH8PeqFFhcbDooPJd6
ORolt0YAoBSdxzDWqSM1oG8/6cbfu9SVgc+MMCTbt04j/xHqYooyROy8RCGSG1pSJ7IT6OD8GFZe
rdbrF/sHUCckOf4qwTPpl5rhStqNCi1DKwK/S1IYA7tgRIQDnyPlhtcDkrEM73AtP4uQWBQWnL6P
Akxyr18j2LMIVz/uS/SUzGAHsB++V1jeRGhbqBEjdVNkc52jSPKVK1DZFcwzXwD5yeUQRXbMAqPA
Adm6/ZGYYwqDiWl2g3B/2CAch0Ncj9/5TTJmqRWi9Qmotyu6WleLFKUlnuXZY7NWQ/ZlNpozftGr
MqTDWfMlSAPDukJnd7YneZlQYGCqQ9/NWI6jR3fCg24/xNWm+116YSfrodg6/h2jG/cQh50Pglai
mfJiwySXtauDMYfxXzBs4NX2JRjQACLkP8PbKcYrUa6r/1yKReoRxem30cx/veGFHfGdtv4ORj6r
jfIWEoFnFd4VFQ73m7ZR7YOHUgkTIrw5I0whsoAXq1iRrDTstHk2tQmzFjMirYqIfV+E6/g81f8K
cdijMiRaNuxNCsbdM8Cth0mFE3upvSTox+rHZXIXbsjXlmGkl4iD5Q53F3uaOboZJREgY/xcLf+f
NL15DaXUpIcenxRJESBg6oLapY8sJnp6DEGlQq+RIK1LIoNukhIuusLjkCArIkwgG7GSCyEM7q2R
B/eOMWIwz+eG9OKRyge6iXrt725iQixCQu2VAHEkAF0ej/EsUB5It5KKXzo8J+B4LZMj6bSHR2Gw
+eaFa+gPt5JiGL4AS4ZPU7gzbwSzvzjKdLss7WAFIZYsYxMFWSQ6Nt1OWYQ2QC7vEirxdta4EOsS
a/3BIOEiqkwtNzSje2P9ACAA+QjkwnKm5+xWvAOBzGTOxVyypc72AipayiugY5dlwi7MiD6DJp2h
zghb854c4ljJFrA3+kH9hNJLtnrDIcCdTe1srWRkQKrg0RibbuNR8zuRqYB16J1qEhNgN9y6ZAwI
XktM6NyxjTZntryAJSr6Vm1snuiTgSwwjpZ2857OEOwSJVIZADogm9H9WWWRsJ0o4RuRrB4pchce
tYh5a3L4ZMiYcKUjycqgCKWIUjsyMrm4RzxNFwIMjiJJnp4aAK6paq6P7eI/vAcx0pciBdVymjXv
85opZj2mDPYpyiRqN3YNBCvtUCvZoG6EGEZ6ugASlay9upyfxbDJTjSgUBELdq93zOQ1kxo1OQWB
Zj0/yHvy3yBbL6pdzBtCqYTHFXddl8UDQnX6wtN2tuCEo2+l8GSpP1KaEgb+vY7A0JzvHEojcLpX
TFPHoJwzNCM/l0panX1ZPYhjmC+HWFGt7AjfdsALO3EYE3Gv82JT1Dq6daQ0O+JJ8xnCXDbzUgbi
d/Cv3+WQM2vqQ3X08YCo3wuT9QNLYNm1naihBgrQgs6NcJY7dv4dagDPVesNr7o2zV7oWt5AIHec
mmVmLHIi12PiVeEjVq/FK9SPj1qZn5vrFhkkaXkFNY7NhZSKWoYX8NrXlDofDopIvM7Pl6MC1LsZ
9r1yMMMCb7AJOv0IjjTZ4zvUZUJ4oGwa2tsfuEWYbmFDW8/FNAWcJ1+bSXMYdCuXLUmcKk7q7XUL
TJ7kvlHR16SPCVGBJxpkzTMJa4svQE0DFxKHPEJlS1eAJq83P4+G1Fq99lFJMTH/AJ72djzJqcVo
ndAF2cnetEVZ/xbsUCI3uLxy1RZNTVSSvF7BpytCYsRmo8EuGoHyc//748u8JbwV8/atKuR/79YT
KSkDKaE1gxZyo9dBSap2+3D0A0/vmzkq9xzmoHU9U35IJU46HKIeyM66e59ax6Jjyw4hN4ApwuT7
HUw+H8XLrBTyf9ADnSuJmRfWxG4WxafhrRvDIYojcMcTQW+umBcMiUMyBJwuXq/Ze5718+aiQsEr
FCHpK9Crd6BNTy8j1CcNWI07R5RV7/LDa019N3lRetDzza9Ra6kQNRg1tm7ZapZlEwlJQvNpB7Bp
N3Ya/LysS1JRBSV4pJjssNKXdxFlDngGaO0N6VMvwfAQ9O3FgZ2dRKtyBV21Pd98H+khHbg46TUu
t23y2i/68kW3ld89TYYe7NKK6NkxuZhqyzE2Wd8Q/9AYXZg5HhyHPhcWvrK85lzr6o9OO0X6tsjS
zBg+qHuxWw0giwVhzPYVZbXfwwrWKdb4rA1Cvv8pfms4+dhjH0bW1yfFm+2CVUyDgFC5cYudOlTH
QQMe2VhLV4yBczfku26fe9ou9sc5FhZ8PopynGYxwNSKsYaFVLMrrOf1aSDevfVz22hQSRdfwC8j
AjMSL59BgOQVqfYsCM28h7pXnWVNNZLj5c7RynNb1laYTz8awm3AGKOEgZIt2a1E5IS0AX7Wbp2s
Ezzsk6hftV1KAKifVSKShayL78O/8x3f+FhfsA2eJoxxw5EpQY7Tt5iHip6VevVc51vubEim5GGD
rrrcmAw7WjvXtUeKBJdoPJyn/aZy8/a1paPqdGmsscaTuEu38swHuFXWVmoCNpRUyBP3E7Mmd80W
1WQVNcws9peKlX7Qlwe4B01KYUo7CBzQ+5pSMRecgOI/CFAnICDh4o3RZQW0mdmPYZWMZNYty8zV
miC8++XnraJ0uFblyCYxsVyNO9oIoX36QS3WoKaTLWHUQqud15dnpXlhSNtnQIPc1Wqzhb9Pb2CK
dTPge9AsfB40fPlzrW6c66DSZuSDfGtrfDo2KS71XmrgyMRirT8kyoARrfBMd1uDsQhh2CvSdkn4
HSN6bNTYZOSFLQmJnhY5qIJHsymx19ZGH6vB/260BGUrYfgUNDdYlLu20opD6ISKYE8Zarv4yRUq
rZQ8jALT9xw18QCMM3/VtiI4iuXkIbvExgMLyOoClYGDFrY4dw8Gq5Yf52K7Q0OlvJ4RwjbtK9SH
ZYZgf8bs5pw8VtxcpSJ6JMxCXWeGb5tdT2f5M4EvCW94StXa1rfcSs3katPavWRLbS23kwk5IE4f
fVhiyi6JY8KsbjQiwPXscKrvQnGY5SWOoUAf4mG0bDWm1rT5dyPgeifLIgQW9VoPwOFLbd/n6ftp
r48xQNAYjJQvA8NZoWeR5mySCCRvOd/0uJ/akt5vj/eQOMLyZREU9XkpUYyKcCOYyjOhMHYIfKrX
xu0svY63dMR0GESXztpB1m43uhyzB0z9tyhqs77ZubXt6bL/ts5pF+wI8xsB0dsCqfImQyTdaqoA
2fVdS1JQ+lRAbDh3NHE4AajT5+7A1JYhgtiaPFaPSCpdDcoFMUzByMRDNj60qI1RAInWkuK8rEN3
7YUCTlh+l9qUM/a1g9j5OC1RhBPUEshk+An+48rY6zoUoPSty7UepJRJ0z91IHVf/1Lw/eI/NhkY
Mk3kdg1X/kk2RgMr2IRCxTc9JETjQZfTk63tMDeWKmF2Hr8dsDkDcUKTZsXBeCjSefX1MG053AO1
jMgQwURViQllje8hYvxIvH6eNVSERYymDbGJXKS6Qyj0Rkk8bfTS/kMaQRYVILS/sypXQ41KaLd4
EF3Cu9m56vTmpbxF36q73WpPX7zK9d3XOPNlcw/fQR+s0gl4pAfVgspr91vzwsdheuuR3C0keboU
CbS3bSbBrqRUCcHm9oW0V6/GDJ6KiKDjeOtpa7DXhe7fgSusS75XFUHsQEZuU4AWjymO2NTXNNxb
C2mKhGqHxP8QfB+g4mDrR5C1PA3hllqxRi8+J0if0mPfiVYR6peMBe1rCNsNZmha3Z0V1z7BYQOc
cTIzF1gUy8oISvCFzfmkYtmQYKOIqLZvF9vhoLMvI36R7T9K7t5kDYhvVzPUUbr+JcBYOfiYcmIp
7C2KMQ+1d25zm861bSmZCtosrybV52RkPvTp3TZ5ldGdYT0aV5pCErZXMDC3zlMz2IVVlQmfTevY
7w3eET6GRhua3vLSUgt0JkoAn9lTGvKsNtulViMm+ZzYCc25MLnbqhEPXEN/CfkJQH0mNFezeADJ
doYBqx0kWCV9E2E8QHY2vh6kPiiecF+Z6nLb5YOv9u3HcrDJ1Kc4GqzDTUIo4PXe0oszHiKCjoGY
ZNsMfknrpBekErvOdS/EXLe4o0iAge7U4NxT+4nrv7sfdLCku/GebeV7wQzadW5v5iaMtM/iyCxh
WKgJYdSPV0JwZOUzhU7PLf18JbAsnFy7WyYfcdcV1qpIyEmJp4D+cUmY9twckohfRXal4ZTPWN+9
cpHvLjG/r9OePKLVTSdB0IMqSEfeUIiNsFNnE0A3reqPsOH5Evh8L0p9ubY2W6PDEwUOtnLR1Oce
qxhftr7+pL/sQIN5UC1wEqv7BOmU8PiKrBFYQCi2kqU903AJN9A85VKRN4eSiifnNeQCwvTDIUGN
+opB3brrkjvOg5bBllGEsp9KRU93rSRqOspNRxr4xQrVdbt6+VS4p3k+BwIeFfvSpZTj6Ss0XTzn
KHDVmLfnDt2b/jijyVLB2z8HDJUyoy6339GjGDvkWjHGvkOMvXHlccllojBK/aQku8zUJB8cu9DT
vqUv5yN5J5rp71OShET9ppFmtnL4MNDA9+0JrnXiTUw4YsyupzM05oiTifzW9KSwgMU4O8qysw4r
3++AsElQNHJNfZ9zBAYkZgHafDqtYd0jl5EwCeMG2oWqzm8DrFWDPpwNqnRtGiDOO8QN60iwmT+l
FBvXJ8Farls0wUkSR9D0c5LeoFegREfIZCy93MolIZLDeYsFwm+PbvMr/jadkCPTGTtYmU3/rRAH
VpVr39Aag6enjyFiPRM1DjBbbqcE54tLntbbDMjaTk85Ta4GzhCecuAGDyzUHefIKQWwtqFgKZy1
+IFYukhVIcJAoFgdJV15zN7Ar73JAbaS4HlEEXpGuKUHr07szfDTkaOZvwBTMOnWWzUkTnw66onX
M4qyvJBTwQXuQfLcE230qQiYF40PQ/OU1phKKihgv29iv3Qlik25HQteAVHHqqQgBAfYwVGyK3BR
xkKpID/MXgzlx+9oKX5Z/59EShvFUzXvfLihaVTI+qQ91cdFG2yeTUA1Ej6nnUARRyJuywQFYbso
02bQYjERgtqXBrCypN/osPmSlRDDwqw5AWpa9pyjXJF4sLlYeN45YBNwinz6V1nQVk07aqyqTE3o
jyk2mSGAzrIFMDuDflAowj4AFHEqFTxci+lD6i+G0ThwYDMzrgSHafgZRBAVqKF2knEIecSMrUaW
kwyUKhiVrKj34AZKhp0H1pfP02YesDbPFbGPMREZWDp76U3WR2LK+ILX+82555G55DzHNlCmSV0m
iHZfixV/4blDI8kaZn/kjETOFHvnJQob3b09VsjRdDRYHPZop9PM8YsX8OElSO6paWzQM9vIxEHX
tRYFoiLaO1iTdvmLhVOq3Ms8tet8DX+ddcssrqr7HEYx1PSuY/r8t7ZiCLn+K3YQplxfktIpzOGF
Mzo29Nidz6HjwB1kueyOAZ/tT2oybE/V/dbcMTa7CsKWmJACiEmDI9bZE3ANK4pSVF8qbICnYsM1
QB9ao1n9ysC8fUUONcrry8xrnY+iTl8szbrQWXrhQj5RpqrjdH1nOyKj77Ngvyk/5jgoMZdQlGe2
WsIr7KNg79DqiAVCBpfGrvEHFyflN6pksKTjPmBjp0zFtSCkgeTSVkmXeJ2ngWYTdHzTOO4gzJUF
vCiCuuZRcxC5BOgTtz2+4VjnB6r2ZXLB1Rk4kBcvecZoGoXHqQ7ZDx3WMW7OPvL/KQc9QyIKKlS/
W6C40GjkHe5fnLxfLkv8sFFcOoU36to6452toUFRoqA4c7A1bUPrpLAbTyVP0qtvsD48v9zl0nbm
ZNTs+KiWFhVXgcBJ6TLyxOVxZC89OZbZBlhAaaV4XKtRG8GMqnAWoP7k5mj8c1YRR8GgSVspJWVj
jlNz4pQq2nGXk/7/Nn23oXd7RhEXe1tnZ2Nf4AS2Ka8pakc2fIDePqsNuPCIMKWJNCPwcD0Lqg8S
eWzs/uL/ArPn4AnYLi5Mt9q5XOqKkTLRJ94YGjBTcJAnmO4H04d0s+0stPxqZ/IDAAQUxDuHf7dN
BH73nGDihYnL+upnOkcYQjBT39SS1FY5cnzhOZEN3V9vQWOFDgCY7eG8DUXes6Sd9NOOxyTD5Ztj
FRuHet43nqOc1D7Ghadge1SpPekXeYoV4iTQZzwNbHUsYbjjm8Un5fK9m/vtQqO8FDTED9wWUWYB
LDk5IGoiYv2+XDeKQ4261ctlt+ZSDrYaadM9mdpZrBaW1lPA8eRMtvLkdYsJ8M9gQmZPb50wUXWr
ffrDarjjK/qN00n/nDX1x8DTtJoORs6xQ+G/qyqiEjqRVSwYaf/KjQp9EFSm4zdq977+Xdb/EmL0
vNRxJqy+1grqhw+MYic+OIImpWxWhWrwggJEh1Hcrt9Akg/2sqTrtWj06YiTxjzUn+E7IbF7/x0I
vmpObsx/RQZfwQrgatRlCirFCkpy0/3gj6k6R74D0z7tai2bm4wEvmbcNYD941K7PduiriLGjAU1
cUvtT/CmWtUkjX81qP1ovtrK6CBjmoha/uWK2KDkBHNaq3rVyMrANFRLUQC1g4LtyZHNMgpOCcky
t5o0ynV+9/qhl27limS+6VSE3kvvSmVzFvnuzLHw4k9jLSfur7B+zN57aNw5b/gXiaHzxnsjIxUd
T44PWEHywSWBn71zyjUSORrtyq0i/+65mjJ7RS+OTTeknGoCypeClLBZl4U+p0Q6pTKTexjdnTgn
auywX81u1MYI9NQlFkn+dUX50C9OI9qtGmGLgMBRfoXVNp3UWOH7zepzgLDMBf3amH7FFuVoa9rO
abMqKmufdJQMT7WQ90BFnrYG76XOXk2NthLrcUxBKFR9ZzDqX+MuyLppjV4marRumF+qqXlNUoc9
nesd9IWxbY0F7y2dXkkYXJYhWVUHeekxwwXllQkruXZzDOVZ49W0wqBA9QNEmVrr2e3NTa0Z2AQl
kngh3yJjooIuO2OYvjJiJdl0g2QnzOLOT4CMx3/420eY9StTCTRQnP7DJ+tibXcpefVezBUeKMr4
3Z1ZI9tLzKXkVO/mVCcxnkfyeIpbmOkWvhaF09dDkkZGeIrXPZDl5nkRzM/omFbq+cxNKLHbg2Fk
avDnPTX3Ag1JvSERKGaDHkzN48+6DzTtY+udpDyHkXLG4UGebVlCUauU5ivT3/X3Jac3Tw8QLH1H
ArSdvPNUd+pRv8iL/8w+aWUoKlz7q1/ZO3OyJswhFthElCjYn+/q1sqkAQcCL0vW76QGmV7LC1pt
8gk8FSDRatwyWvAlRpwvFioPHFYKRzJawNxI25XtfHA/fszTdmAtlBzEpiyj5qP1Ra9ig3Nr3hA9
CxiyBObvCj2L2p7HPeAoYE9AMP5ZJX7Rv8RSaz1uC/0y20Zu3j+KALzfICU9m319L+VejneiZhZo
iaNY+BJOiZG3Fb+H5Mw6Q2w64ZY/MD4wWEZnHnclPyV9xy4Ur5fO7alY2JUXKTkZ2RXtkZ6VkCqg
bOPokv8uOmA3lgOGGTS50xsNvIKxuA5pWVTD8RgDVI4hnURgCU4M4jl/DDIwDqEtBfuS9Pv1D1of
sWWmFyT8mcTQTqVBfItsMEpZ5DwZNbTKh5vMj8SWo6mpCBupk74AVhSzwclOWQ9EsN2D2pRAPBjE
+/fSgW9U3nz36kuh6yrbgoMKocka6D5otCWZEIsuIR9xcflKgvz+wLqAtDCHNH6ZaFaKhRs9VoAP
h2VlFFqKYeRRoHJqJTC+JhS2AAxmCiGoC7Ya880rCKcPkRkF7Q6Rd149DTgifFRbGFmagnXlu+9E
4FXek9sMbMmctTOOI+Hynz3vvhFDbP3p4YTK185gnzrmuzHi8x3RAGtQccA9fD+oQt+TEGXZ4iWV
CeDTLpZ2xCAv68eLwKtn4kZmgLpVhCJDcv4VlQ6hyyxDIhLlCetkdiFrjZv6LGNBzIBM7e5JINih
pngTy7mOoObHOlSmqDY+Du9M2UaqDNEQJsoXIg02yG/Gu486NjJVDn2Vl9kl5I+A6spgULekWAEd
6QN53Px9d1LHA9+JwD3/4EnKMbFnwHit63joGq+yG15ic6hp4/9XZJKj/VTlv+zAbqgTDU2Gl1ay
A6Gk8q1eCWSTPfCy4g02gSXPwzL5B3zimsycGs7b4I/fLbVV9doewpviaa14LmE5A1vVeVKF2k+n
gh1IuFJbblW3ySpIW1j16SguOTXaTQAK2nPtOJZACccgnIlW3xglgWRo+2Spd318JIhiu174WN51
FsHKEKCZEzu+17ARr1a0hOHsSSy2k8QM8jqk3EtlKtI2p+ipqQVyG0vWtv9CKWoZ/A4h7vp6joih
v7gBqb7LJBaC6BEXeCcdFhVHGZCge+MrD0okUXyEgQ5+0coaVC3oOYTIaSneyVwwGQG9CHyhv5LC
X/6m0P0OssYkIlzym1mQTNIVP1g+QaBl/DsOK7m5qMdpyOtxae29zaZVSMtaq7EtU5inpm9tJmr2
44de9vcG8j2f78TYFefxQ9T1tcXQ8akjO4+rWmGGF6F8Km87NfxtHy9cm53Wy7kxQSgnWYfFsoCQ
rqnNdlD3iebNbDhGugw1ft1HMQ23TGTU5r1I4Poe73GYEa+F51hXoj0oGFx13QRnnlXdCP307EmB
hxLC9BhJO3JEaRk4M6Lx7HGzOu+2rEdthx9Ztl+VQIceSljgrFw1ax1MXIeJcdY0+gWSILRWPGM9
kZLDSbvnxidpSI0ZRIKbyxNwQssDoDMkgXT8GT1Q7wzw/HL+C8mLJpbyDX88EYn7xROPR3W6V0tA
+OWWRsN+ycVhNZUDG6dHBH9HM5lWgO6AjnzJ+EPwPHD0//1gfGWfHogRtOWhQ78cABiCC+yZVEwI
GPp9XSutbY9EyRkySo7BlMOUN0v/a5fNdo8bkIflf+hl4ctCwauK39dyMyvMlUshxpZVph3NViI0
qOHAkiR2UMxfGx6w8WjAaip82d7ID1PUuOqwtrHvJbdzoCqFcuBAD+s/jlp7IwKImMZegh4fS+Hw
gumc6iTWBWrPo5AMAB/33dcowHVOquwdGOmRufAogI37IPGMDx3Rb1BRA08xDdRii62D0klxN9mS
Yflx8zWyE3ShtbvVgads8zKinJlcCnCoZ4uxc8f8jKYk3K12g0O01U8XudXThtYVGSF9iX7X9+pK
j7lBlJzKiz+Z9A3nZNgwJvEJsxc8JmUD3IipGYJ6nQmcVbj8Yxd3ZtRkm5xos2EhGdrWHAizv/XJ
3QJUlyFu/RSVyN9LOH4iLaH1HJwIQjWxyQVAYtMDvfA/aeY06DNHoZSK/TTN8q9+t7w0jJn8chSe
/4yTrBBr/6V6G5uW2/EBNjBRWgdJGAw8n/CTGb3wRgp2gJYS+cFLiyi/VOEyilMwGzf7W3sxypWW
4viJMs22yyhMfc9Puh4mRSq7nM84Wih2a6K2wSs5TavGUcbwf2ooYy3+bCF0Y993ir3D+g1TJgjm
tmKlGYLYbb2gt8U7A58EM5M4AorCe5VCRU7DMrjBQhXBvqLlGqSmgih4xHWx6EVFK05QLvaRdaVO
0VRrvzinQQcoClyyWXWIc0Qnjdgd9JjN1EK/x+/BxZdfMk8azPbMUK9n7JNgMKhP2NZ4QgO30WXH
rbmVclVp1wUReUYafaqp2vVpIyueaLHqVKBiZ1WnE+1ddc1x4fxYpwwYwZCKMbmzn9/PfmvGJ4kh
/AIESeveN6cYTu4pYTtDxPpR/JtkPctQRl+dPS1QW0Ye0YbZj91evJIjKN3VLxm1NnJvlvAPwA1z
MlXia3Xl37nwP6WZNgoTUnu3QhgROpkWqwx0zswk4Bn5FDHNqsVJqzHn2nr5G1cryxEvwkpI60/j
4Sm3nhnRoMPh2vn/a46HetF5s/O9ME6B9qSR9uhMXmXHWb36sZW3enr7yxOWlHhdA5eap7prP4yv
gI19SMd3AN4SB2+nXwAbYp2CDQU5iqdxffqgVUbrLMZJwcJK9I8h3rfbICnPmwlTJJ46ZwMdBQqr
QeWOAKIQW+24DVneM7+xMFyDNNlwDFilJ62Ck+RwMaKwuvHiotrH6T8pikujYE1cUMdPUx06QNkh
wyo4Bk5axK9iGfMRjhkcxv8T6CMoZpzaPwnq1ulFjNZeP9OPjISvEJDA48EfSAqa2bzP4dbAaJfF
OCvixM9GI8Za1/D2O+lpW9TdUlRM92BlLh1WH2qoq9hiserRnCsof7FxW56LvK7m/ips1CFyM4eM
czlXS8Nqbn3T80oXiUOc+wyRfJrR3KBca+tLbYMssjtIzLZNZ/N32Kmk6JxbD+mAYS+J5PEDXZRI
Aiv2BBDGQH1grEGtZYO7NtCd7dg+oQZrxeSB9K2kNo1ktI5R+UkOm2BOtRUNoQh7y9T2UOhB4VEa
xc9kyvBY6EfRQ8ZHcNrqw6ouK+aYTLY1BbuuH8cxvu1qpbGj0/ZeAM43IP8o0lZcbCpAG5bK9lBW
RZeahHd7sd64m+1bGGt4bKkLDMAOH3YyHeQEcELVK5JFPFwgkzvRo/ZfJvufvQSXnIZmSWZv/mpV
iIyrjZm73/y8ErgeuwMHRQcKUO2QhWIc46LkdFcOBOIMX9K4ZRBgjLdk9ooojcm78lbIxPz/DH7T
8oQL/iv45+Y5G1I9j4nOupINK5aL7CIQW04hzhhuriI+wESyo3WQ27QNupV2aedMrV3wgpIan3hT
QrY4gv7dWKk/pixspPhryjaFDG/xNPXYwFb9t+fdzZqtiQrl0R3L6+Fh8tUKJRA6c0NaYAENkisF
tUuhlsylACP4kjGlB63TXovrtvGg4mXvQTkFZ+gjkp77woTmNFkazjFGtd1C7IIzpQLs5fDiMuod
ThaAApNxvtgR4irEDfNb9tsYrKYTI5vsads/rperXBFLEuGCPuoaRIVEO1ugdSi6UeFMOqfq6Eb3
fsbcsRN2jZnEQPOSkJchs7iBkibePPsEZ3Fn7SwJtIIjEco0IPzIf/ax38OU0kWDoAOpv07bOWkc
kc0Y2l9OlmrndjL5Ln4FfDDnEq8S7Bgc+zJsNKwiIvu7w1PXASzN4aebUZdcVEuEUAgaaga4ztF+
Fa9W8CKhJTRVibtYCafbBs7NVTdpQ6lEo8lSAzRL32vUUxt2q1XdhPPryzMLXob845KFc3F45C4J
4LZd0wa5Y9btsNYNpaePXnpESqL2dlz7KTRraK/2V7i47S/1VRYNcHiqfEpr8VeGs/43XQaOo+ky
/Zftpphcm2dodYSo/wcsu+qUiPGrCHBVcaWERQL049IsGmqkcLWKfmp7gRXRwsqvDOo2oh6qRKtZ
t9c/hstXRLtL9KyRhIkRza6VsRnr2vqqIgqN2389UlEHU6T9a3x7nzWDoFbpgu0ADS3LsXj3LRvF
4HrBRQoxK479ifz4o+4reKQmWA/SKz7yd+s1oKUBtIyBFl7LBtjR/zmBgjhwpEUp/gPUJuh+2lc7
ZfMV6wC+wN5PBMEDmzoQkvyPUBRUI++OQVrRZ/loCQ2RMINtnowf4OYQr2cQ8J9vATqrMM1rRZjH
xh4vwDs/hHlDaowtfMMQVMFAumjQ4MnWkXSL+XVdNjMCiEFK6PSz/EIqqBDYkhDXXZ9DlhikvfGk
hj7kboKPB2kJsZZi++YDjhaxZ7092L8Ch7RtVIF88K+SBnhqiYmuHCuhI71xkXeqZAtfFmFZSpXp
Si1UcZpl9W2rEOpTEEf/j2c465C+eZpwuVa6zlIlhiHD00XSKwfrD/3b/Sw8urPqQFo02hLdrSEd
IqpGzsca7YtiXKpzgpLQhoY3nMhrroKA+tIz0tLX131cBFs1X6lyL9/3NEU9eUPROD8zL20+301z
Y4CqDWvT0rf/rS+M5781r2KTasZPDWwAi0stj71egbbXzR08cumAWMozt5aS3wwxFP0mOV/dvTFM
sXlGNeKAmd0dhKfdKctka5lrvt0jeJ7VR9hIs3rLw+rZez9cOP4uKMscM2lG88TbUABhkIeZh5Pk
B5eX1BkiPTRS9PaLE4bSRupLhJgVqx9dk5aqizWpKnfIpRJrsmZ3J0wSH6s0XUNVeqxA2Xd7SFzX
RQfadavEA9nJ7mp509ADApt/xtmj7JNYOoWZXN7wDQt6QDEM6GRbGqATfzRd1jyfXTBoTyErkKwv
2Bh+XmUtATcxcTQBZ3NbYbn4k4DSlKvzY/5N7C4T7aJSCgJakAgjxjDEmDRMLe5hWlEgnD9vjb2U
5iwreYJBtzcUCzDjd2+Hdvq7baHZvMFmk+yOuXqzEhQy+5f7roCbrBZtSDDGYHcILgX/EzXcW7sZ
y+P2+F4AeYceT4gU4vuZO9wLEYrIZaljZWMWlGq70NCK/oa0E/9JPMKkC91meaqoOZEKonERRNUJ
CnKDz60ukSFOk+8DQxhe1iaLphzIlx7oJ+mm84U7Qq/yyHCqUZEskT/nxZhUzF4HyKgFv68T2j3x
90CziqH/jHSZf1nNUHMnBlIwro9oiJWZvr9Fa1C9d8wHs+GLbyYzajvB53DusX/7FnETy09vbU+s
hokIK7W3LZtRhfPu2LO3KtSSfin7y9xPPvFuWiNmFJMJ/hlfWzKorB0mK9gI86Jax9ZpupP3Rl7w
POCnrA8s3LGODK6lGzbGBE19MD281fWP0fIBATdeFFAhJEmFxTLw1GL7mLUcmzM+qbxnNSDBs58M
vwPxSyJjw5BH54MWKPnc6IJnVl5mX+Hw2xp9fxVcx52s9jBKq+QZAe59vq3qjYnx97B3YBBo5zQ5
QYg5e8IoynjRrRLG18gUSvBIwaV6It5Em212DyzZta1tUv7tYH+YvDog+K7sjzqwqJTl3aw0gZbW
ybaejs6m7zvK/oshnbIsvNvKSF15iVF3zK6y+wRRaNFMaSvlajEp6i3s5qOqiALCyc1wBqE6WFmL
St1hKdKPjJCId9yWq7x2mpjna/Ut69CIsYkrsTiPMSeuddb+tjzv38Z76au3Gi3YHfKW6e1QOv1r
ykZKjPEMm7FN+QL6oZC8SGNWHOYnmrugtDNGTEl5K3HfyYzZA79skZre8ykGJoGbKUr9+mi+krkj
2KhcZ1956vALX4FS2T2DUFSQEJtpOJqIfYTFtwMW2E0H3N7GkrHJR1xsAMJw+X01Mx91mgOAwfCy
3YgfgqZD4Aj4OMrRemmUO8q5aCJIadas2KGJR1aKuuFJovhmg8bKF6bg/4KFRCaYFrzRgTTXiJcU
ueQiAIZxe1Z/xqKAtgSI7rr8Bu1XrqVtp+m8nj0ezxafDBGsNyZY+ZFwa95IQzHBtF5SstmQpyQG
XtYi51GsWZPtF/kPe1OH5Ec8O93njmI0UHiqM7cQaJPGSkkZJDr+kutA2bJx4cogRLhYGxKTo58X
SeIzqUOLdQkhM7kfriOkXS08+4B7IrRWhfQVwV9Fc3VTkwlWTHleIQ1ZdZe/6gCGWvirfcfS54EQ
9hPL3/RPZOfTgRDgP7m22ANOA2Dq8LE/oYgj8+Jkbu6GamUMKr8zFEd/PpI6OA0M5HWr7jdSBV9Y
1H/BLjC5oDj1czLpl2k8mQjE3Gg3FAA+7glZ1D+oKqgx9bSK0bfa7C59QG6QVNEN1KWx8GlrnMtk
PgI7DQj7Lz0xE7LuwItnza3aFKeUIBwZ4O5C0eekzE57V3hAS50NroigqmWXey7AJ2F/rHDCO+2a
eVvYET8TntXxHzakOQc6ozbuV7zP1PF5EZ17ZB0pyHVftt1aEjrxF2Acp5OGIRk/oUwNQ3hnG0pl
8blgmHJL8E2pzLExPD4HQqUEGE3sYvGfNf3sxixg3dp/BDnXL4g3YeCN6AUS8Tz4BmN9CdDsDcVu
S6yasMuGKBgIzrF/aM5LqQZu/YEGuokBmV0vWUHqpk+zQdIpHReuPZkcINcWAAS7mRVUUSm1dXZX
FFDiFUVSmQ8i2cqvyus8y00fEHH6OLaUBAq4RwHJcCktjSuLp71fxNBWSunLeO/HDYhz/4LpO2FP
lUgvjmPUsqzASG1DI2O/FtZ48JrYRLRv3q5MdNohNGNt+ctxTG92zyfeQ07MFXgrDFuh0GNzl/yt
BklhENKyD6wSMLxjuR8zs0I1rdZCQGXoMq9pGJsTK0BIGFEsOQbg+HKU+eJef4YvoKDpRR6Vnft0
CMm9DOQuQ9fBU+bEPivroSN4q6jg3lnfXS5uBSQE7RAGxlUEPDrPDb3T+fzAa466MJhLnwu0/S6M
NVAHZwCvaxwd8O6EE3b7Rt8uSrP3OBTGapeI1xHhurnvua6lxYkpbh6HEs0PmVz1ndWMSEEZXjuZ
DnkTdCOaRBu77TgI8D4z9nv7FSDfM4xv5i4BZmao0+c5zPPbYKRZ2iniqFSz32yg3VSG6rhNrIQL
KpBVL2fO+fiUhofFq4oh4Vsanc5R1uZCGoTGUsyfmuSVa2RgmCu5o+DSjh9kgL8LvTxoWf5Vq8GS
TWZY7qTrewCfpw288la91eFvkwyn49Gg5uRGSmAGWuRzTewbSFqiOYiath4NRIXFd+/QjILV4Vua
pwhh1R0lneFNBQRecyNNRGl0SWP2wEvcGEpYa2h8lIHLcIV2zDbdzRUqBj5IW4V/c70o0vWbDCUg
+kydsFBuy+ERHeF7QYpmwJPcpatDFyukW9mYSvM8UnZJS/u41FnM3rqfDuhnipp60K7qXqyElgW8
hKBcSIpnc6NvjfEyn7W161A61CslTg+tq1XOl7WjmykCbXp+T5Z/9qdvQr34tun6Uss8/Df4R11Z
6FMxLkXBNikdII6kvUaonzgn2oDXXlacPU9GH4n6NjFjFRvpKI4D92KJSNZa1yJSWkpI1cRtf6M6
lsPLgI63X44+vBcDPWUARiSYX3qqISFCjhr9DenD0fkPIIHqyHrdZKejdV74sGxzFULN2lD37O+S
vxyQGdqG1CTX0d32VQ+wrxAjqGN3D7TG7c3uFy2JSvfaMQdF8oj2RRP2uI1KY6P/oFZqaUtyH7Lx
Nu0G/0RFRqKL2rdAsdlgY0lPhxufSE0vplo+QPG78jiojoG3gDUCmLmw/feEQCySkjVLSmhxVITJ
8R25+EVesWtaWpTKjRrbkwFjjJhesUKZoglTMf0l7OiAV1ol/EqN6S2GQPHidGQOCIij/9Dq0UyX
tLlbas9rKOJhw7cUmfO13fJl1XbNzX3yAOk4vmzOQ1ux645JzJtYsCUe5XsnNRH0LtLntqjhe7Vz
AQRqcd2szoAHoI+wyh/iJzWuPjwDCXfL6EYqkD4EzfFcIPMEtJhpbgc600seAql+4f6RnGUyZi8S
L3l0t7NDaDRE9L9sjT2TRc8pmffm5nris22FEqPYPEIVaLyozlFfynqZ55MNcVYPB74ZgmtIDb1m
sH4W6L65eOpYpIGePFaPV1MpkHwWwHxKg1HuyUZeR/lIs8GPodyVeIh4vUpuJcKxCmdCUi28Od6g
JGLCzqf4/+gk/6uyrjL+q2dhnMGePU0FrzUQ9mL8MawfP367ZvfUtOptPLKt1VBG2dSfLXEfLBlF
wUxyskW5fARj8saFbWdfsoUHn65E1SUz7YH4TTi6Gh1yfC0iBvYtOIiEk9ygDtoRtJ0m7wIOcZ+g
caVwP2qpG97gX9P5Fc6pc3rX96xPlEib4jmLbMmB5oZYPk/ofMp4UwxdyHQCLuG6jNJEfudB/hKW
gPI5B0s4TfSQNT+URA3Muffz2u52oJb7LS4wC4mYTLrgHU/cTyHNT9W3QYgGpgZNM4usPIkwDLCt
he0o/3T1VHomHZ/Qah0k1wkbUCNIQcAotdHv3Sf7W2cIo00blG7FoQiv8x5toWaZCjGZKLn5NmeM
CHMEfwUepaET7rPF450Sqa1oAoex8cY/LLZdpTsTGt1uB+v1EpiY0eNVxk2KP+nIWMQ9kWkKyQAC
vRwlX6EkrvyXaaOTpxXp7Duf2eVE4cMf+ZLS7nC+FzwZ6jNnaO0OG91pK0iTItabKiAlpVlrF5VJ
V6Kie9UiDtcvA4p7cwdhTdf/U2y5KE7zlGpp1wVmmAcMmn5Nugpha3zNNmK5b+BA2oz31mayre/m
uh+fhQOyi+OhQ52sUNsgAiqVMsR2tT2rr7Fo3AP5r9CraBiQZ6axFvMsV92ZOoT98zhyoPikkAYu
m6G/Fc08aYdVDmmjE0wqS2nHEulDNmTdPp/tQpPDYEFDT7PWQpDJmaD+Yto3HeAQJiZzlGT95t4s
lkqTB+VSUgL9GYJ3YkOI8wdmFrQd2u+15s+zsJW2gg22DRzvuQ47eu29aEhNNxJsWIYmKpj96nsO
rKAIYZzuBrhR48UlVWGVuqPwBTUFMnLdSAgpw3HcQTvhNgg3ueP7wzEKc5HA5p9r3ubypu3iqidF
oc9dIlmBvv7SqUidUq+PBpRcYQ/0dC+KxH9cTIWmxIZvo/pihIm9364ZyC1CH6Kz1QkfwDm4JBwa
T4x3OBsfgwAobQMu+8YW0Rswg8t/5pqtn2mBcpX5PEzg8PnSABBOdTiq/v/OTTuG94BALWMnscNm
9qmAq8xvnsbqp6hWStFiOnR6QsHXTODN0MG3MF1GL3BG9K/kJRk+QGmlpdD7hhJ5Sm7sIc2YCyzE
rlr5ynIbFfBkCdmUxixbb1aTjuLb+6dUxJ6gkA2CHTqPfbWBmQcJqS+7TopK5+ll24hx8cCUi3OU
rBUxt/lZXFGRQ9LTwesxhoyGSdwOQnCRQtmBZM2WGWcvZPiKnH05vccRpCxjgAXbrwwyJcG3AOab
3B6FIf1mezCS6F3MUbNDD//pXsdsXbpyzBh4LlwUhMIoXthBVM6Cx1akVI7Bl5pzPdvCCIUsGTpb
lhqvo9bjsZuLsEbHOEQtdV5eC6jzhm0fhmplJU9MQ29cBJxkL8Jyp5A0pqj6JW0ko2DomDrpevcO
G84cl5m0e3pbmxZ0bMl6ht1o/KfXYV8bRo7gkzG5VPkHUqdELTgB1BlsWZc8l8pEWWv+V+wW7gi0
FVpWlAbwaxftobf8YRN0SoIDmmPFPqDlnnrDKQNsQfavVcSIqEQP6clUjndV9kYh4EKg0T2+WQ4Y
GrwWh2ym+gd4bsan4YP6YwHiIhcMcjvJRo8VLDCtOHNY82KNKkntgbDeuGEk9nZF3buzcvP9/T4n
4fW59ER2GZGuVInkhCwUPTbJmGm3CoEc2xfN71UwfKJetKKeb7QYR++TxxBpbSLMUH7pt90VB2+W
GbTKzBGSQPqwz2oSmSsHEx3iK73THiP9YbSDkuK2RgNb8kMWc697Es+46TgzGeH4eH4DBspjRp5c
umw1aOgBFfqV/DVlBSj7Dv6eUC7nx29FNdC0b9C3A+JEOiWD+6uyhKAQ0spwWeUZmdv1YNeQY+8E
MY57WOI7n6f+SpqpcywhUGMS2R3BO4t4M1U1rE/jjAs4Cpn3GqMA4q47OAhBEW+J8t6x6wW1lSbZ
xUy1zUFx9i8PaaCkWa7A+KoLIg8q4MgOvPe/qUddKkzgVAChVkx/XI9BCnQodcjsjPohgigDAoBO
BDdOf/SeZWz89eZXv+jdAPNvi8Nhc6FGhvR76LCmoN7earQoY1THqvOzYIrWeCaKEsmw6qqhVTnF
nLU/Wo9sNxaDrLubae6JZHzUFzYoYaR8NKYrvnR5st3rVCfa/sPRPJ9ybYGrxMs6STJV+PtzienY
siuMEv02pMsreSXL/l+TbvwaEmx7RxdjiLXJwb+8bGK4MwdnQCbUKTr+MmJSfCvDhxjaEEPQGmMM
w8n6evNoX92w8D7ihjC0Y7zo8qi5MBPMny3YxTQ+4vWqdmk6HSjG9wnhexbFzqL34b82iR6jvYg1
VnkwcJq1Q1IdvNlHBN5EjNcZnYF+BaIFpn2K0CVvhpIn7oEWVtn3EBO8KJzNlwk7MTxj0so8ZfFt
VqNkRRtiPI3jeguGWIiGnm8OQKrqfrvoKij8hNW4qjaSLegx5UJO6meycszpfcUf5W5mTVl7piFg
Bqi/OGDTwftzydsCTlcNbvFOMrzZObVjQmxlmFJVD1ZUU1E+yXSIo3Hgg85XGT29nk+USH0xtwIn
uf/twHs5S/Q+JoQbi3nRB+IDIsCapweWmvrpFpPjRc/yp6RTPq0gf381f2bmab5wRqkYmBDoEV7D
0ZA1aQx35v54pmqlnvsRByNhyO458zN2eb66pm4lf0wCpPGxP4Atfx4/yJuLRhUBpJvvldZYAry0
Lqu4C4Woz7UTeHW4p7WO+quevs2Zl+zmzLROqMRdJ2E2G31DbT+TsTk/59948HJD2IYUZoa70MBj
S+KVC32UlW9PtBoWW8lA12BxoZpLfAnFNJuDiGLdeOnAQcPnNF0uP3x1Y9gMR4T2GFHUSq/eeIox
896akC/XaOEQ2F6RdCSus0VSB88oeP3FUrSn5hVqUPY62pmEZ30ml9E47ytk7qUjJepgCKW/vY3m
Nqs6uqx5jvapk+jptLvtYY6anIPX/0RAbTWebgt0cWHYLNIRICD7b5MDQ2jXGppupRrKNvuQhuMH
vefgDVp6Em9FlhX5Vm20Lqp/Fspf2ufX2839eW1/GnRg3wQQ9PWwhF43zley1frxxNCRWPT8DhEQ
WRqB7YuiJ/eA96LxhAIV0aZO2+do8CVSJcENfniJPy5/sDHq1MLB8bgFn2zBynmafv16E0IGPUr0
WBCgjPtN4PdGw65FeJUI+fsoSyoIAwJqzvqwQpO6Lob2BSdHCQQjarcr2MwJbTBAPZ36DFGdaHFh
CtnlMAr64cZ+URlU79+DtySj9zjSTX7rXAKFRlmJA1G8QcgUoupNbXIQ5fucw3vsTZK0kPkCiAV8
V96aQoXTC46C0Ie/G1YmczzK5ho4M9w9/f6aIwrW4sb7ghsx0WKlnI8NcwLbEjOW/CFRRUO9nFUA
qlD9geaOZ9KyJmrx8QRR0SiC51xqSbs0C2q5Vp+uNGqlwGiXICvQ1FmIsx71Ng0YeiENuMY/lXW4
4jlf9DUSIVal+UOMe6YOtbMEmZIbiu2ZXeBv9U/RBuvBLUGwrXgZ85hpvTY44sj4dxuJJqqc6yuv
ZtG4vhnzekgqWwy0zPIWKi445gLPMlPPJpCB7zxXCw1KHJamwrL5NszwrfoATzQNjWskAqJjqivv
kr9Pqqp4W77R8M3HUj3J1SY6uTaotRcW6rPGCpMXJyfzqorA/f0hSXkC06Anc3yPhPJkmHthN5Nw
4XOPThEmYNtyRPay/2Vfa6mw/neNXRJ6nJf34RXbpD+C1Ym2XG3ozYYaUS3gYYrP7girhlUoAOQ2
LPqpRIBkia9wB7H4nkFvMYwt+HbQQxgolO9eQgMK5ZGdDvG4bz2hmilH6ggz2jAyQ5i+Yf4hHZuJ
ENL+9ubO7an2dWIzfFY4rscvYCH63wkvfVGXz7Vkbg4WbEipC9GCVnARJTliunfd7UM1kAZoKc+G
tbAo+Bs3yPXyPlQdtIXHtue1NCDMmgKcTH7FTN+FE4tgl6diCT6cItyL91epGBAUc5f0LNxlQ1WF
Ou3ZsrUNcl51V+Yu77mhLVu4TxlKFG7SeBkX6Bf2rl0GE9tki9nP9xjPypV/5S73JIScEjmgXmw4
a+NkhgBiQajzKLmPCFW2pNF/Sb0xV4YUjemRXP1qwHKwf6xIVcBFKEewuzpv35qZS7h6m0IJ4h7G
04L6OahhHVI7aN7rYOsGeVN/+bBi13Ak2pF81L1XR8EYxotV9guro3bzpSP4rz4faNe6WIGwIcl6
UrdxpfzyISBnWlJgYDkYTYH1ViCtj++3CyfN0e+Q8ZVo+Y5cBDROv4HntcdeCZ0F1pB48x6E/R82
qhZwVb0Jqae1lXRvcDpcdFZmktSD9BB1QXwirebFYERC8W6Sp5x5sqS5ZQpE5mkdB8V1z8BsM5Rr
xuwtvv7nDK34bebcFiVZeM+BCE4DZQX4zqLw6g8eSCpPe6fl4DgFK29KVwg6SGirfsS4cXewuFZ1
syozNKOL2kl/E+OZ0i7NchqWSUyzcJhRaqUoYsdzMSHDGA9G2eTvJQrxfGdktZ3boK20MtIA66WE
Zgi7ixGiX1u3dBZSQhpgAi6OGsPOVfa2D+o8WvwFZqsy0Ph2A7yX6QRK0wQFVqThQRamq72yMBBA
ONE3f6R5/YfSmrawcJC9u+KkCayLx8kJ9gcAp+eGTEDavJXGKIjmWYtjSenATotcGSUS4ufQudT8
gwWKyJtrp2zHMgQgSMOXFzhPOOzFpJ5Xh6CTaO0fxLVZ0cN140g3PeRHU1ngiGWueja17R4Unil1
05QbpDSicwvTzOZyHQBsJmgDN5U03N86NG1YqFgLIOYxPOtpMfzYkaa0Vpdb1usULRCAQvE8yXjP
F/S0vXz8eEsniXrzPfdkIXpsoGQsFxUMCKNkRtbI4GOGeUQmjm1/OkKM1v0jy5Nfv23s/vWmKKYi
ndKhFwZ5WgSl2ZIl5JrWzYC1SZj5do66FzzMGRRrkQQ1P8H+r2ygsBr5Ai61BfwOvQK21Xw5+ox+
tvtX18qBL6qbPwzVSp9kkPHp+IIMMQe9U3YDZ/UpnXaLITz8Li4n/d00o6nzM22QndtYygGHhcBp
cU4Dxzzw+2R7OQM21wNO7IPSUZQfmmArUqFr5Q+KTujmHN3aIYyycazsxXuLluq/5QdcQSNpHUEV
I1Ayf8Kj7kZuwWI1HlauIf8t7wMI8Zrm2WlzeOQnadja17VC8YOClFvCoTKsPLXXg7mSvcVv7KOz
XmDD4lzJtKpwkDoyfWPE07EGrBT4tSZ3FCdrKDYCvO8f42mWOOE0kGAkXzzOydsPQQXe69VyDjDy
lGO9EFu8uflDCYO/DilF6crbuPIyG1q1WTcuSj+y3hFXmyWfZmSfKVxNHppLoxlnuLKiH8f0Ds2g
QA9mv0iCAfcNGC0GFudWW/K5siV4+ktrI39rznCATKiHRJ8t6yY660eJJ/Ukkobet0e30fIv6dh9
HiIiI3np4KOSTL3gwm39fZVwQyzrO5gHEsgjzzRvWP6ZkzyDlM2CJ7pjzJRGNadY2MuaZYev+PqF
r/Jso6Zv0JmqmtyqSWOjDoqgCuU75hBSjZXTCwInL6ee+Vo1a2NWXM1pCrY4+ZlLhjDz4iPnHQIS
3MK7aA7lMQF25bPT2zgCHnPo67Q8qZLMGaCetJuQLYcjPeli489HQBCFHwqyOmIrp4qrxcb6GTJv
AHL0r1MWsD8V+2AroshYscbxmoDbl1+Sbt+wj9oLOqoDR3NMqoos7L0jovBDo6Vv4pcSRYpHCQVw
Xnijwavvi9jjbnKjIAw4Fh+MtGBRYTZI2hHNtsY0vefGyygPJVNsHHyi9Y9fks6zD+J25fmmTQCK
Yy/1Tr4te8FVWZAgBJ0mG/+djpthr9ET+fKXxgenGjpvk1elBU9YmUembiDanzNzTVqh5k7lzjxh
KgPkC393wvQ/xHrSgkAwRC+Zi8ne+5qinCh+HXn2MTeoWvMEqJNUg/csxIudBpNj3OidYPkcMfOg
VO3qPreadAFVjvlOFbl13ywTAiC92WdTnge1G7Pa0b/fTAds01aTvUVzf4/mqYFeseZXmcrdPTDX
unJ/1FegTakKih05c5+oSe/+9ZCmYlctwO6Hgv2diEkcJt3TVXSS7ktFkg9rNbwv5+f3dpAtPyc2
pGrf9qtqUwPKSqWqPtp3rkJ4QWUVgQGmWLlS6EvDwij/e8Qza0hrfbprsHjT4qGlXlC242Olk2ZS
LHU0W1xUtvXO8zut1OVHors50dGWt6kUTIFPYC2AJLzYI94qPNXy+jfyvaVzbB2aZWYalBLrtnnx
yW7K+ravn/Sqz/lSadvRx96GYQZtVbRajh7pS4v0iF9glktSOg/40ZYKocec7hQoeTWnlDUlLLGb
CYBxIv9TBV5ae31t61/vAzh/c5RnZCV10dmAwc16kOAhOBI9zaGuJKOD3O7Cfta9pK/FulS5mTZh
l0uID/lo4GrrSvYET4bBXEYbzmgqI8OrmKabPhn2Y1rvIcSltZQckuK4dIYevDv8KGkfqgsuKURY
1l9/a+tA75aEe+M5cI/vspcM5wqfEUAUWiMCINNGyFD+hpxeVb/ieGOFd9OyNoRvOZ9IG8L4TxEw
mnELzkMHBcIn0Ob2rw2bELEkwoeEmV5uB1hbx6/NUp8d7af12hCepaz+MJaDC1UoqgSMJwN84hvz
1xLQACoBCKXZ4rpIk/vP59aZT+/H4EB0VWU3lvsmK+DxxidSvbtuEZG1XyBYBz/xY7oxaDPmrR31
wSmhf27geJh/puCGIt7JqGRsIpsC0WcDX4hNmLZwhpha2XCep57UHqoE22rK77m04/55k1DPS4rM
cBWVnfHbjz2GO1oNG83vB94t/nEs4t+bwfU8Z5q0osH6P/hZJ/HcQyWL+GjidJqCloVaJrFfjteV
JrBZH3OnF9bucigAId3YegMGGv8tKLhsA57jB4opnwz+o6HIO0btXZeLjAyJ6zbILHNP6Bhyzv4w
FjqPt9cao1C52o5arbIRBr+pUq02FEMHEqo/EB6K9gngGU8nZJFRY+m7cb2OJQPLn6KBMIh/FjS9
K8zdYdKe5J587BLMfhEHHg0hXYN/NcBHMcIKAiOBAd82FU33hY6Gx2GmyadDCOyI5mD8Kzi9h/cH
pZKk6S2/Q5pF//TXKzGNuGxFuoQo1Xz5fY+QRbprXDjhxwingvCbygBswR8LTwz524kqOpLOvGRY
CA+aKK+1EAwSAAfU/nCtcQ1tJtxIQ7X2IdnX1CMwdYB2WVFuiwyltB8kKULzJ1OXe+3EVMTapYRp
Hh2kXP8eUFb3D3ekWc5BTBsdR7XyCVFrVV4FbcgNqTYF9zQffAZ9sAwTcUhPAyh4aBGnzav65sRG
j1eVQQfn2wtqqGYFLogGTUrsrX8EzpU3V70zNm2TWLfJWf04sGMMsKzOaw5EIdQBzsJTpWiEL2hr
But4oFExTl/SEYjVSqpsGc3klJZsDu0+1CxLgzSLKehuLgxXsbcnamKSwW5dXT1Yjm8L5kOlxKrZ
d6oF0EhoQEUk4S8dWO8dtmCHF3v90WG7PCYB0wMsygDHnsfxBsjXwZ+zYxiFuT9kS7ikxfX3qw/o
TVLbQxTZoQP8uV7jq/9N0t/IOgVrZ+gFN4n2wsQ2cp4b1JsO95fwPTyEFCcgWjeiI6P1/j8tafYO
QZmIG9I0B42rlWBZh9t3Ipt7a9abS7R+ov9Qa3AoiRrqp5NqRICC3G4+MPS7S9FVcOJeh48Zb3SL
fRBAFPwePhqNMw5GEeZW5Q1udMo0mmp6VlNswVkEudzfP6ACXicL7+sRThcOvPIfu4LLdZw18KLW
ZD24hANX0W68w8XA7S+V+g4e/RgXqtOGjmufCuqjS5Jbz/xgazo6b9xZb7VIbj9NYmvPvswWJTz+
Gxwr03gSQdWE6C8hIKwo4kwu9Y6kj0Ar4o8mZUKqAxOY2UsfiAjAmKh+VBwz5AfBvRv0MGCnq/Lc
X1+8Wa2IdwEfdEVhxfW1wS82hsgwjB/cVwp4aRZiupjY7rfbTJA8GgCcxbRYb0IoDmdpWYPfSRGc
OiA2b42P3RqoIGXYS4Km39sj5nQrqYI5wH2e4alx9+6BevhA7Rn6w/pM+szlQh5S4KRGih+L9yUs
jqIWFt8eyxr9U44Mub6DUr9TE6RZOfzvjtJjfT7cJxBeMJFJoo4KO54AwK+B20j00BjS5HRibi+b
oHm1E0TXJOkbNHZ58JXcRqHZan5dqal+ilQAyZ2mMdMDBY9Df4Nk+kd9tL1RVUcF8PUBBOqqQvAa
R4LU+gATgenEjkek+fpjB0XsKnRAtFjaxInAl1V2/IQ/dg1rMBOtJPyo/zTCEC6KdxrmM7g+AAF9
iKMM1r47VNaUNYSiWtveQsX9SojxYSj8mbOGv2G65192+Q8D9BdzaaHlSPHnhWoz9tbFpLQ+/L8W
WAxFO5odNqlc/4SenhpY6+MP5alD1ilD+KpPe/95UTN+wX8cNoy9aVzZ0hW/XtBwoa6wa2NQlIkR
fTBHDuF51AckeNLeVLGRovJXqRDdk34LJMV9seRoiRWYWv3niNo5gCbcNMuGnN/FricAkOH0uFFO
zXW+EG6pQg1BiF/jj5uqUmHiieRJ6wlk0GYHIUgap+fq5tHo7AX4Sb8kHJc+03YDeVOE8TgXtejY
8dguqStj2Yvaj0TTTfyuk2YvHTvOzwbbfTjCtwgupsTYDa28BcxMBC+zDyXbUbyG4utA2suCV36Q
5d89uy7+PpSc1hIE5wFSvc0stu4FiGC5D440GiHWMGhQg2Ck2uxibiGeq/KPUvApbknTzPSJdzKF
6E9UWSYTAcjUPJODp+XIZUYjruBJ6jaGnmTILtf5oefHdo1fXUi0U7tuDdvqwCYrjpR/Kxqwrl4W
tAflP+pcoD28nhP2Ec8r6Rwynypjnswa7q3F+2xGLHaG0iuiiDEK9dcS3hf3IyOLEZK/Y5q8X+Pc
zN4UAmKV9rTQGa1RuFzq8dtLzaLyFYOVFAYrsz3gviyPYbLZJv3WAr/+RoeeZMq9U5sgknt3CECw
Zx8xhZZKXsOMAVfaUhQWfxmlMcBb+Gx3qx84vaIHDclJgWLL14R/m2pAwzmnyBc8GEYorJ2OiyuF
D/LxNz1u8UuQiLdZb5FAonxpiIJYT3Ly7NFIqdYS9lmBbz9fQ2VwZ/gBYbwRTAYZ74+ct66hkStA
yU101eKWW0Mi4a5geWrVOZYU7mxg44twkILjrnDzhjHstg2VqYmz7ffCaA8e8IwsgPekH7zmslan
zTcoS8Z7aLm7OLV5YCsAj5vGpaFdCQh/Y0EpOn6bNtPd4z3YfoChW4E+kkPgm2lolszv0++63Bye
z9GMQCJHTXTqxCJ86A273xBDZxQoKPtgfDk8560IxpsTi5+zdXTNLPZdwGVtg4fgGkddWjzK0U0X
LJVpXKlWMSx8pxfPywKUG8XFY5qfH8S1J8WpU4pQKNrKcA9AKKjPc3ubF/F/TbLJkH1vzJ6gx5BC
53kgcxKEK5jpRvhMuMdm4RKQbWphj/K0vDaOEIuCQcssD5gYYC/OFwI31igxXS12CUJD65gk9Zm5
n5YA/tGlu+zfoBNvzbPR06lhs6zmz50uP9t8ocn5wtrA/mL9j8fsYwBgl5NC2ERkWxEEAKJDfGzz
M0oCSYkqYR8i3/bKF1f9266GPh9TTxvHW4k4Djn/y0eOff2APTbed24Tb5juj5e+UbTNRkE+iFp7
yOEMaZxj1VvQzZwz5zjh8Czs+0wuvuD1r/twBA/vVlVUkN2AougK6c0NqfSfeCT+U3M1cP/Vh2vI
Yo4iuhrxyCrtuf85XWEUMvOm5EKzYCRga85HlSckpPm+Y6o1+PzzlVPotK7ztJ3ZeHEsz0H93jL4
u51L5ad6SkVg8+/X/NNMCVt3jpBAgPpFKOlgJHp2aUZIA99XAksQPOFV1HkiaA0+vesMpdt/WVn7
UO4yri0psudCmosYq8cT6n8cErY1QL3+XiSNp/+81e67cQbBCUoMylgEZky2/e9R4KeVh+LfLvn/
d4ULs85s09B0tS1cGDmFjsXE81o/yEtc9tKi/TLzKjehlLtLXgN7o90j6wHnOLFiEQc/4avKFgQW
S5GLj7rQYxTF9IlNcg2LYNm06EnxQWBCK2ZRAJ4SIvCFpFM46ifLhA8wewpXHlO8DrDAXpZ0S5Kd
p6dKWp3jfOWcS/12plkBZGK4G0Hb57oFj8RyEHUC01Pz2gLmU6h83CDOukYmMownzgofuX7H6q/t
WpDiiQFHKPEVDvwsJ/266y1wOVcH2BMO3amWjbQG9RKRwSqq8MrkQvk8ywkKn3ixZrHZRkKOPbFh
dKY/HuzdZ6IWFd5VEusfd+a6gnkxAD9Ve8a4ecfhX+P9kf6Oc6T4ObBGyO4uxeByd3FteEQh68DJ
1ehZQ9HeG/bhafyRY7y+++ZcuEsMa+/kzyPuBRPQiQN5YPlW984bOGgBnBgMbP7OqAjRSoJqDx6h
ySOmXGG1fNUndplqW/k57gIdhELjB00yiYetEc65zDG1Geco51Ex3epmk4qADxpitQqoeZppbLJC
hdOt+5pcvvdLNO+If/bte/lpBKKKFwXdTftGYwokDNDHtMe8LSkPVp31RnuaU7k3jRDK/Wc2s0TT
cejz9fQa3L5n4XlidAMbKjzZ0kZH12w1GPXhzvpoSROczYrqxAok/LpsvlNMIUfNM+7z6m1XEijI
xR/NX89nwzkecJQPpCRyXwkdI31uYnODEzeLFNoxPgH3jHvlQXau0nXlBjcLQtsN6Bm63lXKwv+N
/KVUfQTXoH/m+TSKugxWrtNHSCLgCXzXCbRFuyW+TwemX9ZrWB3rXnX36llzrgYxnRKS759l3SfQ
h6W3vnCyqgQ+3BU86ZSr507Evg8wtk4nvSVsh2yAjaKynSkEuTzqSyjeRhmxmUP0IcJ85f3Iqoxx
Ii7dEermjNdIT78vTLMnCNDhC0TbeX4GTxV1fgbvz96HOl+nDioP3XwaSh2d7lb34HuxbWI/tPG1
nTBhjJGbq7kl4VKCzTk0z2A+Eu8Gd0fuS7Nx005zulO5atqhVO8OKK1skHhw1TluSscyldhFQ8so
hXjAF7B+PZjWi1HQSAXPhlI5Uj0px+jMuKjnzcvH9X0HsQutLDW4wxJl4iS169dYQe+IvHqYC38n
drFzSqKS2fd3mlvX7M/1H2ncZCdaxiP3SdINsB6f62yJDR+tXQf+fEcq9oFD33vGdj+QcHZQdFq5
BhMMAZVrhjTM6SyICTfEkLf9r8Ai0IHHg11uZkIPcSl3Fc4rkse5OnJMjFQm7SNWGY/rfp9xGERG
BCAc0fZn5wwtxZTB6Fm/Jp908fe47+03UtpZ5yLkubb6zmliEDMYJZMyfwF7q1oebWH7Woh1QdL/
Xg5Pfeh78fNHx69fae9oH7x1cKLRNyQ1JX3jf25p+E3imnSs9JffHZFzeUxTO+cgVjWL6Np9fFb2
0ozWbT1MOhDN3bCocTYxaO4LGVSTodc92q8u63rk2yT1HHnC9v15/RwpLWJzQuRoNkMGvrBXedfM
des4KDsWqTHB7qcG1TOPzG1Szke+erja9DX0FRRvgxTERBY781839D/iMYwnfL6W9jL6DOQG8BL4
QwLNmtoWqca/Zez8txa7TT/+N5ed1uaX7FXQWOlrDOCVHn9QVEFNID9OYsVd336UBPvgv0e7gau1
1fctT4B1aqoNNZdbLxGafdoK2YQ0OYFUlu7VMfkjZ3nh7YwdzfqpKqJfKRPN6qmGBdTWQguBCrNy
PPGZq4RL++3zNgF0Nln4XnqNMddEUJ6JPf0zaq/GOWxIvHcCeV6KrdSNZcNKtTNc/RN3aFyXtCcA
EeNFSQm15RtVluNAqpmRe9s+edXcBtqWrB/v7KzCJePyp2WGKPqvWSaCmvS+D+1Q0YQjEoOs/DVt
WL/eGwz3gAVemyaJzT6ZqiPB/X/Y/TRqKzB8HLVWf3GoWSZjzXfBP0UX3zTYLIHkJ94DoS9f9PlM
ZlMEwPQ2A9TkHYqkrRBJeyCcot2Bt2wBnldJhBTQ+uqey7RsJU/ZTN1+YGXdIc+komZli95vCp8n
JlcIWtcxVI6Hj9Z0lNKgxaxgRszubSVedKee/FvMt8PF1QSxUvx3mhxCZ6PiuwrzVyyZZROgKz9a
Tmdw5M0D1a1Z9h9BNACLO+Ax0nNy4u1Wfn0Ph3z3R+H6H1eApg+YaYrpwcBnMDtzvg04cDMzOZ5p
kqh7oW7C4IdB0PrEcC7pm6R9Ak8z0245mC6d4hADgKaxUmcLWODP315ufm/3Nd3GMcXKkY3ys6T4
ZthyMz7VBEkXH+2tdKJfmKZWPTUxRCxmpq8bAV6SHM7Q9lNV7f17c/9NKJrV1iitG/9w4iffKCdu
mThJpmH7EKK4osW9XctJNL5omT5Ii6nD1Ze2KL3my2Ua/ffnwL5jbCYdyxJ0uusCzsE8t0weeeb9
f70fVYLveKDjODLXPq1OkFU4y7NrFgT4cFh/NydIyBjU4UKjNVdyNwlUK9ni/WlcWOem+oNzzVS9
5+ni0UH5Q+AwhOqJldQgiwldWoPEBBOXFGlmV2bkmI3UiVEQZ8WvOVZve69DoK2NP6lsCRcrMjVu
iJLtnk59DWFSbmD5OEhhYVVBNViE3oEBzvAMUx0wyjkasIDy7HTGiqio40UELk9PcBnxkDDCb7zG
jil4ddsU990G24iDUnHvPOIQfVF0+PF6Bt/syXibTxkE5z56UJgJ/j4ceFu0KcYk0YFhf8sGfmqn
Ajsg0a8RlSzhTPbkq7vBya70XNcEssHYJheMU0OyaBO3M9gCyzPpUNP0PH+4FjErVxKkuU4rOgte
oDCqEMFBwRm9JPt2HCNHfRQKYw4BtVDEEux13xa574SQh2RgrmjPemb/JTwQTytS+50zdemZRqCV
G8e4BK9FIT+XoYNu4cq2jOtCS1L6TfnxY4c82wzI+70oDV/Cp++Ktn+lIYg3DxZ/oiYB5JPQpRV2
32w7FcV7x6XWqviofwYbPEtW3PxA2e2ne4Y18CqMJ/DMERsMPg4B8S1plPKQm6rdJ47Km0cg5fkF
5GWV9C5Yo0fWm8BEc7kzxvW04PGeiTB32V26rI560zdvSKowVLYbsbk37v7iCyEWt57fjNDnMSlo
KHW2Myuyy77XPr+w9gxM4p3wT2ClaoekRCK1eBmn0ECVrAL3+aVcnvJsXo2sAl95bQiRnAGkoI8a
VMf9Z1G4OKVV3Wed+z5vGCoVVNbHi3Gx9eydljKJbxAvPocCSSPIJkG2khbHWyfkFPzZAwoeS+b4
aLmnEN4kEZS1Vv7vBHnRS4G4ED/prYNSZKpoKGwqgEI2lgrAdtdSI12urPKk6LfRVSuaTgMViBKK
ao/ziZhGUO2cjlJ2CiIgctk8xE8HU9hAVBARorL8SabJo4Hsz/nr/VPxpWAXLLelIQyZ21HVXRo2
6wO2MfAZvKRhwehHaeoQRCDXN7Ejj6zmU0EVAxVsFY1MtNbSflbPh6ax2HTSy5Ym8G3fd3t1PgiG
COmhlz6BkM3lO5TtFWfjqZkqklO412zGNEa5Sydp3A2H16HP/Ne97fbPHhpkfz1ySpY0+BOyAi3P
tNEKtnoCO2Tni7H1MtZYFDOppYlCVBqEcpGTBrmMkXN1Y7FPzh7sBMg7oO9HiP01imXuKYceJxSC
C9GaWqxqeyLjoRC65oes/zVt3FHeVWiHQDxXczl+I/WmGHeLipIbThYFwUQ19BftLQYeRk6wdfm7
uNJyKBCsphvpExQP784XcJAhda1xQgFj9wyWW+PY8B+yvXArSPtL1PnIi9r1QaNsqarEi0w4v5t/
6aubQyMRdwbRZIYikRi+OvjJek7A7xYDcFMPC/8Z34qLqSErywSgdBje9q20bqb7irf64UxbZYe2
0y1V682y2vhwIxDblH24WiX2AqhlGCv5zlmqS/fIqFE6EJ7ENs58D0kMBZAmYIJ6V4KPxw2Hs6ra
/vRoVwQGnBriOMf87pxfSZzk/lqHAI4hjlT7+bCe1XhhQqN4ghPuf70ri1+8wq3sLYjOaUP8KDGq
7JpsSF4+2+IpLQebcYMBG9UXipizqEoBpT/ftrcVBiZzhrwpUsoIOcyDsfaLZzyjL8ELSoqv5b1q
AAE577zTlnexA2ymwz4MkIgyHGcDfZ9mAh8PWuey9sd60TDYL53OaaU3TV2zE5qkgjg2lHSox6TC
2DiPwfWFBrPCrvIIk3fJ3pQkxv8iuEzErcQ/KQFeVehElIaEHPLKN0rjPEwA0qoYAFFa2sP1rAaO
oFRXDKpCdJjvD3YakIKJg8nrCgTuvg+Up67WJqM8pxeXRxvX+xhAgMadDh0FZv2kHOj/05Gk1OZW
lKBRKokA6UKv+mxBQXIazi1vYPhMjJUI/6r1mB5B61MZftm4X0M0OJDi9MRYvYTWQ7+CQN/4Zljm
Zphn+N1scJaltUYvyoImNz47luIsAyp6LwluTRS7SxB9aZ/h6a+NvOpMfjpyIuHgOKZV6qPMRT8t
D37Pim2PH/nYHGAzH0nZPF8ZOFlNadds64XSnr80ClIYp9vouHdIWOokIOnK8HAmJNDMsOzd7K53
HB2tlJWY5g/Mnq3q4p5JmSk40CU+dm4kWe2lgOw4MnR1Xmi+6VXwuQYB28psZVHPXLMIKc0kkgCq
8Klp43Sjsp2vbSgF/wuu4MmK/UvybRaMZc7OsrCwhlxq8JwoyHZRSAJpGupVqL9JpD69DpaIpdAA
/gWt4VxgkNJA3JrDj0DBzhbFUxSc27Qz3YXJRL249EibFJIXC7I6OA/uFD6qXau7pqnS4Eil9ex8
RJaBW1ME2pNZeSd3hFOUlozKhsO/AzgLCUzSrZnOo1zX9uLWbmEBCvfIQC4svlfAQMTUwQmAAmiz
S9nJdg/SzMeetThZ8So8T6ARP0xUTAy+nl/nbbwIHMh91Rom4UMaQ82zSAPm1l/91HL5GhRfZTzj
+zh36iSoExLX3oReNZ/wGHa6k1q5duDnnAb4K+53SSmE+p5RQNBg9uDFov1xvMQ0vxAit3y+pe2n
hMRpL2kCw9HdLlyRGoNXVDLMxWjCTfRqTsc5TZfEhg99iYh3aN4sX0INT2xRP5EvUYgAYir3kRh6
PiEHNrP9M9E7rfD9XB0I2gN4jgKrdi6GSUSnUluSQb/BOB9OmUxowobQpd9Zb9tjn/QbgStslTCX
1caoHZqC/Zo7ct6OC1hux/Mrd2IooLedJx44BJjSbJcgG2/+Vd98NNoR9UwPTEYSi+OzXAQa+OsI
AwGcHPUQ7CC2+IX78nL8I9LpUBsuhFkMxXrfDn+A5fgnMdBbbomyxGJgaczNiV6m91fb6gmZPoPc
uAolPAc/nejmzaPeXwclOsXRBmgl/AYRjITxRRkKhGwPi6YbhIBLO2lg1RRRLxQ8MFOR22RQhZl6
imGe+SgpJwsUsc30J/BM2bGNSFs5QObyW3IZn5o6DSgPanbeZu+s40QnyhQYUmXV01eaOU0m8hP2
44bxiE2oMzWfvvTjx010JVbC7xyVhp0Ged7I4qLFu3PywJmeWcX5RwW279o54EUj39eWaC/e8xBe
sziYvRjf4JHfz5pjd/av9n6w6K1tDRfMdnMJALLRfg0WAiF1Ke5/fgFWVJhIsEyuJwJm10ISCAh7
TiUHD8tg/u9p1SyCGYMTedcsMPpKFFh7XsH7K9WM8eUD1cI7T3F+aEuBAzYauYLcXv4PhtfT/uHl
YkAjzFriA4micXTgacx6B1Yc6FCK0YmsnSzKf8Rfpt7hGufd1CFR6e5T2lNtP3htFkcqLH6rGu52
9D+VzKi8O2PuHVU0BQwMax1B1u7cz8y2yA8x+UVHBIaDjhptvKtpTKG/6z3kIp18mnwNt0zXEe/u
nmicqUw9LWmyEzYn+t0aFq1EOM756iI/nQiPZ8+J2PKXzvn6ZT4mR16K2U5Xi1+0fKIG8nV3heoh
zcen2Uc5LHy0ODciaWj2m9/AsfLxkiE6woBLEpnr5sEh4kSa7gQZpgGwWDr7gnrEpFWhj77wG9fH
sgkTHnuKHlTHuDBr9sc3RAuPeWbD4kC0OPpg6QVexn1JdBOD1TivpwstUnDCXt+ln06lttgZoftu
qikPg6rUO2i4ki2ADA7znTsYkvfe+HCJVqdtyzmADEaQ1t/bD+qsj1F0TErYq5xefi3Uh2C+M8PH
D5qH0cWY/XIBLHG12RHtYCmK7644PBoXTRfixLVTlds5IkeqUk8muZX/kJWgIpkFjsBU7/mXIKzw
ziWO0d1CvtasWcITjcDSnjbQpUQPIEa9nWHMWg5wUlajvtST70PaOBLjOaEfL1T/pnPRWC0/38K5
we0w5hiFdRMVoki9+3KnI9BftwesLUoA/gbw5VD08ws/VplGmPBW+7EW6/Lbf8+AhwfJYQ0m/47T
eKxogNJtjl+mU9K7+CZoNdfLI9P4G5DaBQjPLY+tlxrZLRbQVkEowALObqAqgjf/ISy92gHxKtVa
RM19ci3nLWkSq0CJ6bVqu9SKuszfdzL7MAC05ROHZD4YLRBO8yRbeeEMjlTLGweeQjbdm21Ct4tn
SmjjWoaLzFt3GB5QcjNGjJZu56n+3edwyltcUltm2PTCV1+9fPAtgZnIWRoSRuS1nrhLiBY3loOz
/1UldUoQcyDMUDdDI5FAiMkppfST6etE154hpKllkKvIamppAArHrGCU7cUjLBCUguwdw2+qWJct
n/FSkAQ34nYPRdzkTx1sDHcVn7qCORgISffewgrvro5Q6Gn40CkbjxygujRYN4C0OgOt6m/Og3xD
SYMFlrr30OQmsOMexXyk8XsSEo4nDd3lH+ykW/MDuAnQJzkln5ViWuwXEidYiZc3F7QDd3pfazXB
BLHZdbLXWUr1GyJ/9cWQSzV2gZFCHJftHf3GHHK2PtveFzHZdZmGLi0BhnuGGtyWOnc7y55oMJsq
I0fA2pK+H71N2TLUatPaVH1+isLOC8dN6dHL1r4w2mhkskt1MzYxQftPG3Sh8+wx2MRkeYW5DYB8
km/RnYtkyxsZdb7hmXXhgnZedKI2HSok0SmJaersdVpAXvm/bz4H8kfZJWkfDFG/OsltJhqkmffj
1Brem/SRF301ahPoaYjpBjHefWIKQcDL45tXsh8SYMXgp+wfO77cEU/+OH7gZzTcSoHPJG70XMRi
jUNAlpxfFppV7At7v3ejMFdnx/Cypw+NkZvFlcXerqkuUiz5i4YjI/RfwBmINCuVBLRgyCG5IpuK
JEpzg8BaCx83rxl/C35iCsTNtdvXoRWhhHuAikPbr+R1izqMt0d+tL0xruaon/62GqXM3r/rFpB3
hnRVSm0l3F5cs09ElLgMap77gWuIiyoyQoTKbiyCD1+aTk9OB6Z2hu5caLJHPn2iRllC9VdI6JdE
i/ebHdvlorFwlTclBWFtNOOPQNIJFAdj5IWGg/N2OIaZx6NHFQBOGyy4kkU+kSy6slFRXVSAhQEs
WtT73bXL7ZKvZ/vKE+vC8mf/8OwDv8qc4yfP/AncvGwkvgerOMxx7Nb+L85YB2PbfTOLt7KvZWju
sU+49zhth2pYn8sJHwopJOCH6OWxBTpJ5rFVZsA/MAW72GKrqGVTgjF1ibz6Q/6NsjKhS2i66lPI
PaNSewcUpxDtkJTedgSl+d4O4Vw4QZHhuTvtTv4pzg3lxWB76jShLnFMck7iWprS0qCbSx2ED0+y
QRLW0ctvrXPlENlnrbwhliw2fPJOPsPi0EJznu8IQIZSNXgMHypquWdGk7XSqa2aaxWLt2/ZfU1J
DNaZ55iQZ9DjrRCgSxbIab8hpBJS8LMN9tHEsYihuM0HFHVgGDOXpFz9oQOXRtzT/EjD0UKZF9/C
F/bjK98oz6TgnBEwx6TBLc7aqtbTbsX9RNGi+oHpjMyRCIiAMa4+u71NezJiUtc6k87RAui0xie2
E1d/njz19+h/MIs+s2FZYVyalLMcbv7NFhY2hmegRriFtKPp1EclIbI/c5Tsuq9nUYcdusl5ZGY0
/FRYTOPyMjMr/Oge0OTyIZi2N5WOBQn7Aqz2i7MFWE3i3enYWs/SAYmi7a4uLWtv5Pk66fWbvdA9
ChVUqZ73om7nWyMnv1L8kzGlrOb9lHR189B3bqBdj6q5JpBIywpUMK+vexpza2g/KOmZY6ZhhCO/
6WeqcOJOUKYwDd8C8NCT2sFTg4hY9kohXqwLRZToolHyrQkvV8a/cVybrrvL9Bu8hMwl36bVgw/c
UlvjzN2upB/l+M8XIMA1Xig569tuO26lc7YWU0Y1qh9Efy/69CZJi8iwJihVlGFnGvIjOeSyctdI
ty6iPOn/Td4Nv7oQkO0qRAQehyMdv5tpU0zdobR0TioSxyPNmzTqbvEE1ev1PTbhW0AGSkCFwp+j
oALMOtg3MM2cfWnTuvvE2KYOnmxCB1HYj8hr33SFlNox4jPhGhIxurepCtyNys8RfJz4n3gZ/536
0MHoSxZdRdxIxi0g/XQ+eppdlt2SPH07RuLgZDPjxWm7s48DmO4PgwEVEoDfJccBgjKZop43U9OL
1RlhCUsnI5Qs9/Su5O1q7LfVD0L3KGK+uJMsISoMO8f0sxYTqPfm6qnVTLlqYBQq9KseFwUcOEMc
pOX3uYhPUm1POISjm5IKKLbVEgi4Mw7fyr+1DYr+aXN29P5wK8biXoLeyFqTL/RxzaaNx5k8OhDg
5yDVPq+Q1tw4FlDvzzhkV1uOg/1iowtIeaBthM8laa/fefXfJs4AKbDGBwSE8JS/3bY46Tyt7GfB
0I75ey4I3KXJB2Xutm/rzgT3xEMIpcUujnk4i/dWoS6QSzdvz2lY/YgGc82MqYBSw9g7ie+rvgof
8EmLq/3yBHt+MbU5sMP0s81WNLAGqQEQ5SIx6KG/uDtOwophpHzmUZMWT8lBMtfnZVnhzJogfH05
Kj5Pp8h8He+GSI/SXNTDeAXfBBGK+zZwnocc69KmSAfVMH0BrXs1T1btCbcyD1VIqTJNxoL1/Z9+
Xe7bnaxvgtqQyu0QAmKM1jk+YJujJgakC+Xtz4JHdOOPCyWE81fA8Gmf5RIT5DyoZ6HWvwlWeTgx
RmKGYL5F5dGhbG8Y2MsoM1chJFsvceVXqYJnkI1rkgA78tihqojqvJNnJTkHqFfvb91OzDLScQwx
ljcq0MYsHY8GaA0Nl06wxWq78vglLBtZ1+Mld80jZSKZ8UsVjPc8ehTza65QYHYTMtzWSuR09BEe
uLLS92LQOYcHUQB0slyFJIBaAFiIipV3zMV42KdmHqXH/zW0KcObZKJ01FU/1g9K4AC1yM1dMtbL
tHwvyQ5/Dni/N37QkJV0uw2z87WE5nj5l0+j/+GtJWUPOATE9bfTDxCVgrS4Ya37uvMDpPb7UMpD
/XUzUJyHNYergBVaIhHqAyT/DV0VGPAAPccrDARiaqCU65Lb7IpjG9QcZBkyXTWOdsh67CSDA4rR
EL16wV7/7dtj+B48gm04fVl7Blof2IRCmmqIMAFQHaD7HocDad2fooAHmgn2gT//d9MmPSEnQp7s
iFN+asRTHuSon5Xh7TDMaVio2R/rEZSPutxZUAwVVmj9mPl2WcKlI/N9nhK44t5kJMyt4qUrUobA
pzlmeDNRswkzNMG8z3HTbKAugIoMQkXLg9dQxnciLABt3984Q/fIGrugH+u226UFUfGcNextdnZi
3AQzuv7cBxRmMFKzbPl32Lhv2FeAszf4Lw435DevIy0+iOuyfnEUqaLbID2tSFrvHz0JjKbH7h4O
r1pmcoW0k/vlhiqobJJrWLz15E/V620b7c9NimYDvK+SXYWnPeiqsUs7ZSkTqDeqGSUsFDcONYeO
vk4O4aLZ0zoNxREituFdq3nNbgvS6DbyRbOR3VOukFRingK2IajeGuFbMYZ36QO7jUphG59ZkY+T
UZ8xMnRnfLuR7XSHy5HtVzco8b7NItG+IRz8n1hV7CEYljZ+HaejC+gkWBV3u1RYcRofMlyu9Lr/
tUZ62jPdUhIp2WGQLX0uckvxPWNrQUrJfqmrwjGGTeh926t7YMOgfYPDAW5CxQ0XfGF4pFS1dhbJ
wOILsbPZpkFN3OQrf8HR7jNjsnM4nf2AOYUgjGtVMm1xBe52cCCDDm3Ja8u2i0Wf64yvfP9UV/dJ
/lnOy4tGO64AoXv2vvF9XOC9MZpY7Y++loFO0noTAaiQnOBsyULd+ebWwXsUChad1AdPCxbrm0ZO
4LeglF7PP895FwNw8u7SrVmSHh39GnmhVdnHG0rxO5qPbgI6HuOMa2GfXSz4xkVH/HhA1R5xSySk
gMHpzm4D0/0mzb4wdQY0nWN6X/45RJhHnDb+eQhpVmkZnn81CZI0sQmDqZ2cwLUN+N+LpiTXVJqv
B4qvYpwZTKrOKWFuvTRmLwBeSOqeAbOk4ZZo8JwuH/4NBs0Wv+XUo9kFHRIHskc03GePbL2UDmKK
uTniw1wLA1CxknASSEopARZWD0BEuZiPE2ReZjY64EvSSRCC4ICkQZWzfZXFbebe0jzEkTREuR+u
LkF7MSB8cr0S60x2aMa7B955wIM8Kcb38D0fdxgTWiLhzcf21srHfifmfZwcDtCItNpIx7ptA3ti
sa3Rgj3+RsdnKdvUPHB8hklSsNuondvKsf/As7f29x/vJoGKBQ13N8RKJqZOD03Kwr0SV8VteX9+
MrrzaWu64Kf990KONGENO2UX1ILh5QO7wA2XgcES0IM8SUSZDIE+hQRtQ87eWavm01ZRUdB6Xj+n
u/meFMS3NtJve7VfzmAN3lCHOtpPHJ+YLyO+ZsghP+dz6FPiULjnEoLQ1liIHfuB7kCFICaxZBk0
Ktwhdx9Db8azZ+tH78PBiZxWQvWDojPdpozpXup6Bwx4bn8+iCJV8vF4GVKuE8ALkBhWgL0ZMiP8
O9AVwIVT0cnPc1ZZscSmvy9j/o15xV7fpXbh86nXVLbph8WuruNQyqKgf4nFX9fQQCqEpm+eMugv
UNVOGT83CXR6NvflBXMGDVsUnfCGgkHTZT30Bh01B7pN9iadKhapLxbpZdfQdxeNi+St/wwfCjhM
0OGbkE53C6F5glDDbB/QpWcWBGuq8GEbBqseTeiSjgr+QQV4xkpanERucYPuD6T+RvKtDB49bVIE
WQ/YSfoz9j7ys3jYsmTlGOE8wsceBHssPcQcbDjvCKUnOdmXiWVqb+/u/ElKB/kMBzJwYh9JzxNl
9eMdXmAd/0ImQ0sfeiSgry1XfIavz9f0K76wQWWD4NC9DOgGxyTVBRnmWLomDQBEDuFHlKGmFvGw
rhhXLYR4Li50v32Z+1xznr5wXa3ZISWpEX8nmZAFOrG+rIPxoSqCh6K1YCsVW9UN2DZNeqIQ4qBP
7sEZA+lDAOTWU+j7CQf3r0DH3jMED435owBYPYZhDdT+aLbkuQuF3o69HuXzUgsmboj/Bs3X8gVF
ZgvHV0B3rXUIBHh+MB91sjQwLDl2t3m24d4sBZPjTafTh9tFChf2Wk8f/XIgY6v8rRYtxZWCtSuE
JUonPVlCn99/4h7q+6ppqRxCKmPV4fHXZ2ykxzaoLRcWoCWIsuY2Z793WfibztAwakmhqOQM+qI/
eGIohkCkLZmygMUr2IGEr8j/vekIHHeKwSTySgOkEXBYZhqhbDjfajJyItqqsla1bamxcH/vXphL
vwQRvyIL/XgeWoG+A8S4XgP/HfhdqtyfpY1N0DcYIObfVg3e0jPxgLYCNifO9IAtHm4cjSEpgOY2
baODa9Lk5yXlL8xR45wXwyeL1NhWJHslZ/U87cAms+cPVaHRndyRsQBXciVnJxA/pGBk0z5E5+cC
ScQqrfQ/Wt2u3F3Pmf2wFHldWLF3BGSNBfjnYTvYgjn7ZoasnGJOYjgeyvTDdX2CmQ/Yy+BZQhWo
Q78CuiNA2h91udpFdE5TAxSw5kgzmplaMae4Qg/hgwJsDBs2/F61cclkS5BUmyNNzj+Z3MN/+/oH
HgCL3H9ZKWa+ho6FPNEBtAPyG5zX76wVfAPoEwoYQTQn9X1p5Rx+Mcd0aAOFh4l5QOe85kQr+wO9
u0+VKZU1bIPT044ITujZ2kgMFrGzZaH1GDFyTtcvV2medB/s9DB+YtOJG8bT8sPcPfjHrbe5j0eD
r/5PFZhDyyZ9aEH5vm50HYhoqcX6x2dwytz8rjIAvXZyZD0mu2gCjvYgs3ZL4LnW31I9SXoUjnsM
l/piQMfXKM3LatY48lRVtlvUZHibYqip5sas2W5jddgSd5dfjjOwV3t+Mym96iB7GhGha6ulppTC
aABm2+wPBXtisotBSlBaW37gLS+aJ5VGczCsJjZqDVl679AeF5MVeUGUCnCyhBGtzfjOPCMci1+c
9rguCbZruJPRKvRmKKOTPtWqEyhH2scJfu8q51MEK5TMMS70AC5MwnFLpsVjLeFvxuriwLs52lsd
kbKH/+5rqMD+QMPDDX6J+Fx0Ws6H13cOSqExIGxyV24iehO3SschrjVL8Ctt6uKZwP9Tnxqg7UGi
uoSQl0hnIckpKkuG2GImXvSV97Y9hMvfcnxhBhoFmkQGYCRniQDPMJFaY0TMEymnGRh5gZFh7SLy
xUHzmkB1Ld+Zdj2DvgiGKNzRD/SK2M3yQWFspiBUQ+pvwj7NpsI8ACdzGfdQQ8APijSZByrZ6dee
TqL1RB2/bKGa2IHSlot35wilj0FS2hfd4uwF6f9Lqix+axEV7KLTi1+f8rzbjzQltzHyzlPebTo1
lATkPfuSVWmOoqX9zc73X7qJr2Ey7mE718u5XZrUavzFT0jreOeQx/pImwljO/jdtr59kiDD0beU
9ljMAsKkcgeVFefJYe4mEXT9Uq89rAvQRXvW5RTyPDrjZdIa5BFMBWZHiu5pn62gtvFdXsf6HfX3
G7RZnIfigXr12BaAOgdI7tK+9tMdbM44aihS4+g6xUHlBIzNARGLe0ZNFUGfajOiuTcnlgu/Y2SJ
aNtialYUB6U4nYXHNfyGOANgCUxZodNPjXQVdvMiO/MtGKlE8JjoE8+jpqfoFdSXjSeTZaO63rjF
1XcJjWMQ/hfIdGQ7R9LWbOKlty54b3Mhf3qpXJT+5hvd/bBtf9DsJ95fwXlgJ122y66XnxbgP0J3
qYfa1m09+nRW8CmJ03uU4pFm4Z/GCv0Xg2GcIdbhCmXhwwWJDWMxgpIZhI61EOFYnS1gTNSvQy/S
pHLD1JzNxRf5zBOKoEuA7p++TvQX7rMALNy4V9NaHqPWwPxLS99iX/CjMZzKo7ck9Z0x7JecPmBN
MYl/NAF7puFiiInWsqcVvMydkItKiC0gulE4i7Pau2fGwSlrNiD+Kuo5OykSNxkUeav6JwvFv0QN
jCJO8JjRoZ7AtIA2h5f5e5qjd9FCSH+iEe6U9o8n4e77nSnTJFGO36AoQ+Pkc2drxrqnJG8Uqt0q
wMV+1KdX7sRO2njdZ36MkERkXIfXUtF885/J2CFbxvLnrW74KdsnaQ/26NCX5+Vcva0njjjQ1QDS
WGxN3cEHMYE4Gs7HII+3HBvNv9W/kOU3aBHiPelHR2CmKIX8rK2RmVERJTgTn01BIhgyvOen1Vbx
bZdbITif5ujPG6VJu88JchUZteQ1Zu9oHzcLfsi65WnfBlRWYVz5cRhNYV1o5E4bdBoAgGfI3Naf
a/p747gUxJ8hflKESpbgOqSqNePpam4nxB5z4sLH+13wM2P4kmjT32VR78+u3+Q4gcyBcay4OhSi
RTJhWkXzjF5fRoBQBOkXQ0PrCg3IbbOkycEKKtS+tAwfQnmf3RDlOIkxX1C2shXxQ/4a/WIRBns8
tilkmF5wqgcGDm8Q4J9lIivh5mL99/jmyKyZvUatftVd4K3HWRF41lByW2qs5EFWoa+s9xSZI6nx
eovwVZz9HwVk6qFWv0TJxcdiBOZSX9rOe9E+eYZGDcHsRdRJXuQxe85XAh/oVQE82bqQhwfvw9c+
xaXGA1qQJItIRdC9TtX3cVT3e3uO1Y2ontGga2pEV0OCR5wk/ImpBIgHrVWXHSGSl8gla8Sw4I2M
F3u9J9IYcpVQKTYoxl1RZpLUXx2PSZ5pZ0DCGbcF1w0PZpIo/gCE9V/0acJ5NbfPLYN+mAI6Fxwe
l0dpSv3TR7fS+sLSRmvVcApdqCRufIY2IL13uE/ZvgU7GIPk9O4fp8P/QpF1g99MnvMwtCWm9QPq
M+HgBo3CUe7cpzNYjqYPizXm9K3nbApo3wi5kToKFMdjPi047t6A5nf8u28NgE7YCUSBexE+DzWO
ayxAb04GheN2WQs1k2myVOAafCQwC6ogcXcqyeclvi9MAoR2DCQDczIMMDZHAHd47N4UCfis5jgv
1ZnmEw2hfd+eYZyvTCai3JWz56XXmROVZuxbW0BZ4h51SkYVznPKmfc7ffsVUL0XGNte13tU26DW
t+k0XARw1Bo7Nmmf/HEUhb3I3y+2RKDfamy8JuLMDjB+OdXJtzfG9fcB+LrnfnpMhNIniTUtgibM
L7Vq0ojoSaLLDcTU1rzlI7wZEjZB+rDcMS6FYukW5t8hi7k3ZwPk+anEZMmza6JBKHf3qsvePrDZ
gG02LZtnLNXx8t86dSBhgnRsDudx/B5sv5g/JVCX6L+GlXk/F2b1rhsXUFjattaXKkDxBG1WmAV1
XurEsyyZuBdrETEGr54yH7TAXMJ4ZebQWf4ENzoLcODaR0vd+JDJ0ouLtX4d/XE1UvQnmbT8/yJu
Lw8UlZVhkoV+6U5RS4wjT9aMo8ZGxienz1rLJOVrtdFJMCYHxXi1u/B4JSw0hV3IgRumCwGKkddO
TNZW5DOt8aRbtQp6driSk99Mb6bqzCYJS85C/TaqXR3Ons3lfjtnij7AScuF+XkwsRKVsr+fWtat
TMi5BsuDFQ6vE9jovzO74tp596/7657tYuUN7xJRfrmj75hxPpumtIZukEyWrvnJICxEQPosDByi
7YjRUkwAIEY40t2Mw0M7TrRyKGvGQVKKgH8yz6KEPy8/KplHj4DAcZ2RE8q1MFk6xrcBENX7NT4Y
Y4+zxvHP9imaetVWXR+XedYuJqcOkNxxT5JB5wHts/H5bgRvJeP64MxVhE7Q5S+OE4WVev21psXX
xHzxPuI+BLzj5aJji42RsK8bJKnkllI5EdlK6wXKiH3YDAUH+N1n73mXReuH6kAxjQISd5WWuHH0
4R88UuPxdYJBIHjjf32Bm8Hyseebj9Finkjpa2HEsTbl42zUI4NiJNNmjPLE53AJJeNMkwyeR7bd
33lM393h/+Ddyq1N9kiWKIz9YOnFdMDmSLXQmeKEwLL8g9rjuBaYsEQIbUUQrPynCy/cjrbSzwjz
mHOxBsT5C3g3cXT21hWbqND4BSZZ51pI1iSixgrSAk5g4DQMqfYJv6u1y3M4SgMPC1hAsCIgC5fw
tCf495zTyVXx6Bd8ouNmWaTZTHCLNYnSErADvM3w4NQD32dGV+EEIt+Wxpa+x9xER6l5V5YqkUoj
uAuEM4y4yXPyDpf2uN7hE0+CK/dFnUHAq335MfTSAOKdKmpelH1riLzF9B6UV6998YIQapt45Bod
8N6KJ4hPHnYXvzFDV1VoEbHsve5kqIZ4lAwQQMqWevy4maSZnR5FR/oo9oL+W9nmhTBlgJn9PyO+
qhfggUy3yxFgrq8GhqfWOWlWKTEcpPyB2IpnwR4o8NH+OOKcDnSq+yjOHFoN2rhdHk6mfGqFSTyx
c04VVtohSgn6fKCJtPAd8C3G20X5reUWPo7XlblwcRHcstdsGzNBQahWUobIKz7CAoaJANHlIj7a
5udg1bXCqzZNHSDPj/Y6xryUQcm2COc2stkkYmV68AmhhVJBXvjm2IS90JZAjnl9scSq1LnreRsD
a+9vmZzMplf5jrdnTIai1XzbFk+Xb2lv40xkgB5G53jn3SFjnpwucnOIFuqJPjnuhh9BQXEg/KdW
Alfmkk+ZpALLwZdWNMvSlx/kXCzrgfoS7O5ZwmjNJDtbFzHK3tvVUdoGoqPFbYNIu+vBpPEAoZgn
IBixtuT2SsmGqpQg5Mi6yqV+AT80+RqO6JB5bJ2bZx49JZCiFbL//1H/yNQKcxTEJDMFeD+Be5DA
FWUcKGfwxgYG44VW9iaO0qIpYCPWqB1aljOhxCZ6ML1rlwPcHxTZ6fx790iSFUYZT3FssF/ftDHQ
s/0Nzy29t1CxgkqZpLO142Q+9DYAARUlf+03KjqlAk2shB+NmHtcC8cAY3167gKBjOjSw+Jo/S2y
HLurBVYEgSIKdVGkzc6iodtnW1Pq9hztsUYllwuI8ppgwXSmfN5poFurgVxAHulGhZ4zI+4TeGz3
OaQN6iziETgEWNaYWOD3PFO0dUORNVglRUWtGPnGCOpmbY8CohEh69NGFeWSZSyDQlIRXMZ1pzgw
k9rnaRVrBbH4h1QQgt+fvo9/WCMKZyDyfiC/Lfzs3sluoghDH+YyFG+58Rf9PpSPDxZvadNLGUVi
eUQAJbrthZpJNSmIUjWHc5vKozcIaqHpS4N0RYPEVo1FAn1Ed+FqmR7hl8894IS3Hcp+s+qjcTFD
Yxu8VlIalCCKSsxwi6eLzdBYPHUMqjtjUB5RQBAF59lDmAUJ470sj7cvVM/XcxlGIl6SyV9aMghs
jBVgJa0338p4hXQgg92xDxlFVANKYFSmMgJnBQyi0lvbF4QFnDyQEJF4akLe3BRo9aYxenivBLmn
SZ/t5ZFcwpS18lCUkAWEVZ5B+AzJoMYv4gh6IjeeeXCYNNiA0XaGpptwNPC8crknBziH7sZICTY9
5xpSvyolawmd002NMmkeWRt6fK0iIE9P0lv1X7WAy9ue0mWmH3EzemCMd992E/EpZynD+4A3rxRa
QRaEKzPJtTOjHarf1c8hkTTTrMh7f6VVUWmq0u3Yh+81IllpPlwr2vCNhgSIKgG0luxc0cUJkxKk
AYwWjYAmK7XK+BJrWn7Vzkgqh5Eps1CLVpqEh/NeGZUVEP17m3Fvy4MNgcyCksRYC2ZjyzagLztc
qLUrb4Wa2hqFTa0w2P96xIxG72yN/UQ++ZLAGPFs5tdTY1T1G9PS75coC25OZ2tkzJyINNN4kAIw
rK7vVTLlKAXTxNS4JH0jl8xVa6RD7x/Z6iTaoxYZxYn5BfoDNV1P0zNno47yGWLBfOMs7ll8bvFu
gFu7DdQDeRukyMw0nr6lbzTEtDLJes3X34BMEf9Nrt8DdvglIWOlwCwrBLQ+O2vsj6TnX+SEC0Vt
VFT4i6Fs8JHi3VjFONvWdgaq3+V8ROy65yf9o2NdqpxX5vGQGfq5UYgPE2r23h5yN8ZTxQv91sIl
2JyZe0dKIv79bKNqme/z9dqY5nIJM+0iwAnZvdS2BvfkxTqZcFhoipbKYvxKdaZSY/t0pn5ZgGMP
MTB1l0awO84L3XgFveGYJbbMzK0CB0z1xRHkQ8qUt2mVKiVYEcdvfoGfEVILsgAheDv1I9RVaYPT
bIkLGF4weRWZJf4VXiqwnjvdMX5ct3N7acAo9ivcnNcpMz3KJswX158QRAnNakcLlFqxjKjXRSyG
doz8Y1tKnpg2jjSGWUb3oyf4zdtkfjXATnINhzJXyDnYtGc2vemWkfnK3J9qhHcV6gI00unAkTb3
mQElsRu/1xzsACqrvl5vvSxC7kiLm5Nj1E8xaTAuzgGO3XPVO4anEnc991DcdMAYQMBfrI/yWAsD
Ue1TlwvO5BvDQaRN9/YQxn6hwwyikBN7y94uwfIRlUSJ2V+E1vIPJIMTMcvLUKi69s9DFVPOMwld
5f1wBnB+eJQP993UM+EsUloy5WrRYZVftw8wGDT8XHnE1ZWPBm9JZtbFxpFaul8QBZBsVlZ8lID1
4fx8JxSV/mEAkBsgDHsUEkISH1K58lnQmMzPi+/QJXkwGhyEdVQ8Ohmn0h91RET+PmYR3lnJ3zsb
Ww5OJfn0YhySeorO2pT1z+TNwpUFzk0p4X4UYIaCfM+HJ5qgLNSRJ23whUNGVWAlYMj4DXWM4F0O
cV8pY4ONiing5b56j4XeCGaDfeaN4jA2+5+UgyZTXJlJn35QFn09YUcatnVWnynm4LRdRLfvXLmd
0UNYkmBchTbamomDdXY3L1tHIEMqAnR/JNyP8kARxKZE2rCIwOJ4KVg/Z/ChUQLUVW7RJuRzv4Ib
0U9fchZd2v7ssDLllk96UI+2LAqnCPXa3GJLx9HUd2xG6Uq6czvK0CJfhnX6sNVhgCqthJ0Q0Fkm
BxdwywNBCXFY20i7cYjUpuEdxftQLtCiWlJIv9eh/iHqzLVfKZ/HAHeDIl4lcqiEma4lF/3atdlk
BQuEWkdZXoyipxEQq+BrVsz7rpWUBdBMBEdaBy6bu91xDi23cO+M5HAOntkn5oz2hAJ3oU53Rm9S
wMx+ID9lUnzhsl6ziz1rb3BSmRYiUV6fej5K7yICE/u9GA3hWsVUXfLWf+oRKQZwcOse9TXKj23v
uvvOdCWfiYVHKXEo15dGAwt47hetRv0qDoc8E1bEM8bGu5eovZu1OdgFEhm6az8CjuuyGc6DkFze
S1YBehD//TEmS7b9JaMnwyBxV4UJJskEQ5cD1GeZDrZ55wI7FXtM4SuylW9Ne9exrmqk9jOvzZQ/
n6ZfCliJ3H41i3JFa9ItRYVmCI3vZ9sE7e+vl530Bs9Gq0MPr/5kFOjUEtIQKdDW+N2JDSj+b3JL
dQbpE2M/1lGHv7CO/gofSNqAqkZBpjKp0FIGha0hL4UBStaMCDWs2gQmVUnBifKR+tDnLB4aw4qJ
Ijfdswopsm8gy16fBEgiCrKCjsf48Qx0GG3CGkbVz2m84hC0Vv/hcEonvtjPDh2dPJYTuuAGPQ3f
MhxI8QyfPpkNfNTVN7X+m9AP/h0oPBYn0JJMAFliNmJQxbNCXVB8HcjTVxNYmyo/J6t0zODQcYyo
gPstc8/et0T9vtieu1h+QCQnxJli28sCWwsgDLGhzcKenVJgyNARHaRC02XbchpV3QupauWtsOto
Rw5sPykI5eygpSROrR4m3LkCpuypRVIc/s5Yf+l2b8VkZlXU9uP6v1aOP+Tnm7RiFuLwr16xUQq0
NHjFJwcTlE8LPdD6RbIPvaoLIzxtsoMvw1VG4DwSy8/uEXpI4uq2b1gbKKGAQC09+b/bNdi1lai9
OSOznvgh7BCQr7mHbJ1jJI6mwF9jY6WmixuXpoQsqHNsK7n/84f1J3lwZpWVe+6IgdTMxaQ7pfCc
O6c11KGSthpvulClv35FYWhe4QdqadWvhOum24BKXgxVsAxtLKC5zZX4QPrMd32EqTZE6RqZ8c7H
1Fk1lWf0SLDrpGtOqYVnOlvXSK7GyregaQPl1qmEamMwugH7e8YUcqlYMNtTOGcm492DpWb2m4nN
fc67khhO0atD1A1IgF3gm3iHp0vG3kttX79Pcb1GLemcLDRjW3elLN3SMgZgtGQDh1Ahef2tjsdK
WmEZSk6m51DBspByL4KUhClRYqNj0OcgyOz48crsCVI4akB8jZkq+b5uW3xFj9Er/MOqUil6FgXn
FC9dowr94TLeLjDp/nO4n0lBgwUJb6hkaIgainPkfDHcIhilIsFqv2tv3ERYcFVgLDIfoAF/Qd2I
LB8KHNL5/0zGBHU5WUnnBvPQ5nYqjWiAA1ieho2W2OatNEj/5AMYKjqulRYxeCUXmhuxqvj9nPMq
hYpgnslQutLzJsslPO5MHA5ANvJ7q20JSSfvJgGwO41ivM8fIqyg1isYnkJA/1D2GEgoo0mSChvY
8a704DQ7c9Tsv7OUYvuhqJgZmLfRCv5ibBo3qXHO8/9cpV5KDN0JEPQrq13utZTxVPy1+GoGfQPl
LCHFBfib+Am0gpyOZ96zlL4bW11NhAOEUk/uKonTrzV09drxKHS7RHx6qqbeIdmr94vzUmaEY/vo
r96lbGyimDU7yea0tuxaFLVe+t+AmZ4Im2Oq6T6d8vnegkI8n23JJzQY+bPagWyeov96YqASLKX6
ROMxE4KS518qv9ShatRjAPxThas+YNAnrrlxc74IOfTIcTlFiY5CsrUTuy07ZbZJLCDyPcLdMzOi
kJE6DWOI5p/9S/SVsmJbGDMe76CH9B3dZzmTXXlUFv4uWTZcdMuxW/jMD9eG0Nq/7udfeFY7BhsT
VLEDjaDLr4FEUUKdquntCL68KlWKPqYwPfLuINY5qoMJj+pZybx7wF/2zVjcQQ7z3BIxQfHYAGAb
04Pfzk66fFp35I/ArWYK2VtqISAAZqkqvr+nB14HuQrmdY+emX1INpl5R2/LDpbBDgoj+K82L+MI
rMKh0fThfyAVKuodGIPkVj8Rnv8werR+zA31VheKId+tmqxztRmR6CPSZK0lP6FtwUPGcL/1LdDf
yeqNgBG27k5rdm/lzqKka0YW4m+gZAOee6gnPqOL2kveLCXLS7SXNz1k/v3q51KOVvH0wn702HjC
WHPnkk3tB7j3CSiASWiZd0lJq7wg3bWii10hxA064l3XzSTpNcOYkwZ/KynX1ZgKUlxuyPz+q58Y
KVex6nLpvWV8nCfeXdgZPwtnOECSWqNfv4vmUlrNKZiMR9btqcY1BIolvI770Sqw2nbtnzZOEbZo
CXADiXPS4S1cLx5oc5YMk/wzzcNwoIrNfaxdmGzeSwyunLFodaoUT5ijQXF7nZTOJfpEF9RPfvRa
6CMxkoCBCq6YURWF0s+ORIZH7y7S2IKT2cyKrcgUO6xICrahINQfwAUQMibw1wHZh6aOBPiEZ+lw
6ykZtnCdq92J5mYGrzONo5mm2TL7vctEKhRlfKG9TRS103RVRc1tvykGyhoFpRFdIXhgMFVuf+ne
GZjHK2PkNQR0pwznGOW/u3kXGB1IWwENLZLlmXDQMYggEhtrG2xqZ4Ut7185kxW3TnmEgdmqvajF
zHuAglTbWvkYIVzGklnX7R+hWM3hO74mdadbn48RVJQVKczMPRtNSc+i45FsRoLv6f/Gy7nhiZRH
6/c5xBbkAJWvJLreb1JyaRH3TOz6uUlm6/ZgNup1YNBTdAV5isdy99TumKp2O1cAxraSxQPRlnUA
aT0jT5t6cfazF4rY9eavDz/2nuwe8DILEK/o5aT2HGXQ88RgU9fZhg+eZyPQahhvoUwtMjaZLlcx
of+tX0Cskh0ClXnCYo/V8c2CR0khZwGTpANXwuNbNXCh9iMi1wmaB0os9FO7KkpIXhY6xPF0umGH
VaKLlj4GhI6cXWjwJgXV+UVwuUv4OlChFFhSd9xSNLrj0qF3Sk2vBVbOH0ZV7GEB1Xp51C5RDbDL
P6QJ9jgNj7Ej93irty5m6/jf6Sk1CsipccK0Mt1IfolUmNp2wiorv3Po/4mJCKvTYSkk+iaSileK
eM3R3LtlKTdENb3Q2TJ7rIvBOukF4Wy1OGIBryP3PO56QBp52i5QkRNLRBU9iAZWUsAmRLPDeT8M
5plDbNESH8Wl9EzpcdERB6iOdxUhyUaARTuq7h+l8dQ+Mk+b9D6e/GM1RuUwx7f9rGhUfHe06j/6
oIwGf9jm9ZMlYKUuMDM/93HPFdM17xTjOgudxKLusN7OATyTJBVaD2dSMKF3ZIWDTD9+JImJxVVz
VVeiXWsgyUqqqfNRBg25unj5/3UdqVRQauOemjGZTHJBiL8zNpoZ1LtMy+zIEiF45aICloRS+Rdy
l2DcQEy/1P/uxsEPMrCe6wn+r8pIX53FSAgJoDl87jBOrlKhKonr+iq2mvFGtWl1w8NM3pArrPYh
g4dwdYEFE/JD2slD/ksmOuNI0/NSnVJLQCf/S8SO1In/iOwtvXnKgaBFs5CsMOEvAvJlDDoy7pcf
3x33nd5wxfuCebKeRCxyXJvuxS4kqYrJiVK9+/codf8Bran/mKVsW76ehPKmWXznq0MaeoY2SxsX
vD6Lbj9ykgSLxkc+5+P4yyfXq2Sq1Rr/IpPgW9v5rLtfWfsbhfcSRmJhpCPcaMtlbOIVch+kLTaw
xIaFEdK91SkYHHOq30E+U8LkDi81vTS0ojtSihd7JFxT6PBsXCeLgSHstYzMI9bTCzPHhhLLsEVI
9qUOGUkvF2zJB7DTk/kggDA1l23Enb9P9RnzEgH6fyNNJihOhwhBnJIWP9Gl1GXwgpQFFzwUScDJ
fOSwdaO6eMgXOVcL5HgTzA5f/+YPOXptZ+UBK7a36CRNqU52AquDsZjN/2SBXBNv4IWcSLUnZDOR
oqeD2oqB4M9E8PjWiL8B+RMprmRCya+JpH/XVRQngdxL02ImFXzlcKtVa9sRCUJUUDyJ8C/MRW+i
VFmX0cilVkWjCPzXXhpZefeLt7b06yfjZsuHEWQe0kcSUuTtu5offXG7gEjaSIk6cQOsawFdnKfS
h/9cJwXj+U0G85BgAzyfPouJBrQZo8bFCDotNeVJQfaZGlrsQQV7WnKhjTAT7G8x4M6U/7YI8mGR
NYMd0vkpCL+XUTuALX6Gzp1PAfNOnHy9i6FHvo1R1W2nQWt0jHG5ezPJYG81sTEFWKE2Acixiu1E
iomCrN1i4gcaZyQV3mWFtO7DBSw2rU0RQgT+RWGl6ytcQFDdpIhhwr8EGq64103R4NLWV+jh3DXG
dhSxxMPnufZfG2KaXAdmN4f01KlglX92u/a5hCUKqtXYY1by2APHuxUXHQsdSqUVk5HBRIio0ISe
d6o1EAYLWFpsgrddw36QQ1e/OcQjcODwzoKhMJp7mmrrOgjeM4V1icGrDus5z89ckeOcIdO3SMmn
rtJgvw8UCiuWFC3hhc+jX+d2SGeShPlvw3Me51Dd4i9kV3XYQ19hYmKDG9n5IFzeK1rS2sGEuFyH
qMi6mIP88iRSwJU0hAGJ0LoQ4+fyMzLcjtnipwrtUzWsapVhraVONvyDndLg8dcUgDZ2lU1yoJ2+
EFZFIKs0vv2o0swTUvdUbgmb7USj6HA4yOu7qmXvSL8L8FTInAKpyxfrMjvg75LGhPpJpkNo/KsS
DqhJ+YAtL/6nAbmNRw4qp8NoUzdlk90yOOzoA8UhIYLUutjOzuPj/stdJiNXnPNdO5SrTSKz1TDS
L4NsXtRtngqvgxD3is3wFjq1UJYvkjZEAG12FcWkY3iGiXKNh3ep17v+fAIzvW+IEvLX6N3R0i+/
FFZKaLiX7VVEWKLmlMgj6dTB6GbrBSssYN1fK6F/2xoXfv3m6IsmoLHCQgjp+fLG7mo52lAUwzq5
0VP+hwe7QN7FJavRELIp/ewdifmfcdJwmvzlpBWBNQFpqbMt/k8BTL0UvACXt1YyIlgkX1Wm3qdt
EnXGLysf1J9VL0+32GX8Hi9S7eV2YL5RRau1Z4H3mTMvXnEJgoQ7htr3xlgRrUyjr4rsxvQlIKBc
PQHiHSSeNVoDQqOIz4J2DpoCErGP9sBJjNp9mrJNNRYQ0VHd499VFY+nAKxi2WPFBTZBDfcYHcME
3IMlaiX8tWvTbwGrRrXLtkALFkWay44YmqpfAxEtRsAiK6fktRYYx38TuYfnCbGsitKzrUxBGfvs
2QdV84/AaOeT7bnNpGVgONbpUiPkIBn97M6NMUl3WBKv+wK1Pmeeywj5Easac5qrDR5JUiNDLHlI
ohcT68h2jrx1MVvUIXAmrGt97y9TBTfQot6Rs/0sVx9m04NXcjLhN5HUtRMCYSlEgMRh5C1uCyOb
qf3Ns6czyhVluUR3Y8n1AUqUms7vfFiVkM0ST1YxlSnKZ5cZ30HwIGE8lzplckIP8RAq3MmvVuNJ
YB2HcvkETKQCQBTaRj/nis3EYAENNDThTOp9rzVJ9c6dlPpddr9PO9ptifACKs9xx7ZbrTUzMtXa
9Y22SJTq1wICD/5/0xVmQN/Nr7eKYQ6fovADy3yHk3BfGBlUdASs4t5owHrJdCjBLUB+e57WeJQl
Tcrt3nXPuLEg9xohJSpLhmWAzyvmoBZxAQlHHlj+DQq58u0KRkg4Sp+3qfQsU2N03XsjOGqVYhoW
OyEa8xo7tzXOV9sx/ErQznZq1aIJssB5MXtzek8CkPaCaNyDTCICWvjNuQ1KtsTGv2T89lk23W+T
yRc70fkB4BteSeOfag2sahmFLp/HOCCjgpUvazBjm4MZHzahU0ZYCb/Gpmz0BUzcbrikEJCXXz+9
KVHMGCrw6+8Cik+KxKOU0a4TJikTA8FCeOkzwfY3KYb4DQNTpdMPy9vH+IuElLwlXJFJ9DXIEn9B
ad9tmBaVEgF1nace0miiEnz6A+jb9AgWd5uv1HeYaXIrISj4/BAFKqxse/hRDinB+XvTkn8UK2aj
/FwtRdMI0JbH0kil25ySjisf5/Hr/MVMXXJ/BOYTnzbkuDs2mv9dTQVHnJMG5bK2gU0qhj9tpWY+
Hn/2kjxlVyfZTDj8v14750wsoYgsnEa8npzIIDQCrPVZ61n8aUYPPmpUK64h1RygLX65cpJ3nVCY
jm7vKoGQ7X+7bHPuycbRQIHN/jJncWtg29tX7js06JdNwTcGxJN8j3ibavrZSa7e8OtWXJqb0+9Q
arrzs+xo/K9TtMi8cTALRzqoudQsZ/4AWnbXv/Eb+ycYuDUkAR7G9i4tyWfJpB4Mwrn3S68owC8g
QrOTWTAdbvWkQezgsyhNqvsMH9TVwX/Kcjs1yLuSNXUm7MMats8bgdgQGQEu8ahN8CeKZwBo9+3L
q7E4cn4kwhQoM2zN/A8fL8YzrMMSYrpX/dJoaNSP3tTGDlkxPPJS3B11SxkvZxCY0O4Dzh3VnPyV
wQJ9ZKgWyVi1iH4i+vnAEgkExmCZMhRqfR+kMPl6LWjKbAjyAJMOfjxgqpIwewowOn50ehTZwiTX
mkpRqMIkVW8SYx1odJc2XUzmzpNqE0732bETaUSc7MzA/I5IFj1Nom11H45bulZ6ygQzkBOig0Kh
KfBOZMFsyT6qYhrobeOaDTyGxLVAM2nAu3gxQ094Pu5cOJznzKfw5teqshxPtne0fnwbVYPQdzlq
CHnnOc8AILAciJQ9ymJX3C3fj5SUAJAgvxBL+ujXFTWOGDKj2QR2RiGccB5wYxrPMfvMTWrpeedX
u1ammQJqqDaJ7FO75C5VuX+5w8q4vNgonVy8BjOWsDNUHMHpksn4bgVuVo4jVk09HhdzqeiBlX/T
vBVgcWpPfXfIRlFak7HybsaqaTyC0K7FDDhcT0VUKlgmxCr08SIomG4YpvCWH3Tcfkv5dcluZR67
BFxa7oCSKZUtweO1JP+RyHAmBAXMqK1NjPZPoVgno3TcFMfP28RhoaGt0dMCUzlmGi4NRrJi3GBE
iV8410UVu6+qByU6CBme2z2G7k3q+F0bnmTbmpgyNN5hypQ45nvkFroK6NfmdksbHwsHJJJ1nZuu
6jY7OoNy4mr/SAicCGcJ898rktjzzIclqA6otQ6N48WQ0FLdGrWL/nXl+UVT+OLDJphYolJffKqP
otqvailPMs7RyEICP4W3YyekTzJ6zHBvjadxQYQz5uP1xPr0xSWKQxRSD/zsW8uDQsJxULRxKir0
ElifpNn8c9aype5Oc3sX6I3Np1cdakzJsvN/p3AgVG2+WBMYPMfTzHPN2xkveflRGsgMHM/xJh8O
mYuDIXwKNvRdG0TG9AduIJcKxZqwlumkzQ14xl2LRgamZQFhefjKotXTFac8UgiTIIjajNl56pbt
392etOKwRuXjcb4pBRcmmpOKFT0WEOupm75oZ54oKKo1hJ6IkyYGtY4RroTIhz0VUy6QDc/7ZBzA
0CF713V9/OJ82nmZfm0hS6UZ5P+VMD5OjHjgxnPcAJDP9izmc2wIkGeeh86H7oz8XiETMqo7ueXi
lTjB2vjlg4Kq1kzMozCC2p6uEQsadw11dobrf9mTi5sZuTztKZmigjYds8sKOD7gMw8W8vyJGiHz
KaU05h2lA5Axn/423NQZlUaGW+xoeZPnWZO3r7tsosjltQqA7Om+pLdpDlBq5LPqzVIRVYRW7vx1
y9dDMwaCfrZu9TN7H98cZ4P3zH1LT4N0Z3S04WaLi9FmbgxInjlSM2Rr+Pn0T3evQIBGTUmM37un
JUhfbAo4+7YGvoAzh2DL0o3xBkgpbl2cIuOlF/I6uVL7FbwjctjjldxCQz+JfMqKH+auGNZyHMzs
lwjpv92z2p0pUNof1DrN8ue3GOSbq1vmuLvCHWASpCx80cFZsOwa0JH9RBq9sRdHw5aI1nEtFzXm
7iWCfxqOAj227EEy62UxOpecLtsB6ipx53crKSd8s92mshBx1Q0sGeGHbN6mLb+tg3pxoQ/Ef3fl
3bysWJl7OZBAL15XtZhqmNS5DRRsTdcO1bKlcK60PfFQFJA8185DCMygC2sA7vytmGVMKUgpLh3l
qIORGYGrGfVQHdwuF5hL/ouJQG0Wr1k/6zJKdnec1TXYv+kxCaQFzVZXeNR/Dt26zh1NumuAWJ9T
lGU4WvlkuE8P3BFYag472PF90PCfQzLAM6xkMuMePisV5Zby4BIa/IrexptRpnWcvNjNs/0ASUW1
wJwUagBcHp+2w3YMjKnbnR+WI7IUdftF0h06i1U6psTuejZSlV4UM8odsZVb6gyTiTuGB2FgaVZn
E+tdrA2rFx7O2SXdALuO8BIwrM2HC+um5LLaA/eu2Zn22BpcU23uCdBBbfyE57/hetkE4sbe44OR
sQzDTOsO1BisHqEUjigAMZA/iHYy88gfs0Vo7IyZj7e8H126XxyXEF1kvKbqbPXgfST3L66Nmn7H
/pkneyfnI4m9yXgQImdB6MUZsollNdL/MU3iGuULiJ+vtopvfkg415rWW1Hqi83gDf3Qv0RHlZQl
jIHA2jB6gxkOJXzMMIstAxJEp5rS5dONzxdSrdK7Wim+9/pnPwaari/qErJbMfcBlEQYTSuInGIC
yi2TD6BT4LVE96+Vy5yFatA/EfuwDbunaf62JWbMc8zS4ZtELV0zsxds/TuAVXPd2b8x7RpyuOpi
BvH1uYDdWMdYZiLjHwz9VYepAX1dMOhZ+USlbbklSMMNfMgpsDDurEakMppW+O5xtVHmCpE9FwKS
lrNKMJE7EbH2fb5T02N6wy3SYyDlQ+yXBkGTXfalr1ejhvPyhyUqDNiIQCEl8RGcDFUDHEHnSIGI
tt1EoSBUePDeEE1ICRCkJt8smc692DZmfnYeQ81cawv6bXK5aPZFF6f0LCMFcdvhnHT2UcYoTSOn
RecqjhK4GDPYCKveKF7dIq5lBJhU9SUvWG7EtA0Yhxd/Oa0RYPlRocIaxKQ945xUYgyjTrktuGGk
jU3Yr2xnK95OuBcJsul2BPcG/Zo/652PluIbwKiz+E2AIWSN4LVFPmzybYk3R02Ql697lH52l1Bk
GtLV5lNACNHOtLQf60ezwRyCEGkr9yeTVDd0Wq4R8X2YP5kyWYj+rPdUSXiinLPxvEoIqQWYGtdD
SHzRvUGJgFcnCJwz6mH7cjH8VevJl0sg2cLW70RLBDQqCzPzwvSpbKQF+n1On6mejIn68A0QU+WD
iVladkVeZhj27hhYM27DNp1sZiPmY45UUJwIQALzRtxiiFYF0jb/3fH8pcqgeo544z86BrQMtqgM
ltTPYQRCZEY0S5J7e2gzURxe3p7qyg5tBJRSTW4lcVmkWaYJVClXo9nelnNXhv3UjMBKKwoOkn99
Q71Q44NukWftUIuILAIWeu9ocXtYz80a/z8gKvRqPnfQHvWGhYuYxSeqMWDGMHvwCGypoFnoYghv
fPUr+YVarOMQI2zE9XkjZQKSnUnLCzNuxqNpBGLUc6XhUQxHTeVagkg/DnlQhONy04b8AtfoWYpL
5bfUXPppfR8Qc4wJCZW5FUi5e38tnjQ/VN5M83kp1e3fwY6B3/94Wrfbw0N9nq6YV94lZWkIq4X0
yDP3Q/Z+bPz28Z3m0IfYKT7bMPiFjIS0ndKM/cHjvVNQNNhcjifVO3Efnjy7LWbnxHGz+w6EN3pX
LMQZCsQRiwDgUd+fTweNkGzj01Cr32EQ1lHSZnxDqcVE6DcHIbMSAHzLFtEiwyx8YIy0pP8DInA9
sLBddRWQq65eUOT5TTKrDoDzzjCZkxfgkYD+1MHRs9b3D8v8X6FD9FG6xrAfUqyhEAA2nDBOVRvh
r1PEuLYQ7/L9PLdOSvloGZYymDGgf/8oo0u+sD3n9lV38jnII2iLnKyVwkPt6pjlkKl6jGoieJHQ
QynLT666JqV8wCGBQWrQDvo2qRqwk9WOdQiebj2UHdsDtP60BUj+R3OmhgVhoMkfuZkA1tQ+GqPT
xAFEHNPaVhM6rriQepSDBNIvcfb/lPf8xRN80FKN808qF0Ty1eIlGJwjMeQ/YdWr56EDNx1nY9AN
nn555Ix2+58QPfAwpc+xRnTG+cH8gVp7AhySP7D5BhvIzXA8NbvJuFt1sL09HYWWhUd9oDxIhHL9
3op2ybrdt+LNDHvstkDd7tH9T0KArHOtDF1R78cZw1E3bwlQQrTbnEDsqNSMOodBWMeH3JWvA3yl
XUlrmskyh9ZomFyPCtllzqjU0mF9RAfszUxXe49NbagrCisgYxqXWH7W4ZozvmaZMjhN9Q7sHQcI
ReHUXwlzDD2FNYr98DxSotyR/Xx+Ips09/Oqh+fD7bqE9OJ5x1nRrhrLmMtMm5l3GJNP9mFvXt4e
/UvFcIt6Yu1e6HhqraMKjAFgo/pesKh1jneLpPInEPPE/I/HXQbUQ2GRV7C+ydZgkAgLennr6OcK
mWzgBMRPsbM6H7xFTgAqgrDYQ+50c7kgveKnnB0MKOCsDBkiNQ7PICHhbjsd7q+OapvDXLmU8cJj
k618soUPO6+ZSRAppw4nq0FIWd+9gzGDF8v5ndyBjmwuV/J2rvPGZYhjeR4X/cRyZ/b+VkafFkwA
hiNwOZF59GUg8TJnu5rynPc8bwuxwG2yeVyV+DTV8a85lkYCwyH5qVm+TaKlqwvktmsAZjtH+2NM
2IjmXk0HfZnZLixaybPK6DJsAERTgFxLrgliLAGVhhgvjFW3MIi68V+0BVSBZQQEFUcoxIyVg7oN
3hLBgW3ZeCFVe/id+B7u7uX2Kks7P79elQV0mB6zbkYQEW7yNwkzqzaEnQCYulXaNkUWfUaNGEkZ
C/VDyFYCxod6lyRD2E/+DLK57CXCcDnesIQ5wKw/Tb3V08xTJzh73aqoxmzb7TTPrLA9HPav8Orm
jeGAwK5ASkCV2i0fUIzCiM781ffJuVUZq/gefgQJxaO+Wq8MXgW+ZxzgcG4I8GWg6qLN3PIGmPDT
C+/FshidPCyZbyiOKwzm1JabdrXVPfftjpHKHPg+s+STcrd20D1uPpGG5l/lcsO775JTo0zzb4ek
+WxVxox9F7VIRBfHX+peNBbqXhBQVrK2ecg7O5hBBiDyCMJai/ks3MVBMb4QpS1dYbfenWL7A8DG
52+gf8cZZAdNyr3IaPfjdFS29afF8qcoa3uForUpXe4ZM7D+YIEWdgWDdG9Hb+9vg56P1evtXydu
bcAig3CedYfo8eBY9WT4rKY82Pvlq5WVTYgyFMQAEy4RTDg7c9AUs7Ri55rek24t7yx4fXo8xlEj
umFENgqVreXwK8SiogZQ4uxE47kjTnxWBPe1LGZFmgWxHdpfe7W0hTaoDBzhp51JkeUqtDod96uV
FwRUsMeFLMVXk5qFVkrxAzuIDNn42Egw/j+MSrby1WekVYRDwJY6/I+4kf+aj7eZOIzA33WC9a3i
fe21arKcbDaydc067XgU0ZqrLY1NR3JuYzADqPA/7pS9e2zTAejm3cGlxA3A7/TA+rgDywWUwtUq
AxuClb9G5P+qPO9RbQxusc4Xc//a0gmnQPELvNn7weGjfYfjD60iuiN6w7zdp8AVI7V1bAa/vpg9
pPpPz4qctXHNcz1PyVxxwT48NAWC8AyBAGSVxT562c4Xj3hDlPh6J4u0tce1fIf3Z9R82ReT70UK
P4gBIMokwBkjEJZ3Z+x2ynnoCAHgnQPjb3/V0ufnZ9aH5Z3qh2WFW64lkVppWC4o5GlpPRlC/3/I
8vXsOYiFmS5dsE/0szH54w9fB/FWsf3tna+dcO/5u/+0eTU/vbaInWS7OFpKemHNotySOewjK1T7
toztrj5jVBosLIPl7E0meKo7LkDpfEVttn4N7V6fGC5CJ7Frupr0oCm8Pee+fksM37r8U5xZRnXa
sBClUAyeQlWWCJOecoXU+aoiUadNaoPLbIpR7v7hLAA2bcvjSsnuaWSIhprsuMxvddCpbO0tn/qf
2K88RwHO67P/gDggL7VemynR8VRjjrPUV5kPv3D5vSwkQ95xjerNyVhXPPt0aL9q6ZX7yQ/FClDJ
QSNkYwnZJ2pTHryuBet4SqXzTcVcPWtBqqUx0aOytHdbTUnDypV2Q7Faq//mGaz1jbmZMQTYrTUB
FwIZTCX9M4dqSKcTnBoiCCJSUOx8CSKaH4Yxy/srSnB4Cl0s2z0LvqEx7lEBsextDIqG3duh4XFA
ZihS5tWC/wMyK0rf1eELHIJdEAnPJurUK6HEDma9jw1Pea9DGY8TWaX4K81uwsuxaaalneLHFLt4
IvijEgGv7jmqd7vi3jQt0hu5S6wehmGodrHvUOyjfx3jBVLqKQnEUwSaqsjQ5fottFqRLkEG9R2k
YiM2QFyZ1VvJiWbR2k4UFep9EMBZb8PDaReN53Utd4dYinmKOGjZAL9a0T9uIZtx+0wZRE9XQtw4
Xd5uWG8AnUPBxbjsODhONNHEhX8AsCXBEA5tpFpnHuBTGuYdItLTor0Ai0wwaLBdguifpDMyMmX4
d5jTDBNZadXJOtHzi4wBLY/HWsxEn1f/dnqjhb32euBYht+5/ZMAsNIoRp4tzQ50b10qnlJTmov9
WoIYNTonmV6F8xIkqv7BEnvfRUeQNvFFY7ih9xCFQpBkkugKSpoP8E+UdY/thFYLgx5MkHrzkW5p
RY46qhI3iNLt9lr+xb52ANFoM80B6aAdYjGJ4apJHbpHz+Iu4XTtZNkx3GdF4K6CCsJBOKdDF1qJ
k+uHNiAK3vE+04DLXk34mjwgpt2UOEGSAdWLmTMgMX1tte8VbQO3Jn6movA5JR0cyKITMae0chfg
1SEWPV8SQpua/fANjkp9Ez0EEkW932PfSYm4Hnjz1Q+4rZHravL9nrq0zsmj2pRIx7qunzdluko9
IxaNGnu/9ZcDwMiceIL1RgZP8sz0XdiP4Ddawgxa3E/VCqyjlN5nmKejIqJF+AG3iERW4A80zzxK
dAfSpONBWcslyqRdojTNhC0PX3BF00fWHOl6giKi138SZrNtf72+gccAEB/fzr/z68E1A4YtOORO
79lTbTh9v6z+s2NFa1SC2EXH2PUXb/bPUUnJ6nLCgJhWPu6JRZ/PVPXKgrricaH3cGLQ5cf8tUnN
s24NV41Avd3ORQGQtrWQAp6DnZMK5prGds2Kl8QOVk49LS8VD8pLlvwW4XPhvh2bhFmzCGqf/KvW
wyFo9nruGHQWP6HrY2UkNAERssnHKcsOkIODD/6Sv3nPyZluHrDTtnqEeVgdmz8KGXfCsUt5tQkk
a4y47Pcgp0zXFN0ouEqLfOWzxm9zFZR1b2cP2AjYc3Ub529ptpw9jQ6SDsVUzbwPX0GAsQSj/gVd
SzjzSxTLCuc+0FVhTrQs5y1uhN0biL4T8V173Ap/OzBq5Bboo9I49BHKm0PatVHbtw6mDAw+oPhq
ehbsd+Zee4iQm3BzOKTAex7jLsrDvhVdPQb59eVYH81+sh1jVmZD7BTkxuU7k7sakklsaAQhWD33
n+oG4HnBmb0O/+7Kjw3Do96baJL/77QxOv/rc0LbPaDShtqAzz5AtnbzdzbHiztfwqE/XqAcwuXg
2NYARC4+WQQqCOpgD6XQY/kKI71I/pMfW2nhSTScrBAZfKqOoTeiewKapIQ0gC9itsjg/pGTUMrd
oWu2/vKL6ZaHq3UQr6N55NGz/50HA76hnrBcPSfZ6zGkBaZeVke1lKcU0lWoODsTodSTpsFCJQm6
bj8lR62afeUwjoGleQG9Y7txwvEIt9JueYKZmDMRh4QbvVmffKS/m1WLUH0F1rXjt1E34c12hcSu
t8u5cu8hL3JIzvVASOYdFhn0FQ+JqUBsVWKwofC84o88ghyenyqkI7RKC9nqz/27i0UrMbl0lOs3
M9xJy2Podt7YQtDAZazb0cT09U0DJ703dr4eqQK3mZYe0Rt/QJ2QF/mHoeanuwT4YcZ6/MavZGDf
V/CWvU64U4zwq7SILhEpsz01y2CZW4F9KdsuAZbgJZZm/haVrINpL+5WOrLUyXVOvugjTvwHLvwN
eo2bCVECA69DcNLqkZNrilVBZRjOM4b3lHjie5UmQZS4cUGkGOQeMnlZukRo7HYMSnij1tzOu07Q
B8yley/X29iTVHJKrVd3njkoss4hdql/fbs3M4ePEY3quvMBAhxvfhMHvcSDoG4Tc1QQs6v7r4VH
CnqjXOJ43mHYIwliPDpa74T21ac5S02I2bzbADqKv1E8koU9jREyQ0CiDtLHNOAYbECQXbIgU0R6
MO8mVM1JG2OtGDnfropq3gj0bBK++GqrA9EAqYaBG6M2XSpWJgryKbQ5KEmLHQXwkQbgDHhDBz03
VCKKORqsoy2vDVmcDVREEQLtDPLtsSGLQYSSCFQ36+AFNzdw/mZCrp99xdhtHd7YyXvux3rYJ8K6
cgIyaVJ/RgBVDLDmoIgtlnUCDdGLDvDeoYyAYP1pKO8RCMwz2Jgf9JUkxC35HYanEc6fTJ4W2mI1
QEJcchndLkPDi2tgDjsm8Ez2a+O7N/drfrLpvdKiWeb8cCSD7ubcouhDbOpRtb2LdOm0qvvpGRv5
2g+J9W0NBaj+HTRKsWJXBwDqg9yPfYGt70mIic7r0iwqvNv45kuKKlpRvsi0CNWxLrpl158Wg1RB
HTD/aFWTe1ia9f64v6c7odfu7t+8zwI/xGqotTRpBWNFtwm0VWGTYb8j+VM4W0nxErIxQXjKxICV
qboFEXZTX9c+tCSGzXY1C+vZlgyrjkj9MSpoTz2v+UwvCNGhOTjs5oIIuZXfE1BpmPiRdviSZ6Ak
ricUlpIHNMYRmXDX1v24VaycLaqj62tzo2VaDQroml6PNZWRgEiYzOgKohVjGRCc2jWrHs2vC5K2
Djfe8JQB/CtFDbnu1MEypWhOahKu3pjw5GqsKsLvuJy3WjKWREBMSwh38uTGyhf41p7/9raTriDW
KPy0H66VProMiNCFFbCFMMuUtgZASIeUr12+otIxGXkViM710kHpanoCOTWRtuvrOoOc/faEkFmt
K/dpvZX50B9PLl5H41IDVxcv+NloVZDJ44mmtnWlsdDQasEP4dskezyZMvUM+nCCZWtybKk0Pgn3
zOamENn9HT+jwh4+HYewWxPe8SFfkIc+teBTTluz/H4uWkdp3Zmc4G6QBGdwTJVLdU5KAk7NCigT
HTpg2yidwsjZYOMgJR8Or1/Q2s3XfkmGJ3UgF2AHP5L+t6uy+/9YWesEGvysV53bPM278bf3mE39
hF1Bx6Kp72njRLyXWltTi/QA+Gii996idoAPR7QmVs+EsbfZamaTz5rdkbn5YI+qzCcuKn2/g2VT
sbj1gcHwybcgAvo86nZGLu3CZ42VOlvPHqu2JvpklqDATWzv+pxNHubbyVnYYDUzvsBlcOkPllRO
h4OcO13bqS9H2Nmpeh1GZx+NK01HFCKDaD+Qc5+I3UPLRZbF+g61YBiwBrC4rlNk7fuUTNRO92T+
wfYhiakdPE44dlOALQEpx9MNgnSYwuT1MYWOQa4B1QTCTa1S5Ga7ZzLfE8/DKhVGLU0iGUy5e6JL
SybC3JfcsRvbAD8uwGAH2ocOcVxdPJn49IruhXnb4Pf/US8615dHmrR2HiaFSnWqkbR5G5YHEuI9
SH+SQnKSl8QE+0JGorT/NZv0/yfWf5ccbnpAsRt1soK07cVp0Y3CBJYgMspdkV9tpoETVKvO0BHV
IqRUd+s8y0B5x9cCsS6ouBGJXLocGn5QpBqrMoMHcrdRSsIsocug2aFp6Fu+O2+3bKSpVNA3t/6W
7dVrBQxGgr+zd7kD2Ol4ekkZdq3X70aHh3sopXa6LBAQde8zc6Q/NtRwgFCaXa2xVebMPCcNGkgU
gUQ3F5rkPX4UkuAeUXSQugjJDDjnpT6GjhrcfCP6KksjuVsKoxQ57zjKbkUK2l1vSyQxBs3UkYjL
rNc+Z1Yeu3jTo5wWylvWfYoi/vhFWrLXB5qRrtE/JU7xkuz+gpTLppkBD2fFVohziya3Mx+jVeFG
rLCiLL+jFtd/VUqtnx0EZcNA0Tcb/vvK29qS9OSyl6pPEA10mlENyKezf/D454bQ0/x5i0sJ7k40
uFt7pqcTHQ25mM+fGHDdQi9zdNSgMdgHt9RzkZpYZcfqfI8U9rJxSDv7llfZFjfuydt/NcdC0VbQ
m1XS0F8AefH2y2r+S5/osj88bKPquKTEFQ7lUFvMpJiuYJo6x7axIxlyqN0QtGjxsV9trNMy0I5g
dSnFg9wMc7y4D8OrtbiVpRkMCqDF0SRmR4ZTpst2B8quV+rRvrme480fdOKtXdaVWhH+9jQMslHX
ijaB7abH/ktO20Dih7ObebIfYw4HvV8a3fI71oJioU3jo3sK9F6fjrrlh1w5qqrKmqQLiWGBXvG8
thON3R/BHHH2jbytTLeuMUnC3cA0M9fKADQ5f7gXW3MHaPrJsXZSPeEQO6bl6wvQC8tU24/1Tc9p
GAACnlBBKnysMFuCLQrj409ZddpAeHrOirNzcQ+kRkJo01+H2Bf5cr2cWNAgO7deSOHnTTDx963O
O/vZCs94qXrTlMx+D9AeM+DN7a8k0G28fzN14fUDlw840v6WOXpicVXiGAypToRa3s0HmDmQO9SL
IvC4f0vJs6V86nCm1wMpnA/DSGqwL6yv+fTaH50alcWH4PN1+45T29J21el5BsG5WokzVMy71XTz
m/50Umlxb1I5kY3YyHki15fz59O/USWVMv4iA4dn7qmos6W+CC+PW3xLTm6IJtRaRklQipSbKoeg
ZvBknAu97USvBRm5KCF7EX8AQjzTViuHzSccS9eR2P4lSulP/QEL/Eu+DU6BB5WcQnc1/4EcY/pv
XXBpqeWegMcHttXYRKZY+9UnE3CNuWShZjBNmAs9/JCa2Z9Z1h5h6S0zunwqYr6M+qAVepZbkw9A
Gx1jiIVkmpMTEZeysEnbMpCv+Fq220ike5cRRAtpeyNVw/Rt7kvbVE0e9ld/WYBnQgmTbDPbStN3
/5LGZT4+ig/x7VYud5SJ+haVyafS37DW1CcCs13+wXULbXT7zuYNLiOrO7HGnlkFzKV1FKPN6qAV
0iRBmpcs3PycVt2faAM6gjvhjfS1YQ20woxVqEHqkHTO0dwhbfAdpwynYHNoT5GOTeuxX4oXuxDf
1ja7kgprYrVeCaUP5XLtC2TQHrg2bgetVd+nCNymwHkWFNOYK1EFethH+2w7sCLZjYmoieSKyroF
MvIabHUN6SMs4jCSEgAiCr06eFZn1b+y4FRB7hVLOFCCTcOZkKzY2oPQLNAFHBuN6Kj1GGFDR4hx
RhHhDt5QxWxuen9biMattUB1w9jl1co41bmfR90jtR385J2JKkZR2gy7PYGGb7OyNq0fQAjOYDrA
1bzCosSDqcPKoc3XiwjQuSUz0bi98S9/wN7RXIAINJWkh5oTTkbfvmHkz95jVYZAy0nU6ei6gXl7
yo3UdNuOONncw+/pnN5pb2zVNsEwEKQ/7T3B2pQUbNxCm0OKHRPTvEJVrQ413YgV35pC8virKpvk
2uaZq/rLiuurXJ2HlPlMqVxLqHbC+nLU7oJ90ri87G9gVi2UQjK2oae4wUJnmFad3MmjTp4X4YWW
Zvc0F61QeewPT8h13i+69zIYgRmnD8R36DhJxcVJGVou+yovrQNlI6vcEJ2D887xvb+GLY+h3SU9
1by8cQqvMfrt3pZbfFpQN4go21p8PJ9DFyMLNTiakpHAXbxXUQCsF35P1A0JzIIuFouP0eCSXiYM
Vg4V0K/I1la/Pj6KYmyYKHJoNX76HcB17TzOzuUroutbeKipUH8E4DJm8ioJj0/8tSt/QW1kbAuH
peEXgZtUh+BO977ZzGV8LpU0tThfqSSGDhqTbIGGSnUVVMZG1U9/RKHaxtA0WN8zkmdGUSfdq1Hg
LwuPGnDl+/QML39bfkvlUHY4ri2CesnnydMx2Li3ZnmZ7k8GIPdLrP+HeWTiIDSou7VhnuLHLPdE
E6yfVh9TUeIKdaDgjzdPRtdpNEaBP7PAeQkpTe1fCMQ+U1awojIG8TqVS9nYLUd7y8nUWvlH7kBl
BaRvctpuQZ3JqbTSlXOXTzaNQfZ45XkHvBEEOD/2yKDu4802JxI9M8HUxPc35byPAfyQnfTmj5qS
OVoAfCUIq+2NfTmjA92LQriEZXbjok9TfwB9HYv9o3iiOhwsBZMtVPoLTFLrZyCWWYgqsHFGbYH1
pX0Bah5FUlogFdJQzQ9Fdrwz6Bq2N3rgPY2x7iVLTPuj/cqEH2X79EqzY6i4qqmQFe3449yUagMv
W64pGLwJQ5NDeA6fBNLMpVvlquLmIe2UfJCUF9CJ5WUu7FKegso9qVprMPChwgMWlEWOXInenIDf
ATUHR/Ru+aTkdMiuHkUP4yffWua4ebH2mO7r1Rkua+V0ErL/ibpyTlfQonRQyjlP3VjoCFpwS0b3
Mpr3ZKnF2apmDJWEwyy4eLrk35RAUSyAWjBcnnP3Aej7sAR/fdVinacf63XzVU0JLveDNUqEbZEl
4dxqPlIraT+1BLJrB9JVUqshvtjQ/BhJe5YXJtEOEwwmxrJWuF5+qNBDRea3ufwz4Rv7pxfGMOUR
tM+5J28XcFoSYv0hHjmBoUH7o2UagetGTNmsu8qXFPUl0c94UGCW/EGGTZFiHj72XzDokCFazYkZ
HfSHYNcjOYmrWpl07tdx1Zb06Pz8mKC5FcHOjFk5FdQ++ulADbNbdDg2U4qAiyLXmk4u4xJOqbY7
OZNkV6IOwfphnpeKUmw58DpOOgKiSk8GXAyP+JnhjYI//EJ0XJ7DTzmNmK5Vs8lI16rzI5LgGkZX
GZWTHXdoNO4ngouUuOrSsBWFtyMYxP/8PXLuLVMQcy+6uKr3O9jSuB0CXtM5R730O5hhS3VidShH
/bTAO5krBQkTOn+atGJHBK+WNQG0ujZZuttJF8M410vBMphZ6ipr6LmfJciB+UGkcfCGKysjOcZL
y7Z7o9KxTsCGj4t0Mdbol2i+tjgh4oxZ6F+aXy2Z+WoSaQYCKrzkdx90xYNX3C4f/fKnDK/TDYdN
nFcrRR8M1NOb6oPhojOKjJC+E3y2qqcBHe8yp9nz6AFMxOrpI4oKYU0AfUFXap5gJeRVrEdhEwYO
uZtyQJkxCkFIlKhu4heoNa/C1M3v2gYsctNs6XQVMs0F3mAh3j2DhMdPHJhxpTgH5TNy6qahK/OE
27a3bt5bVZFjts4ldCX86K8un/3FiL0VNiFna40NM9Gv0ZLaCjom+fy8Iwu2ZuN5Wpd+ISsDlY2Z
Qf7GHsFzlmnRzLHkPzZwKN+oGTAwGerBYD79f62Y6jjldI61q2Jdtlp7lsA3yYfv3L+1wgnrZigg
SBypJ1MiiECBZYmhHJMhD6xjqwvi04QH4h/vIQy7Mmrduab+H1mVyxLBVRSON6M1TzqTg4GOz3D/
8rnTj80FjcOLFdoXBmx11LCX08n4zNK89227TTJoyuzYDD6/RD5fhLWqPaXEql5A1LTKIQBgcxrt
GRSzdVAlI4oubd/tSTJCMQNWladpS6Qu7sM74XmvCUYby/RKdEYwW32VEP4IaaN3kYUfABa/g7KZ
pCeibQ4tOdg5OA5WFIBLtUfz5E0VTh67UhUoFKO0ovc36lAEHe25NCrsdZAwfx3SRD0CIiHfbbNH
MP2+DBUX8SeZ51gQKzDnBD+xNkPJ4rp/hgnCY/ZZ0J9AOndZXhdLTdrKWndoeAuO6wWKJx/RpuEz
0ZnVkgNYJl74tcCAznDRq2Y8buXe8WtSJctHWS32fmDwFKY9AyAgaVklz9ZF1oLmBerAgIobXnXJ
qRB0CDGW2XXRbOuV5H7x4eEc659aD5uw+dtoKTOjjecXrjqDfb2DNFZxzn47JDgFuLm9c2rDvYgm
N1J5umppStQvWXvUMbNmc6l6d98Cgx20CC+H46yLtzj5AcqMrnbcNJFdSJZWDGtTJY9KVikcr5Ms
7DDO/+pDAAAW2h6swx17xXnN7lMxPL1dswX64u1m60GvJVr7GO3Izkq5qO9l+Mz9slj5y9mGaCsw
Ys3XNcsOpArERSSfdnO60Wj4tonS4Fkn298FqTCDqgR6KcxoyGcXEKIVBzIOrzKxfLWKEysU5jdQ
Kf/9x0EZfgivcQmPrs8sVPu8zRdgHKHzROzXBAZ8WQ0DcM7m3tWXVOiuRxZTYgcvoiza+UzgDwUF
rcVFwQTcvw4lsGz3fRcLKZx3PWOrABI3gMkD/5/thTMJP/nrOJ6BMfTg3kUpleIMkcDHU7dzlqp2
jhQSwYMTeJpT3gErCi6GaJuA4U+ODNCEqbDuNifBciEkAlhwV5PwRCVjggn6g0BeKzx1oAmvb/Vi
rDX5a4jkyKl0ZxCR/kw6onATEdt3Cp3GRCYIqC91qXV1WRF6YmZeymy5wKF0JsTsFvA0Yki6rOQL
JUp1Q3wUHUYW0M9UCjjAxxvyzcYCU4+wjTL1XsKHFCZIGziasnnJiUUTvdzV2koAjW9mNEfrh8C8
TfePB+aB+pZRUc+hZAlJRJ+1imEsPEc/Yl1AoFUfDuUFRYB+gIE1A+OWREhsKJGH1DYgpP7YV1Rt
kwan6OzbV90Egr7lMu42L6nnkK5qFjbKEwVW6RKz/ZkN73S0VabJA5nby9C7O4cExb+wEYieJjqq
a0ojvcy4w0KYC7LX/2Nxpp2DW5yfoeL/9LPxuHn3oeN8Yp9If+kk38GgnhNs08DiIBIhvr77EPVl
B7ZRxxqKzvREX9tdtTLCFMsJuXz2nNV8uKEq1rW8Sf/xZwsZk+wtFT+aRJksgEr15dbr2t16sDtZ
mh9ZSHwCFa9Sosqc/TCRd8HEzTSHb2O34TeYvx3gqW+0QgZLzzoOpT3n2/F01CwiLi3aDkmeXbg0
DvY0wrXEVYmzlgPJb53fJ62GXqJAmA8rnZRYt/ox5z/XOKeLznrjuNwd1JOv/8EEma34m/jfrQVq
x8VOwYynXQ3Hv2oW2C6f5qbAn86J6+sKAbc8o+CpxrG8uRQwI4v4H426l4G3YOxj4MMJ9JetXHNp
wSQes2cZjUgcVmcnTdrspYibyW4avXH0TQy9AvcwUEpx9Ok3NPAgSiMK8UDCOhv8S9mZTEpfpTiN
duqqbrg+gh2zODiE6VcqcyeYOHByk/LL8Ng+CP1swO5UdNoGFdcBPtTXedLGf52vp0dyfsMoUMNz
PoPbuCFKvFpFrf1G4imNflKsfmLMzraa0HMC4OTco1SfsT614LyZ/TjGi+wqO8oROU9eFTulnpLM
5nhOmFTK1vPihSdxxRQeRanv6TQirpXKwSkhVytXUqxboc9MuZAyji7IO00ffR8eQFze8ubl94Dg
99eZ23JzES2UUH1VHg26J+UhNSX76GWN2heig9WjfkBPPL/hHqp+T2fGf2xs3wXPFfRaXvMFt7QD
tV7YL1S3MREtAtYovNP0VS15doJIDfkllhoOBsRoWO1znmvE1mJuQCltjTlE9UCA9OI6s/UceD8d
U7iSwtlqhNfG2LZou4az9b4FqMC6g7uhMiDQOHfc3FSh6dtE2VORq6jlWFDxfdv+i1kCystuy+BN
sCo3UAscfRSi8fgVrW77Hksvl2gtuIHntKHEFprTXpmJPLRu5rpm/fXgsYd7hJk2JdOl5nH/fKQw
p+si4U2/2H4ftUpY1sud+F6T1Pzk8KYtCpWTZ1JJqHFntJRFQhRbKxKn/0VyPiGQUS55lA6wA7IK
GBIs50DbPorn+tbLKo3JxwWPA9F63IOY/yEo5SmxGpanIrFQdiOeyutzicmHoZ9Ey/+7AAE8y9HP
GEldIlfqRjOaM3Tj0OdC7H8GmZCwL5OHsLQWQY7h302p0WEonkvLJLlc4MxBnL80a0fN9tSg/IdU
ID4GEVzuJKOWSUyMRe1MHAvNaq1XrIZQtrKjg2mj4P4vaxGlpCBQI92aTF+hWSVOkO9OGgswkfgB
a86LkgV8VjhJ4tteR+9yOKOSOBYXs8MvGyn8nz+EPlS+FGahQuXSmspLvCpwfLeu407iz1BFXViw
dUiDtMGALsnWV6qEGENuJYu92huQKnZSesnrdO+OWDxZUV638QjxGg6vS61BIo/28hVZWBBfynEW
6F5GTvGRmtWYkQxHWnPNYWQoX9m+gov009XyvkubmvZefYtzo8eVHcq3sxP8SC2Rqvu/u0ngllex
0o2oYucH9EV/NRnLJgkFezc7UWv0k+SKVw2yjvu6bkffJpXmc/3SqYg91WTKq+rhfVHw2ao4acpC
o340n1TZXexuk1h4BO0qHTVxjKGjgBmyET+iYCuPt4FH4ZvUVXjwxPCZD1uYMizRvQ6w/1fm0flY
RgpXN0DhLKrv7PFz9nBJb6JF0LPNSZOAerjXqo1AUNFGUW4lQeg1uFd6Frm3KywLSQFnzFbK0DGZ
M3kQshWiW6IH+xuGkvzaC4FKASDEGRu6oqUEQCAOuKy7hToAqoOPyGFC5M9jYDdy1fdre+9SNu4+
iKqMV8nxVJjng8KB7fYQ7Uecot/FqSP2vaYiw2BGb72EBGFZ9Ee8z9swmB62e38loffjsX6H4Ejr
7j0aCxAU5DyNASbRCgMd06WvETLezGQAMITRP00vs90elnCwOuY8SjtyaGpB3yf2xsu+l/MTqjkq
TnHYUHpmnTGzaEKSXEFZh7PI/BNPdfNNbwhoBCD/3yQddNHhLOxBd3t0O7Ixt6jdiJ2KCkhZtDff
B5BFH1if8fcmNxhP/eGtpwvank5eAaKXnAPPZEr1JZpIzPcmp6v8O4eCxVXWsGYn3m6tjwPJcIW8
yb665QPJj9OrXf2Ue0gKBJYgEMTCQI8NjXDbW4L3PTXxI8djFZyjneK3z8Z7V/S72pJ5W7TDU3GM
Z4BO2goy4br4enzyKB1YM+sHnjvXFlpN+n2AhX54ALpZhV7opsolS4rrIZU82bznpUVJ+wX5cmII
W9cUOlqlT4d8znmrIsI9y7FpIGYwSZYqxF7695IvmqwNUyT7Opfdruv83dkIWz5J5/ScFDdn80sY
GzScAbcPJpvfC4OpD/EglTXok3P7Dz43kDYpZia3GMY9irSfZwc5Hl5NCwoXMk85n+stO97WF6YM
w3S4ctYoyd87r8jOc1Qt6vtZtuMMMuBXMZhuoPD1pTpuChI/T8vQs4q8/tAzaZi+duMVJqqdE02E
eo2RHaJBRP2hbr2gJyIpuDFS2kqeF+kWpnWUVcWmL8fnd1hwLG0NdVgkQlB08UYM3IHHgpji2A/p
npNEYepll1hZU16HiLragRP/+ymCUZ0NsmLo9NI+PRmN/9pfP//scXWPujNcXlk3WC/ce6uemvgT
puulCmpYPSTB6yFtDwfGpTP0m6TbsJvCbv96r+0wa6pIuRplu1Sn3LUGxgygWwSK6u+ZebzFz5xo
tQM7Lbh3idOkEthSh8pCu//U7Mrus56KWPaV5fOZkOVbiW4hY9sEZt+MveHGI0Kqr6yW40x+qR6o
hdeqdd3b0faWaA13IJ/cKBx7paiuxLYANg/71QJ1SJQpRujKyJvHBolbRJSmJbHN2Hu7b9A0A/70
mZL/qOjS378J9NuOe1FRy+p6Sy6uv3WhOr5ocDA6sPzYogt4QfCf51jzUvZ/MIzCy8N2pEUk79XK
zEMcBkVlw1HPs/mD9HPFz90ME3eP/rLUon7utFWU5kKaq9bJcjzYAWdDpWkfuilO8DQ8GPtP15zk
hbj+k6+rvbbWflIdJl3Kze2q+TOsH59HXCW6hTXcEnsOotyWFbTqOiUn9MAT9H0YZ+ygXapJDmLf
OOktsnC4jEMTRcnzqaJ9jhfwS1BZ1THr7D1tgLIr6x6dGOqtqehDHjaAm5IOVUoWh6bq31SJpdzM
YFVb41Fac4v5GA0wMRRgYDLarNLLH4qOv5myRJjQgxWAXLDfVrdFuFx1un9SvyrTP9FpgqC7Lpa6
O2NusOKf5VXVbGa1NxbmxM/jrnrXwhxVDk9DyKTLhYeG/GOt+4iMUgGawPcCg6qaHRae6+7ohZVy
i9TVR9npT5n8nEvYSFAIe9afiqxEd5yiK09gOqAka5Em+s4/80dCdOc/YWhVEekzRuQorjfyYmlM
gzG3kJgIMBJ3tKxHCpL3QY3tYO733C15V6BLckVvZy4DVwXSsyJDgR9uMLuxit4k5glC9YojpydJ
G/DRk/4zmi/LL//SVPsSd6+XZf9yRrgMOghKjB6nLeK9KjgT9FmCpqoEsRpxSE2dlVySH0CUkxiJ
YJB0xncdhyLchnRIYA4hNh+jjSSj3FJ7w8RXPYUWFE9Tzm1BWNOfR3878Mp/BeBLhWQu9CG9pAC7
NFTH1YBvJzunBifx5inyqUjy7Gjm9uw+cHIcZYlPA2M7fHUfzO3XzFYQYdjC2CctdrRqOYFVVmTO
4CwbXgySmrG+qQeX6ZrXtDWnZwsoV/8O13nt0idK1Lz1C0O4XcD017OJ/8vgwy5rMiRewojlM2cj
HketMNSMIzX8InPbW9h7l2iHtABLIXrixOlPdhwnBRBzbT6sA4EqdSdcFFkYqN9C5ry7dZzlQVP3
zry6NAHnc0xVw9eto/3OypEvkwbBaDN+Lu5Awu1tra5VUPQpM1tSAzWLv5Rlgr1AuzYLSflBbS0v
5XoH8jtrKk7MAr82qbnCZLqeNF2UCjXNzikFDaKRd1NJoNJVXGl6f01qG0gV1WPffXwAPbsHPuTH
dFVc1yL/KPD5YrdQQxDXv2p4WZTCxRcXCGlTEIwBGRsjUi+WMM+Q/ZIe9qSwAghKVzhG6OGfSKzt
zoxMu8Esd9PPi1n99wwrrJSQfIxP35GOMN/vsCzDe4rPE7xCte1pHpTVh/Z/qGKtt7AJ0yecNJ9G
8XC3HR/sRhcqhKbSzpUbMu0ywKK9oOo+Sr5cWWYSXXnklLHw+IG0+nGAzePdoZNSmdbT9ZtZ3poZ
bZlSNW0AL3bikzuKaIpdz9JQaTqyebx2QZkMnLX/UEKD0ED9ngMVCyhYRB8xPkyN8+kCjywFVfdQ
BloNnleDLOZ1RmEJtrKzGPKQky7aXpDSJPsIFpp14QhsjSbjdJ/BODgoGZi9ENKykN8sK1QYuatI
lpJIerYoY/2+ir+NdTzKFRhEjMLfViFSCPe580Vm4aN+abRi6aj0HlmjCxKLoNXJwMRim22EhFTR
pG4XPNDiRzwP9adQK5NgXD0xCvIvj8iSCWenK7PfO8X8FLijRSwtd3EmVsIHB+2pHkc8CbKrraAl
0l4cnIMJaGP84224VlG/txIaSLylzwf0Xoda2U6KT/8DgxUFQPeWzU15LjJKtzrYwYpv81bxYy0k
PHEim7ndqYyHimum1Kpx3bJ/r3nyJ80F5izzuZa3AUs7UN0XWF/yozaY27r6zsxpjX1mZ21xuqsF
1od6F8A7nlhJVye5WjzjzemKomrK908yZ1Sulz5lnBDAGBn19GwyghVvoEKTYzRZ6+yI4EOGxCjy
ldErKI55l88IttwQXi70AUxcD1tND7gfVCAHj5noX0HDN3XQ3HWPkoSEk9LM4JZRJv705j4nqo4X
jiBNQTKJJLO6sdxb8KEuxripPlB5wTEaEjycqxAopeuXoFjRk6nsK/+HJ+50ZQ42RQ8TkQteR7n3
LGPnNxe36D/z+vkxDVcxA13a4CRDKs8FmmreuClHOLNVYZq7bGLQdduKV1gT+jMR3Cn7Omili5h5
dnutuixNpZ91u4I46/hUFBbSIaMuBUxJsInj2KKmHeMT5BmskOMZXUrnILD+HTDKaZJRHFUeiyvw
7FXg876Tu3SDTD25AkppnO+c0LwcNByuk72EJ7X9w7HXPpPWGvDjZqj7SexcXh8FSpDZb4FAj1J6
AYDMbnT/q3NbErnI455WPkRjZy7Pc31mw+AvrhxnDlRyXk+YasvwnDbkL3tvXV4pm3ZjqvKVpxJM
AhTkXF8CizkRtLVCcjTOkuKlVqwtsMJo4dL//atIwJtQT7Ve+iVEIVR2m6wXM5fWAy+56kgDxtZe
WQZ5soxXAa7MMXQGnxjr4oTh4f6ccIOA/aj36L10Md8NlLx6CLQkT6DPGkECz64pYm6P/9icdCv7
OxVFghuKmCoovoKHjh+LUEHmApJtZPZlN7ftNbe0980sbs/NxnvlKcpW6NzvIMgjo9rRYsMW90NG
NGvsUhsvzcvEiac+BvB/vZFdeDg5+8qT6A5nIKeGU+UqGfgw975LoI6FEXXM5fx9Rby2n1e8skhj
QPx51a3iWdPyTUqmE43+KV1lvXkclaHEqb3FX8W2JaXDsj3iNjCMX1NQiThVLMt9lgS0INedammP
Ad91dfQWqMkwEKtjvOqaxjYJt48lG5qg81SpzfknnfxA88n7FivakrV/nbpihzLb1TnWMalTbzUO
zUhoZxtM00SRvNfsPite5063kIiRQFuIkVyb1rmyzyBe+s28gIoLI3kiY2O5zeMlPhg/BgdKE8Cs
i5W2jfBXEufRdCLFasJiC64ehkqE2ymVWwEC6mEjFraAgbLewFFhE7pAjQrIKYVwzTY8jNcYacBp
s2D6xjFx9TSiSK4W43qQfJC7XC0M0ZeQ640bOMlRHGV1WckKEOVHykPP9BiJYy4EOfBFq8UVIeJ7
CzxfLP4fHyB4vkI44ntS9+nLych0keA6ov5vCM2ipBtcuAopzpGnX0TK0dvN1Lw1Z7yvJjtW2jUF
59VT3VkfZW4vDeow28RUXN99UIK8nSv8D7VscoIf6cXnYEB8kNX3oX3ZOo4oN3uKOJzYHgSXuBrw
mub5xVWNWxLqthjzT/AxVaSKa3phXLnbJxDTn1yWnbir/JSugJbpOtkIjFpgkrvh7/hep1iVTwzV
2HuhyuybtT1VyC4/eL88ypsufvcees0O80uUPBkFmY0KexVvTfmb8Nzfrn50FpYizOld+lGXqIji
0cSRFE5pL2ROwHE3QuMJ3GQD2SYkGF4SC3VTjOHdC+wPqsBf0bSw32LiKTY2uhCNqID43vmOk++t
XjhgAAFLvVd5uIAAMtCKMOwGo20g8LyJVU1Pa724EhkEWPqaBoIUNa83Ulsrb4IHbMjbGpTg3sax
IbW5Pvnsg8DOGJezrDDxJnlW+0EzwJ/Jxv1BesnhVjrmYDo1DaHDQIUwO5/cXxC6e5JjTPX7S1zz
7GgLHfUoxlMHr5IP2FhWM5QFhV0kbZt1iz7U6SNHfYi2gGRMmHV2h3p0jTD52zO/Y7E+/0pIJR5D
ydATDHG8br7iasiHPOOPTvgjfR4OaflS6p17ap/Y9RJtLqCPXYzHx0mPjWZKH2QMgfqn24e5a9KI
jUi+LJG8yThxZ8WnbIF7ICl77wHoHzSqCvCC/fuFxKtfRidevDcz+/MSeC24nE2yRcoDVCm7LSlR
tpmhZbQlOOLU45SB+BRR18/BpqyF4MQrHHjqMC0bfCeTVQnQlJkwXx1NKmYEF9viCc3eWitWtN6T
+G/M2Jme/lJnjqZJLq38DWOZuav9CEWCF1Y/MGAHhwovCZbsqh69z0sOQ8iYeDBHwrFauTOaAeld
zan/u0o/6+wzvohe0IM07G6lOgrtiHAZOlRkaI27b6MPrZg5FHwEaIn1FZR1lWP/SvJ7GP7AtTdP
14kEE/rO0mKUcbjtChpultBhO0Lz1zNUqhnb1ed2vnTre/dZw/iPiYLhFZNXU7LaftC/e6qpndut
Q1jkDfCLe7ZtuYuewZQ8JSLxZFldF/Fklolt+Cv5H7857D9pw9VYQ/2dS5mcNbpnoQKpyiUTfN2B
6vHxfQ6iT+Q3eaFv+lspBC2p/rHLsKJfPri22C04Cdp8zZ+Z9acOhNqu6s9kud+7R4TRXEPF8cDe
opb8j6DjNhYvEDnqyy6t5x6IAGlsKgDsKA1ZoWgcOyIvDx2SrlVEssLo+eWwj/KKs2dUvebWkKwZ
Q9bBxo2d8E39Xc+eymuvvXlGt0XZetAOBibpiwE2zPZsUCAy6m8fzckdwr2Mvnd9bCXDZe5Pv1x7
zTQk01rhAORGznvXxKeut47rZdoll3foPcdUo0FgtmupjBTnhPGBEdVNg6VxDFkNXSClX/tQHAlA
EBapyU0uEh9/tN/Dua4dHh34VXirNckbOkP2u8v0S6cE8S9fdv07bXNYrk7Y/1/unBnJANCmXEaY
uceeC6NzAA5AyZjMxxcFueowPSI1rSxDKR+muqqINzi96DrI5oDkEuFlLZMSi6pZuAP/kZOxWRtJ
GHVnXedM9pQ9sBmRukuFJZwGaK4WzvgrqF30ylanyfVbWXpTQnXcyKpeAcYjLxF8GZ+dxd0au2YB
Mc7RscFuUsESqlDMnawjn29P0IuBR7KW5AW2h2T08g4BNnNDUltl6EsBMuE+rZPIO3VrxEtAApQk
SRXug65Psne7Q7QULpVq5Ly4GKCJhxFWI5/nC5u5VEHq5yZLULULoX1axSWHg1kNQEMSJuZ2oaKA
4P8RDYtNxrkT9I2+oj4lEPIjz1ORZyC8Gzj/AFl1FCdTWN8+275sId8vzE1WFW9gznLVGhQldFWL
rZKmR61bKAKN4L74Gtu61nlG60IYzMxkqdyVaPaeVf4wX0TElrFYcPiRvG40BdATdT3mVJR3ICHQ
byNxAQUrpahHKgfiFZrXilpJFGHGP9uqsAarT1atnoGvq/oqoJwM+S97KUEVwixgmwOM19BVJZKw
/lkWKNzw6moRkbqfMnsLEkqKL+fvds5zBVgQlG+Cmt2F01WrF/C9xP0oU7meE1RTwQOEsXgcrsBD
x+DWc0IM8tpqoKgrjRBWoUynsJooRXwNUAxaSJHDhBLYFGxLTwxAtE9cCxZssRHHVQZVOd6eMXF+
KpIN8pCSlTmwJ4pFVKbRj13LYE197pUpEqfzrGTyRKA3NbCqCnmx/PNFfufc/oujBk1QTslPNi6b
KGtDZRgQ22CKoVbatF31CapLyIuUmKAXpbWEoFbHW6OsS025761kK6oLzEpMgynVLTQ/p9NcSLy5
V/+GuPMkxJmXYvQ5c/sO8LhJ2Kkmx1AbokMEGRVkMzux4wPEYM3Im03YwavLPRfmZi55tXDmP70r
KrwhLYussaKZiA25GsyfNwz6Tj53vxjUA9OeDxgZH48RM8KhtcfASjMAlm9Qu+jMurnTFUV8Ge2F
2YxyQDhq+vv1gDuW5NttnBEBF1tyH+JGhQpnK4l6sC1ZYk6eHQ+8rw/HDPi4ucP7s0zJO7c87J1q
OkfgNNl8YcZhJ1ouXKChhn18i7JI4dXYh47SvPeAyiiyvjGJP5jppwzTN+ROZXpIS4/xNJNnqiFg
EvcR3KvCZxoQGmAvUHCWhnmvAiNOgV8NsQZzqqi9KTs44NAAopsTI6wrkKnmtx6kIsWmDshh63mz
fomteisHCpOMdHOJwrmavx129iB7rVFT92hIbZsA5a1FiR7YyIuQM2sVJ2tLuUhXFT9BeKo74jw2
kpq6N/XOeDa1wcr/+sRQe8JpYDWUIih0ROI2MJM0UNdjv6+gNQaioRTdTERTzaaj8SN8wx1tSK8Z
TPmbP0KzIXWaiF/IZKK2961enmS3tUnBFchoWrYoxjmgDqpctfZcC/Y4b+30w9r5xe7auEqER10v
Qxdip33WYFm2f7VT6xTX5E62jA08hUmv/ggsLseGPla5RQf8R0q2eUS9l9px5o0dIEIPUCqkJHPQ
EIIJr/N2qtkXm/6bKpbkTTibIbMx2USqeT+iSTVLk5EF3yr3ROmXdY9fRJeGUAKvjtylUGnmIUbg
yGJW9jEK96eu5o9odtbMjs0Mr11ZFMMvH7NuuTnZ613tkzhfcWcxpRIaCnGNvl2V6I5VEsG3O3nG
W5EcYqju2ft26SqCQF5B6uPOzU0235YpGralqRxJqRjdRj7S/28Ozm2aQPIfVU7YpA1xNn62vcvQ
IlyCxWyxYFPm+qi1o33WcC7LqJSqzGXC9xieSKQwC88BpITILHMwYtoZKLPxxP3CCDWA+8z3xsYw
zm58tB9tR7O/xSLBz1vdET0rtx7H3Vge+Ea9u9edzsIYQBwxyHXj+HCjKOxL3pLUbON8JIJOZ7Nr
a4Xl7fF6hKNblXTBMXSwmCiDZJHK+KCbZlkQw3EBhjfbyzn1vI5Eyweo4RsqRcIv8zXhfvg+OcIi
2l7BRSlfyEpmkufkFKYfVEyozpX0BC7rwlzunv76M/gHaysk0A3KxG0QwrIusHoOeWKwVqkH0CA0
WErgPxu+ReJKj5B+Llh5H51oVuU68P9YVevT2HkWeMc4qCKb9wUJirDsUucqibNQvZKg68kfJq09
AFSvrpEUl+2n9a7P65QJx2rZ9IprnTOR/6tKC9HXiEHtCFGfJ9teKf5vYi7SG6L2w4j2m5Vv1YsW
uvBBkZehUGYk1VgHjgDTv/PQtwFhJVy7cIJztcVQfxH6sti/eGKnmNFqQsYdf1wpS45T6bJI6/jq
57fn92G6t8K7jSpA3d8ulYXW14HB9vaw+FRC3WUemCd+gHsCU3jOV0Ef+8uJJETh2pZnt3h3ZR5T
Z5iP8oI42mz/HL9MdBBgPiyEvOhUPUr3+hNU0MyXRLd80DwBdMlf3buhopF+5sNwfQcBjAvqddh3
sIk3Kd503kuDaC6/KHsEehv5gF8V2sX1bRGzpNGTUHOxUrrmf4SafFj6yDknLlbAq9XBWBxqFZiX
F05xmwqWJzU8q3GxIocq//341FW9TxRIgnUWolv4L1G0c24OmGqlJ/oTw/wWYMvJjmpV2hRlSso9
XMZMVz8/6nwaOIhT3mOXqwJ+sQ4hA+VWRfiKhspSVFRB0+d5oFacNoJxVxc2wt8RzAr2Du3QPku5
/0aa1v1wtv2XXI/XYDCv4G8ogurJEuXigKHAS9pwQlxbQYA2oekeEIR2SoZMiVS7Kpso1D5FNZeL
8FQg0PosY1md8MrCnN/DJXyV/RdNWmHNz1tKoSnLtpGEQl4ZhVWZmfohhvHAlnFBoR+W88VA2ri3
tmdtIKqS9Mg3hDFp8vc5XKu/f1Pi/khdK6iVTnBMJ+IYfMcEtNw4YW/G02X9Zsf4D641vMdNObis
Xv1i+z6ODL5Zll2kyCoTRTs3D+Lwaxeb4PZYP5CO11AOWUU+fxQmu/TjkaT7JWferoVObJa4FutR
02fxoQcnE7tCIGU6S8hB0kDLZPAq4L2+Rh/MZR19EJU2JEJdYm/aM5LGPr3vDBc/hk54atEKrRKt
0MjuV6UulyjgtvsWDY0QzrXgtzZzmr9G5AOLbKAB7yycMTRn5QqBzD66Or1hy9hRTJS7weNSC6Mb
eQKq9E00t/QMhXXidTdHqf5eHXCRysRtzVfaUFiMMexKRXT3x18myDKKUequGGrnGMVjNTV7+2Dm
WuUMIWlZnKzQSEccC2UDepJ5Qyj1V51t20YdCRoSoSzD0hxjiUmx8HRz+DBD5KP1jS/02vQxEk22
sSDTFmZg535q6GLIRfXmPdLLi3mztSb1d5zSRJxHL3RJTudTxWsqRI45MUQzc8GioK/hvd971KqG
xIw3x7aS5ZWIOfEfb33JJd3zvNg2oRLFsrnEUQPqXXGpuxwoYlnHQtgbJcjcjBG6wLjw7PBxWxZ+
+TPriVFstqQFtkdE7YQjdGlyYIS00818iLzVc24vF5ZP/0vkr5Z6TYFfsEU5aUc2bYPORoAUav7X
ix+VJBpjqe7REJ4HfLcd8a8bYuZtRNAykt+gcs1vzqPrAleYnqsvpHF1MAXp7MOoYj0xihopHR9R
9aRO7VE3gMk8F12VHE1qs5sFK4czULTUbopL2Y6dhNweH/a8adbvfFnL6O1ChFQVXECq9oDQgyvf
vvx807zJ5ic6RVNf6ABtYPfUC6hvch5/TlPNfu+N77zDqVuGhrNKb6THx/BdCmDYDvzqL/VP4vq9
DSKb3Cxp9J7U8ILeAEoksA19D9FqDewcwx7Lk2dxTj6sAN9SK9UnjJ4c0nVZ+wyGfD6jF9j/M1sO
QVe+J8SrkV9jpcrhBrgLjPZuXQTCdzkASHCEhm7++LPTGwSAaiWYgYcKcTeAWkN3yAGbEHaJQpCP
IjZ8ioZOBgawoDKtJGb498LuPVaEwhS73nLc18RwxquFtK5OnAPNNqbEZocVFZViVfOJtg+WLzLp
JI7K8JAhSoEJyF0sApNNm79yGGv+sNpPNMhTih16eOGmonbdZ4Ad/yCB7GeDeGXSlEvwg3kLaw5z
oy2mVnGaqzMCiBp+Yg26pPOppy+ydvZ4Nrf9gRqpdDgr49jdsoPd3NMpUzeA7ONP2T0XyJJxkA12
/1v6zCYh8CSrZF4iTFU67X09Een7FazijG7captG3GzvN3ODh2tGk6lCUB8tDSXVrFz4EVR9nsJl
XSISNwf8fn9Zk0ykb01yWkdD9Xm4d3fHYGP+OX23Yb+KawVkDtALqoTjM7fyc84vDC/77UXMY59j
txqxNcBAxcH9V+xGjPZ9Ae3n2kSI8UUwuDlA6gmiK7xectOzofdag8DOlUqXvWvg/hVTOtxuUYzW
JQLbi88qDRav+q9vTkUkGrekBp9FYfWQnmcpgtwfIjZ2e2aLRphDyULtftswPPbbsCFzovQ10a+9
HB3MzEhbz+w1Bh8SYMuTGhlfcMhENpImgfjrt+9nYzt+R9+jQCL+161/2t+sovjLW9HQI5fKtq+H
kfC7ugmBIVAXZbHhERTMGLO0fOL8SRJJDuEgAjPXDNZIKdXzw7WArm8+aX4hHXj7f9QOXNfH+ELs
u9MC1c8uNd8opXXINP6io9eoUbMbPWm2qHNVNr5lvb5AUs2+CbpZYCWwgRpZUjOpl3b5s0rKxtvn
YOhkBBfDOiG9Mc2EiSbFYWp4yD49ss5nu070Mp6WUDHQa2P8zHRFTZphqv9FByHU8Nws/yfNDRzx
AfwwPyrlrGhcWdUFA+FHr3bdpS4Jnhw9GxIKGAEaQj3X5dEtmoBc3GVXygs7N7Lz1BucWC//Pzw3
5OntPEI2Er7Ly53c/XX9NAzQit1GRrGRIXTVkgGPkGFF4u2Tbakt/K1aIbDxPFwFFBY8z06eQCTd
wzkPB7NycnGeDyuANZRYErdfc+9RZVMGTkYhay0B2yV4EofFRsl9IOKz9fbv6VnSrke6wkFWDRks
wI3fbhpO6C5ZznpWYQNdUioE1Mkh1t+U/4Z1rbZeD+qn/SO/OGD+AGll7DeNFLBiVvjZDVHT3nQm
epXd4k+BlDNjU3vvOMT4Bblc8IalyQAbubco7zMb02WvYo9JdDbUQJhjUh90xJ8vQZvRyE8IT5B4
uYh47Gt80DxPi31ILkPzpFvvQRpeAeo3yrQz/lQCbfH5lY+3VIAAzaH5ODf7GG0Pa1OKkQIc+chy
SL5qy55JiKBVzOJ9xvIZe416xOyw9FmXw+PbbWmOwSyvNqwENXP/ELLTH9RJ2IuY2qSc0l9MxLnc
UQlfbi+jySLwX4uN1yUADnC2RwIxDjsYfFk3ZYYHpTRXSatZQProF+jAXE0j9JBPHqz8hWY7KzyZ
I76GlIOoRx2emnpcuzYjqtJhNmf1B5RWSTkjmniqPtakAeKhVrc+9oIuB5Uf7r7MVB749Ysi9NWC
9czFI6TSFOf+aG86aw/BATl0IL4uPAOn4nCW8quojmB0weuyST00yKxvtJwP84NPjS2mxNcI3Mru
lBR7W59rkEqYv/NSP3WdHATOYA8OWOjUU7xG4O1yKqzYzSOtJclRShfneFGdU4wO0BYCNfqy2JyI
VOQxXpnMouIu0lSD2MkVewK7gsYxz0d2icr4GPjgp2p+w7cuGOfcl7jstdLlTCp0UhQP2G5h/CXN
1bi2vunaYMpQH/YI8nNJ8CXkF2xbiSlu5imbVZJln/97sOFlvsCxZ6HXw0s72Z0NTCilVSQ4xWgx
VtxfnqfCaTJRaydEhDeTwGt1Ter9ifmZj4brjcTTvWdgRD7HrJmby7tyUPpQTgCVH2+JNoIQZSfT
OpzVHDwIAfGMqQvdXM3iGBIGh2vhDd3gmVLla8FJ8bhm+lY6yrtKBgBm0YfXaID6ePBko5SxVas9
Qi0W7LFQpGBiYE7739GhHlay5nyaG0jIRN3VsrmAaPQyowd31+P8L0imW5huBnHF6P8kCFuqZeVH
gs7VqG5be+llWsqcOGEvIjtKXxG2Ta2P+hdYaHiNKxQxZrARrL57ZebIQ04VZqSo8mGRb+jp5XuV
HHdJhjCtQYmQqjZzIFJgJ4fv0kEZTYvonFbdLBm0nOd6oX9+UQwXaAVOfHXzq4jZcogMtiaSkhuu
1YNXAXFRozEKWN+UIQUN6hl30LEr/yNXiN/hrLZFNEu8+ntNjj9LFZuE84zE/JjY0lPhbf0r29vb
mRzPjNlcbYFPPkAgb3UrKcJo32xY8FOU1105pwfYMSnkq2j+jXtqMDTvLJFNOzkD5dJvHF3QVgcH
faXQuYBfGriYqy6C6x4Z/niqODsYKcoWo6WP1F7SqwHZLvp/Fh7oSbwsm5ebo9k/RcxD5kkO/Y9i
3gW9cSSTHm8Wm7F9WNbpOO3m68B5nvMlJF9DRfLarYMhMe+DxGksh8Mg3M+wy/+WVMkvZuUCkyDw
cFyLzx30xPdJ8ZECjxkLDnxQ4PIO7ZRN+0PsYx0dtzMuO426qiePpuJuQDv6Oibqcq+AexqsEZxp
vQRCM/XxIIEeDOR50YLLxxH1sVjm/KS18UFF5j24Jhjw7Ec2SLVTIHo5XhdA7iEZ5T4yENgkMdG5
ZooaE6yOBE3piSAbPqb8TC1iK/v2r5u4UEIMbB1IRzTK9tnxGF4s3QJrOLtFI/1m3AeVlIe9KY72
Odf7hX512Jq/ScNTfmCqA3KINJkbxYPeSf5jZQJQkyH91KQVmhk/L7nHY8Al3Mshv8SpkhGbDDHg
P0T0SeNhhkTfyxgdqfjg0a346XVweroPQSgIeRTfgl3T2k/m87ZafTwt2XKE8u4JidJkA7gY+1jx
GN/pluNq5p+ZYtVveTC8Ysxdrbdd8E38Odm6zTF0NlTZO4vPlmqssuOP4zP/58xV7hr4SEA5tc8S
7MGZag5Y5qEm35JNbmrEzqzo1C0mtQXNcKgCB13d5bajGyPwes8XdncyQQPzOGZrWJVi2CeZhAsv
Yi0sl5SriRKeg+YQoOYBvf8CIQk61Gi960UDKOeasgHPRCy2lz2SY7cqIvu+iGfoC4zeWAGZhjan
LhcksMBSSbQHJWTgi3kv+J+wtLPRAblRy3b5YWR+ajJ310B8cLvGejHzfEAu8DxImuvVcR1RwcBP
0oGj81V0wpTmNaQWloHGyqZakEEyvnojjHIN/GWtFd1IvGCJCzuecJCoyHAsfsT5RM5vOSb9yDrq
8PoJOcBycZGXvyuJ5kAQD+thZoxqEppa3z2iTXeW02n9GPutkUKQ10k/eQJp0PASRxIFvWqtdLQz
qNHOuTWcAfZpIJ4/xiSgs3+DbktbCaiX/6SVkmFflaLOpcFR+w1nmMSzO8ALDMpbHthqIvaqj4Rk
59sZS1pCCwvdY7O/bhUDE64LTU1gQj9OxvVvBrQXcrlUm5oMEShDNyJb+f2YZDqk6G6qzZCX1DAH
nPgpL6Oo59ImkzLCWwup+cuKuViabHqykw3kogumRg2MSOB7t56VftqtPsGELyW0RhgImfxbXXuf
WLN03P+K/TuLVRFUb4MwNLgMIsZuXtkkBsyS+h+H5hSSbWQMaTA8WCn5ZWpXoUfKYO3BHPRN0mDT
EnFRop+elNehlFsNaL7mqaLJ4oQYGtddasE2XkwfsupeHgemUzcyu2aIf3aNtXKHoBCMC4NMKGUB
6QsSHutpVrPS1FdLsY9EmwZMZu2/nbhYmJMkx4Alsb/jcuC8RBroCygQfDAI05Q0q9S2D0MkYXIP
G16Tw46QvRtPWnWP8m2HQr3I17Mlnl3+NpbC1/eJuLVWOc5aOZ71KXX9sbiY6tiNGe06FnVMIK3A
/sJf3ShTvx7DI6YzbTp6Fwp4FURNniNLFarZfq0l6n+cp+mDZRaWY4/GsC89ntwas/y76Yy8PSte
cS1Si4UUF1d7nMTQ3xLrGdccZXICU8337MtVN9D7qge5UOVE2M3i4D6WYCB/z0U/QEILv9h588Gr
sZuDdmfOCzF7f7M2QtWD+MRBcoGQVLxWxNNBjohumWUpOVTgANt73N1wHJkukOo6SbhY6VW1XokK
hdm1p14UOCgEDQbsnt1c6A3o/uE+J/LglnkYj50txy5lMcxXnWNhXrzEfwEMQWIu0rDedWsQbKh1
IOrg4DDuJGXPloMNTDUmC4vZSuKvn40AaIvv0r8r0q64pkk1DNJZyIxskeEiYk5KhaZcZ01XVUP0
VlgohI6bc9KMJjkXwFEIw9BCZJ+/Pjg5+3qiPX/+SDuP6txw/WR7gmSFohGIurDKYHDHkqsfbEJ8
bwWPstvT5xPEFnVptjeWEV/AQgbaIY265WTvCBcSK2MacJmzNH7Jg5oTySV7mpOeseA0VSeL5XDN
i9xaC4QFevyvAn8XXS4Q+GCZh9ns8iByPjxPuM9zzvrbLytp6ubS4IRuxfI2l20b3Ssy457mwhff
iYXeIDIhR7Tofm1f/Mob38XVYb7kof2lq7oz/IlCHUo88LWygslP70j8kpxUsw5jdnMef4DwH59V
RTMVmJgyRF7sy4h7UW2OvvdrBpSwjBmfNRrOYnzBdT/GxppqmeF6CUAxMN40olH6Na3wMrOK7YCp
NFHil1gTpKhuqWrF9sQm7FeBwUD20mubwrMwimOovNLTX5hQjJtHwAuPgMrVDbc02l7r5zFAyHxR
MoRxBv42wC1MFgVZDD4Az02Q28RM858XJejB5m9xCidU3h3wRh6pULMMai2zWp4g6+7KH3PCwvLH
QpERe7rSmSO09xn4FkN6oD//y7okoHaPU8AeWUlcTFOeJFdh0g9Wc4IB0K7elndLGSlCb/4tf+1O
p1yo0W+ZtBV26D/8IMNgqIPmyJhqiB/kaMpa+mUBMs2XaUQutGwvindOTzi6LL4ThC1rRyUwMSBA
W9IWmDFsfAzTDLxkbTvtUv232dMyamAhvBRwZBLEF+JPMADGR/F4TxH314bxElSq2hfEcflU+Fie
xLZC5f4eLBVTmngx3W6ta7ij/8yozhK6821WmtCZ8Wgk6S9AdaIypoXR+l8U4DPh+v1AIINmvueo
i677Y6QCpzyJhF1IlwKkcMJX3fZfVYm6czwpYSwEdLgfNdwO7And2ERwFqHXWAKu0CJxgn64gLoI
N29IzjUP1R4g7hQ3pm/wznCzJUptsWt5tPm1ufccXo9rSJIEvfGW+sqEonx22Nscj/PtRMRJjur6
N3Fd0H+C9Ir9iVGouBo7UdCDQqwftNO21NZPQ+0gOinOhG1kF9R3SlAoxmwIdu6UR0rk6AqTJAQT
zZKm/S8pAeBuI37GsgTYU+mY7NpRYXpwkQ+ZoMqmCZRsqjeXNwyB2smgKN82CF2vF7mx5y8WeeqQ
LTul/Ze1v5miUDECgn2mMgcJEzpBoAqHOBgLN5I3AKsP0AhhJsGlvVWhmPNqlv1OO+bAICK0qlKJ
22gQUs28AIyvANyC3wMsGTCnj9QwFdKtwGtosF7eaTFsdS75/uytnZGfLVN2p8pTwjbkjlMrlp3w
OPNTblRly0ZoO2y2O1TuFkfCI3VVUrtuL//ymOqZOK8o+1pZ7HZa1LZb7isxxmmTyd22vzv53WRO
bpofq7yVzXvRqwIenI8KdxjkGGT5lG/qDx9hJfNBsbXcLUP8T/oBVUYeMYGbvmH8IB/DlweIbRX0
O3Tql/576NIVUJ+JHD+za8ryoBpaTAzdLC7D7l7+OvoZGSxX3Q/FwQFKNrDcfs9bDQq90VH3B4ms
5W6KC7+RzQsqixDX0Sjvhmxj/QDt5KbbOIkBrrdY3VUDIgAs0XpofGxDzd1bYmzC7os2uhblUsxZ
ODg2oCKB91rM18QTLPk/dn3rO43c64PzVIo/B1MoiR6T62RhidLtSJJvsAKX804lNeMTXEOoBs1k
7Q6TexGPhVNW2JSfCqCQvjxzw3MTzZM+6w+++cGFRQUWKJjROBvNnvyoCsUd8cJ70uwvxWOS9WC+
7ot0TdSnt9o3G3ZOINYtmnmCbYNXp+bEFubA7EogL67mKvdlWXDbmo+am3GPSQbMoz9D3GbgYwEK
Fq8lugwfMXz9QYyE0JpNNpv1/RLqlbOukSUwzHLtlV+sdkboDVmHpmbuPfAXxAQkue2KamxXcLiU
RvXPmPyQUCC2kXXStNQjRHTbY/IzDJiHOGkc9XvMeOm4EHHYNaBH8PX47T4kx5CX4RyvUgm7NoZE
Kp2fDsisEyZPO6kvsSuOV/qOr+gGGgQquyMNGMzVBeAogIkfP3MBzxdqw5gN0D+GKIcJ5Ilj1Gq6
CYl3Ix3eGBcCYWuRSKbF+5Aki6xO6vipfL5HsPby/xrS6k9PLsa0bhQAKkhtcPyNJafehDaKJ7l7
GdKyYizvbbSSv7OzCdmbn9NkLPBmti494/S4SiM3nwqSmljmWql/tHrmLkwo0eWW89a0twdRZbtt
BOZrqzhtnEMeOPxmy9FR4deWhpz0IG2+6m6Us2I4tcPkZgsuTWaaHhOfcp0EARrIF1kyiiUVzTJ0
Y8iDJaJqtyPjPzjCQ4HREjZUTFkI3D/6HQSK+d8vvikymOS+8XP2sFrLQfG+vjmje06fi7KE6Dxl
EGkKOoe3/VNTOLPbnGUNCP2BdRnGfX/kEb7CXY8Pm1cc3v6u37g8enMuqy3FBJkY6vpfnrJLQzQQ
KkFhJLWJ1AmpkBjJ/z7TaQnwTslnAJmUyhFkp7/u9ldajEoNwdqNDfbz/4DC4Wg55j+mP1yTuyZ5
YOuK1fJan5xZ8R2wUIOhTiJvioxPKDjSVkEsVfaroWzx6roRzHZBFrlEApG4BejvX73zCwdGQwLf
0Mh5i1CYC99QdRp5/+EiN2gEg9yehxJiR19z5PnQNeHkvJ8FymmBFrD7tkh2qo9LODmVELxvknk+
eRMSy9XkFi8Is/0+rSZzBV+wkGjJA5BACKugAqW6IojD/6FvOe8F+Oti00ahEDxg9t0N9/C7iSV6
UTousUOHdFzSAuUKduiRkNd17Ng092K9eEVM7rGaT6+NFgxI5mTxyzrYn+vjgK09497t2awUFNx5
Gwoc1l74jaSAIQtMf86ah71SqsZbAvqSZXn7aCBddvPBjNzNvd8ydOBzyTL3DpdLXYIF0ukUhJnP
hmjoqIFvSzsx4xrJwoisodO7yNrYNxk/eP0uJctRgEonVqF900ynKYxt1oMrz6FjVPK3JI6dHm+6
2MeaI+pUb6El6udZ+9S5cm14d/e2MVa3iHUNDBxE4bnYh7bA0bc5wMDz937aou1gUi9sjYbXoq8c
rpxWoqL9+2amN5jD7UJJhdyDYl/HhsB4yaHtIDBSN/afW/WqNmzUhy+DYe9gCLiXKVJ9Kmtyq9bV
/1qVz9roo1HQiLZlFdG3ZQJf0qovY+6ZCBUwMww+B5BUZiLsnX7F6aUa+AZBTBKjQvycHEDcHEYu
bVcvAlsAuzJ7gJ5tdyu4Kit+nj+3hwzmh4XXVkQ2OzLut/46uXdLmBq5k/dwc7RYtm+XXsFfiOO0
ywuZ4NX802WDfWIqBMcTsq5o8akh1WYvs1n797ji8AxXD3god/07l1tvq+RoCJ5sJZC/WQp55ucp
3BVAcOihQerztwSGdpzbquM/h3u8i9hZeXqfDpwVC+7WLebF5Kv3BCzh01dRPN0vVcKacVEq/G0n
jSXxuhIbJ9TtCouJSYhBsR8depI5+aWTR1qquSiztAxa/l1+ILbFGiZN5LeUtcIGfp57+xFlowPg
6v7qygsrjgSehOPV7C2nQDtoBWSUaYwsLRhnhvGQnz2zvQpSsMwcuCqenvQmRWTkuZU4Ulfl3CWn
vJ/QEYh/mLNlpV0bhXCfdin8hpIkm4uI3tbB+SOrb3VzHUdCzRy9vIhWktNeZV+T8OazqK5yVAkh
iiqghasZNtlT+gokcHA+tfAJJSopbbQaGTimL/uSoC4iNAHPFn8FmlT0Zy+rHc7x3DFWn4ji7s++
jr90PILBDjxaCuSLHo/LGgzJer9fVoUDogNrtx+A2lUu5/AASIhZn+yWB8/ZiAY4352F27MyjWli
KXiKvyuE19GRELbW5chQwFXK0oE9jvHMbiTsBXYDDq2CmHgF5uFPWxmey59ppeU9bG9pr5/ZwxH4
RwasNBhXThJ79xCBT7uIly2dnYeeksEEgUKA3OJnTVK27r9Jgy0C8/pnDVDBu7jMPKm6b+ezVENJ
dSUTZQ3ojX9SDzgQRiqNoSMCG1T3u/X8pCJVYJId/v5LWY5xP7aHmXFaFOBWyl6gzKGPMVNSVihU
oOYURbiO7mzUEhgfIapJv++En+O3ZpWSh5TRoalNb5pTSeTpMvM85QQXzyxULtTNubMF29qeM+mV
2gan2QCkaMg6t3LkbU7x+K6lK5q3hdjlL7tcLERcyPjCnL8GCk8QTwSX8VMR69aoTHeFlw1o/8Zk
7/xr8DHTtPSM8A2xPNAlLLjWX1G1oTTh3YeLnfpYElovmUopGNi3dajUTRhhAyV73l25vwSieybN
bHHFFvTXHofXXVtPMf3eA0dJIGPKv4GoxiU2Nvm9FkPUJ9Tr5w1shRtZDDgsnMRy1jZMYEpNq0oQ
mCbRwerZHf52andtEsg+t6bvVLrNJhbDNBsycBrKs2VhQHrs+p8m9X+ca7F9zAFeQYIJsZe5Osoy
mMcZvKxM6qNN+499WT5kVqcjhM9jRloWxaVBfKT6+vKsGqiJgMZJn5UzQZdYAj40RiL+tnoJM/4C
z4MeRS1Cj2jAnheG49qWuKNO0if+bLRSq2OC2yUUqRGs/9Df4AVudSpoNAcWHblbuQ+MkqCUTCtX
YoqANLNbHiFjZHj9MD2BwzSbAtSuQKHA6lFmTterIxK7OApthWGPhTmgZ1BzL+axgdz/J4hvL3s1
OqATqChrSZLIImqcG24bHkWf0lHcjRBku0AAQ43DuMk9vh1bNzGFXQXp3AFaHGE+/TgRNX/ccM8w
Rj9IrhS1AqYw7/I1Gz04NydYPV37p3zq39Uu6mPbGLON/03hLuNqbX/MjQs/YhtPUCisWP/IZGJx
NwfdLDg8BLM3gHuGaatQfVG079QNGfMQSjfghjrjsUr1Q9VpmKLM9Ec9TZSwDJTzy0+7+zpTWVgG
Om54Urs9zp+KYnG46vGkNeDXAOMo+aJoIi/nzxJPVl/NfveN8IDCVciufqTrnrvdPsqxmaisqXzD
uOsSmlenrpzfM1TZ1SjODEKxdtHMlW8AzjGf2PiZS2WP5mgA9mcUFkN0YceB+2aQC/u8+M1s6QGp
wv5AoOHeuUJ5wJRS0fZWgrRbwiqnwiP+4ftLeoFvhMEaZ5N2XysmH1aQELu3dS6BhhnsO9iO3/q9
ZQlEpDSOT3V0j9C6Sqrg99153zt5/rOB2cOGp+oBzbhSdsqaI4h8wx0uBhm0xWXQn1tP+n0I44jm
nzAd4YEgl1fO+vEvWBr4rMI7ryyE6pKxHh44hX0YTJJ3H6ql7trnVHgmrRKdV1Fc0UkMGme/6XIj
+TuI61vfaGO3eLEWtHs2nJv4PMAjS0qiBCXqXcawwOexrvaYPSTzE5CNDaYi3Pvt5cCXjKNYSB1X
tL8Up0SxfrAsC2Kzxx/WveE3klQE4EnCfzEBa21dKaBUsNvXwvHLVI15gKlqSvqJfPWXeUGqlIBv
e9jcnaBdLnPZOZE7af6SaoD/3mvZw62iC9L1ok28ZH/UWjzyq2NVaI0ik+qgS/kJ6sSQqCRbSb/D
LAeEme0DH4u4wMt5FwdJ8v26urrPUMVwPexWsWQcTTICznWYCBR+KfnMpmwMyIYtJSa250G/kvYH
C0fFdQzPOJPpDuZEfICkokOwws7ruIxHRW8zYqDCV30qZckr83PqDgFHWaBJgAR66oatWv498u99
6wThgnXp0XTAzzcuK+y/DV9x4U8AW3l/VNQ29QFxV7rZlMBrbgVDYRUKoO4kM3NhhmtMvOiHJPxh
8Vg1wXMKWpQoSTrIXuZIUmiEnUbxXDoumOP4gKkvxrqkhh9K3QmoV3f+EP4f6cU6Kn08s/nv7vKs
MygKwYoSbUv9z2yydmaJjnGiz+nnf0Fp6pxwd7fDSM4eaNVlZ/lT1Hz5sy9jWC7pr5hF+bgOh2gT
8iuCewSjSke70t0qjdgsXkjIxBmwSJA0hqYYM6SEjoIlBI0hnLACryEzWVYl6GVXa5BNQFmn0UH9
siuHmGvzFzk+MGwIDETauuXp7+v2ukXKJGMtORlkEeUR2sRRN5r0Hp/yW1mFpIuDUNk3wNA31XSQ
hDgZb5NwO8t69mTu9ATksqDkwFouIVuIAN/7M79WnXhzoKw1ijQHtw25V3nzqfStRVtW3SiZycZW
KPgLlh9yj/hTOA4tunx55FH2naaCHcHVhn92l4E+sGAgxytZXNsQwQyozMBDYF93tufnyenUWQoK
S6tp/wazJU7H6hM1mebdz3VS6+Upl+sqUNt5vT2oNcY/lnBTh1VJQxGx639H6Zb9gBaG6oA9HCTk
TETXAaVjZQ12CMYv+ujRYr3LGdCq7Mm9wg3D6eXj0dWLP1S540OvLNpPGMVj/Pg400S0u6t7fJo5
dy5eim9r54cr7+jSc/YyMR5oLjkCM8RJBUnVx7dcYnTq1hQJ2pmKB2aQIF/8pYjBxqVDIA1SwKw0
gqOtwC/0gj3n814A3m6oiaoqpfnf8oLahnEDxZSCabmQfpv5O/5dQZ5wNCGznuk2DLeKA9JUfYCq
sDc+QKAZbowa32mifK8y1hcENd13GJ/syOhStLZnOT4erNFX6k4Xza2wWv5GFElFBN9oyBnbk5Av
6cnqFtcGDHyw3O3Om5O2v0JIDfu0WjdOvwx1n535s90EBM0SXai6UHPQ1C/1WL+8bqJkTcNlfGa7
w0L2Daq1oETSC7mUGJrSbxPetCdY2jfF7U2F2kJtsOljwK0+OhYPE5qUyWEmahFsD/9KJr0/XrIE
DVMe6Vb+eK2rku3SlX8Ad74ADJtHJUzxHvJT8b8V3NnzttbhBYIhA8Np/9xJ0Jjl5CLxoEkNNXm8
7g+Jt+MVZUGCCz5btx2BUcUQdrQ5DzeYHpmZOlwzdPKUkwn3JcCZv/YqIoyBJnWiIGqQUaggVKWx
bTJVQWLoz66bA/W0P9Mn0L0AK8aVVTmWSIPcJoXIerUeJ1ZwubR/v+Pdr4Xh6V8S6iXbH/fTmAu6
KUKPwEGBjp4yp8xlx7XWCaOySeF9gMP3kL/X/qVRrg/rCQbeWoCBWpLlRitsZk3rlAMkv7yx523C
VR/RrTZl40D8NBw8rCa0b9YvWRXhKPuNaClnT0n8WuKNhHhDKifmdNqiP16PFXYuJnLhW/kAyVe/
oyOGZxrJU6dRGDtbTdUFJQHoXAFCawcdEZBIvXGxUjsmRD2CsW5ilRzj0POnDmBEvOmvKK0ytdrX
PV4ibhOGOVloswt/SZOrJKjqle21Vw/K+7JXHjg0ysvq6aSoCAJZq7oGnc2Vrqeba5Ew5m5wzUMM
aoZpwsvSWTFkp/JPIjS27fNLJinBJxmv7LXpt/XRgHGU/qNmP/+RRS/3CurxN3+lkG+mc/5FgPU5
Im4C7ov148OkzTFLREmC8lN8knJYKO/xw/AF43pl4+oU6kXaVkNsyrDck5RJbMD+L6Z4qFek9dZb
SFrCHI0UD/12KPY5r4DTvHXW18TaUpTZVYZ68nOJJAsL6mMdMGi21ZmzX91YdMQFbcGbnCk8hkck
0N7xQuxeOYsG6u9YNa9FqozN/W4DZlr6f6APzzrC+HTpyrKkVUXmprMt9688HfGx3nuM6t3JK+bG
XXz+yzU5ropqfhbiVQe75q0wUTRm8pRwdJMGMqDb3G90ozDrDR8fRX+fQkGb03Pw6e1nRGF/25GD
h+KRF7nSxtXVDO53LUG3s4akaFn8567jsk9Qiz6UerU4JJg0dI5co7zfoEWtmmosK93CkxDEzm9e
pv/+omM1ikP35nAnPQdeIKf/JrEDKTzOeHdYSOSXhEAJE3/cBWISmlRDUe/1Rlq9JB6B70D8cD7C
4adp286ze9J8+F/KrzxatwF1aQDTAvq21Dc3jr4OKHlu0h27UHhidQRPBjbYaZ4q4m+PmOupBsKX
5t4PE3KuM/FOz6ZbAAuQYlnYXd6ILgt1ofp0CPWwzKdL7tU/AAHdFQzKxqnlrcMq8etfdFHzsBnQ
yAGmYds8GOqZebh8M/ttyXgnCb03BwO0c09WnaLj3kjb5awmOboDStd/KcbXHkmU6p5N6BnCzhkz
7aeFfi7lCSnGsXeGJavDpsA2+lBaJznB6Yh0oKgsodnP269pEK6ZyT11sCXwbNO4htnJrXNikL/2
yk3eRcHyPImv8aHf9aAvv6JAC9llsGA5clj0alqrnC+TUIM45bDMVO+3yLv2UDy5dtwlArBUfoDv
t4KGlKPx/2udac+/WTgKdFsrqeFWbZiv4O1FO4LOkGnAak/0I7gKyDLiap5o6wpftkCsq48qK5Ui
U2UvxAjdPskmxwUjLQOdi/0EScIVDQbTjkGc89qU1hqY2cyBRY7/FyX0xEUxW+/UBxgsWdLpTQCM
OaQpJL6jxeXP/QSgsccHja4f9uoJeI2cYKuO8YfFipSuaom4HSZ+AtlKCvqnApJSBKUCwOe3URz/
PGHB23Z1umZ6aLHaG9OurFHiih81FMD7XFSsocBQlU9seTuw02QcYAcmPnwYf5mOL1g73XuwpsIm
I7Vp5LhCfVG4u1eQtn581xzp9WFNpu1QACb47e1J1Iev93gtR7q8fSsba5fqMKoc39EQDkhbT/JH
A72RY97dBpgCaY3HJrf6hAjq6m1dXy2unaPQPkpC21c5u8R2YYUDeup4g3eMdJQmAyMogI7JBEvt
sNTgIIkGpiKJcbzYPm+C4OF90MafDvys5rxcjECkJBqZvywOoffe0lQifhM/XQR6FrZ7F0ZMRpvF
uyXtts+Pw0w+byYcjvcdFvJO0vUXvEf0h4Nd8ik2Ucs8ypq6MLGjl4kaP5Ntt7Rimj9GgTilSsxT
DcE+Kb6MlV2aXoGbtvyqN0aZtS2GMIyAckwQINRb3K7w3yS1ZkAgfGVF7/MmhNDqNYg1k5i0cNqF
MIjZJHlTsoKs+ujL7wQu5oug0UHUU5ef0H/rGQVdfSBVnfvcqYNZJFOQ69O+vy+6GWkILLONLkuI
bD4P7/YcfjT6k96j8uTi+0t0UwvF4kRA+e6qMPWp8SNQmHKX28j/SGV+A7OGkEVVlKb1hACDKD7z
+1bQm9TH6Iftyc/FD968oziXvH2ZWkvaGsxGPaM9HjEl1vcvAdl466gW4jPl6//C+snxNwKB1Ofw
cMaUIOVD2njG+Xvt5T6PaSuL9Ty//JUtc8kun01XcRjZzm8Mfbm0XoLb389VzgMR7sDmkwTHM7no
WmEwIkZl6Ra3++DjASCyAvgwBvvc6+zMPjUvc+OjUMw9BfeE7qkrmJcg4NbnrwqtyNnkB8NFdKBt
fqM7uk6kBntsoI6O/q6tVqDuHS+IAXhCvQOVMbBAPybNI2uJ5wPBob+yBXt3/yqrnYbu1ljaedYS
qTCXkkuPJixwj/NK9KP6VNquNa84D0e4kW5rl/Ct11vG3jqycHjms05AAJYXqnTfIhuC9VVJz9f2
U2nJ/TnsxAfDjCKvN0cgrhUc2/F2T4GJaYmHa4cMA1+lAR/DYNq475qZAILtbTVeOaM2Akn7znqq
PNCiPqpApTK/fzZmCmPvj/FNByQDw+jXxCD1xy/5ysVVWcwdZkk+Dif+2hSdPTj9zlNPs8SWHDEo
7Osj0xqSgWqdPWWewQaXR3nyA+otpgI5+9/jG9Lzk0uNq85PJjAjS6CsWBVxVbVoiGKJguBPnWhz
xqfr7r/6jDV5xdzKSF+SJOClg8S9jYxrf4FiS3pAzspStbeqVLlUXE63WhopGkZ6ZGRLlKszPPRq
npgy+SSzqL9V4ECd/RAzDLLghdJQn4kH99na/ugwm6S6RAc+fRfLrtcFYcYuWZWrxhEcXN/oQ437
DkZwzPX87zy0WhSF+SpA0yB8+WmjsqsGR0vCdSiqmYCkrSlJZpZrvUuGn2r1gRA0cvAMYF6VfosV
+oE+sxEwQjdzUJb+bVtBX0J03/nZbm09LNu3JS2Bit9isPjmFbEMosA5qfJI0KHPlae6UfIlJJcy
9SfNuYXFlGPMa4i/jdJHRIqUTNNTP7pHgDryHAZAvawcjChIGVxKqlSi+bKe1LwSjn8vpcgx/7NZ
xv2MKZmIdpbDrhzmDRTJnrzJU9EyeSK0bL/Z6absxBFjmlj/KgGlRkiJtzpa33VCD6WJgmtF04oT
Uxw3Xo4OUXGp42tsaeGwwddXpSm1Px/xetsJ14VQj1ywBfsHf5r0uC95vkpS0mMaCiU+hw2DI9go
tt98sv/gnaOisxf7Weuwu0FBCG3X6fhku3aTt3y0lc80UIGNPuc4/vn7oAfW1BeuVNaZEH0dsXDh
Nr1JyY6+XK7b8Ado/VWmbqF8asIQFcLyPP/SP1iSzBBQTCl09F2DlT3gkvv4L/NKi0QtJSxSG78F
zvj7h7TgxTYaEj0D4cRrH6SNU7GBYEXK5z33VhiArr4r5yUfpDsk5QS/CC8FWxbTGFEktnmeo6Bs
+lOswUif0Gc9Iy3Hymu4AhinPe2nuuKZ5U/ekAiJE7kbZbcKe8wUN8B6qaOBT5bHSz2q98oLs9nN
SSBzEu2bIbPmdlCAxK4f33BbADqcnOfB1/4mA5XcnlDlJFKLc5EdxN3rdFDg/HPgDH/GE6aule8k
Wa/oNpvHPDSEfRsbgqtN9VzE3TAP8Dxg/yuD90Ye8KB6hkqI9112+MNhkmAsCUFvigJpvc3KY9DU
FZpnfY7RlgBmDKJiunDowic61KZpkz9DaLbDrmAW3gOsby0fQGzKTMl6XOHAWRcQE7ssP5t0kkB5
8pQYAolck5wSRrZnOfJL0IPGjYdSLFeh1MIwFv4+wbUUuGHZZ/FRGhH30e1JGn5kWD8Zwd4hrCo8
Rph0ZhMplGzbP4xo5UfO162r2y+FjQ1WRuRbKKVIzq1nIBiAigvbPWFfFYlcbtoUSqWHx/DdIaa1
F0kwosgKj9MKjUQXN3Y4bTI9CzKBtGzOwO4i77RnK3eWHczeJMY26DfToWj+StH9SYRbCnGXEjR9
BMqvt/Z0YOZENAHMZVEzkb1DjB4ttthMyMPGo5bmPyCn8XxayA5W9mz3gs7VjI3rst6hBzeY97fW
DQUHlKwYO6qURvMiP7sqPtZRnXyQR6YnXm8SU+lC2blGSl8piAZDn5f3iX4Uy1SiMkmqoOnCr5Vd
TJaRUi2s5ysPg9qCzqHQ6+vstFXxJPIIbJvgtm6BRHrkxjYNnss8YVMNYbJW/E0OaIObgkyTr83G
sssUvWQj/bygWIwDiYr/AoEPLBCXdBNvPkFgTquuwTrMIOM1USdaRnllNBXpDJh1kLBR5bBZ+99+
tzZGoJp/0nXvw+QMadoz28iBX6mwSCkutvQIT2iQuZqSCLfXizmsovaViVuVSE+I/ilqGp/5U4Op
oh2GqzlcUdFj3fr1w8VrWEfRiYBgPDBdq2GBiuA58pVHl2nzCZsZm6E4CgHK6jzAIqh1jTxCXaxO
lsKT4c8Atibkz/A7gJ3nNKBAUn4byyYk0BCq02ZBoYYfY/IklaIroB24agyIX0w+sN4wqNuMAq26
YbbXjC3F4wfHf1CVLTbUvxhK6bFKnc7hzKxe6STxuRKfyl0oVL1PlMjGDnjCrFnSB9hEpOn1GNjS
7Sf/TtdvaO8G4eO1aeNXsuq2nmkt7K5fqi7FUfs08IT76zpMjzkMmrRzdMku5pB1ZaTJd9/5sc9D
Wr9vLG2EK4hJGNQt5wBlwO6FOmGQ9RSkY8CZIHDODftLSB3WZ/jq4fDkEYdpUDTPynYPi20ELIBz
QEkSRAv0Sn5BbzJOLg9VWVXzQX+3yeXdY7+06BeDD0LQIlNdv8GADR81ROVpQrvClhyTAlzEHMFM
HSxLJdNqQm09SvV2wwYfaQMv00dQj/BQqXZlalO1JC9nebgRzyS9GECIhgUXxWRepyenV98nZhtF
reCpSkbtQ0GiZzNJuTV1m6DUbtGGPs7ati3ge5PpjYmoiPD3UfZMTGl8R/kqq42q7z6g6n51a2cz
9sE3AGK412YmxD+d6m6/iiRZ/A1tQk89jDmkhB+GBzulE5Jhaauf6rSRj0WaNGcoPc33UmrzwnYI
8sgBNmNjhyCsW3DQRx5pw6VPVjwIppPPeBzhhtw747iyV/RA2SuYWQ1TYonqvXHaOtcN4OE2BmVL
95hITZ0kTVZdeIQiQCUyZZfQuoT+ZJLk4jZR61ZtxUpN65hkGjdbfhilXKtJGphOX+lWZAvVLkpz
FJ32uxTCjkCKAlV9FAIsPwMpEjsXdOH6nuVtqY0jSseBoA/Mp4gTDlyhuiLbxb8h27n1oC6Pb2mj
WlItqS+Q6toI9iREkiUIj2uJ1fdYr+gj1MhjUs/qjHl7FQo0ZTW8UdCwbVWLXM7mOrmO8aj6lP8e
fTyZcndHTvdF3B6SMN/QsIlE8RQxee/l9q689jSozUVUZxXft7jTB50jkI8AB7z/T5YG0BDRxI2d
jIqVop2fFkH/xg+1uf4+dQAC8hgw2/VpmmnuBGZG0kQGSP7kanHRuDB5jofj6T0dWbCn8PfZOSo/
frXeR9mRHi39yHx1jCfrGk4ZFCb7cqlDM+krdXAUqy2faIU2sqym0AiiyFnWbCjBbSZwFLwLr+wO
Z+RVHD5wHQsuQbPApzNN+DYKPoAokesYJsxJjN7fRR1Sks8cqtH1187BfIeG0lBClOsbRXWnnNU2
yC5sBeBXXTJ34QBabJ1HvUoRFx0NzxFcdRESfTh6ArWQiEi1IV27347429CKYwIq04LUfTvvUL5d
6szlJ6z6xqlDkEwQGCCVqG/NbxfVMBnSDGi4svsCs2gLDv47eCq2nXfAfU1kfoudy/xrf44QDVaa
m5pBlX0++Se+E/0hReeVeESnMkO63ztgYcQlsCwyi2D6jWVRui2tPwjD1Fwytil/Fmo7sDePJwJy
YOZKRXI31dVNUMXXxdLACoYlCgW6ZJriESmkerfNmCodsilmjX8dG/psuDgure+mWXbvQYhoV5BS
dI7Oer9CbTH3mF+IU0rPChTNkfLnl1d3keb1Ob8uo+FBs44ydHnasj+Agemd7ucTWOMceyZG29sh
GSpEbQSMStQuGGp5VTOQ5dRXQ5tyr8aB9F6JLkzGGVQ0WQohHIv2D06cVWrGtic7llIobltlawuD
NACk6h4C6zVKExPx4BakzZgKDeImefDYx2+kJMspTAaftPD5L4S5dvwJEOrZlxYROEbQTBt7RK24
2rL/6W/Xi17ux4QWjbishLx2lIAs/+dgQaXAyGSJbi0zZOJrS/m9oQoDI/Tjt/re/p6EiOcKE4Bf
FwW55EGNqO7VnCDtjZ8wpEYDZJkdJkMS8aZjXJiPtMyET/hmkQ8jvcX+M0h5ZvPslPl3Nd/0F/ei
ptB1FAXf1y+/dTwFB1f6lnD7ju9sYbuyJqfQrJVkgkHw/yVjypUQ7N1DpGEPGeaV6myfpS6Wn1X2
5QZm5XOQ49fYn2SYsoun9SHgMbxb5XJIDDQX2QKnL03zQmcEe8r9dMpRBSY4rJRsEKgrf+rBXuCl
cAEpOI9Mgwifa/BVm90SmWI4071Pr1z/v6B+R9NV6WNaPNDh9yKdjZ8XZBk4Y7MvDgN/mPkSekMx
baMxkPeckijplKk3/Yd17q6+59sHk1qjKvr6Pvl01WnnGFfJGL0dOGABytIz7hGPprL7lRHT6oR0
muC/6AeVcVKU1tYdUN+C22zJkmlO2cU2DbGkF4CrdzxF8Du2CJVS1c5gOS4N2VQPT86+xY+aPEdY
+S1WbQr5es0xssPoOq/ZBDzopcNAIZ4gEROPkLTr3VoDmmdycwBEacwrKrsLIuL2Q8+OJynxIluv
nFA8avZ+aaXVULdPTCjegr5Be2TqVpMJjBVWDGbHWFQ1Ni7dy69KIKLpc1jXIBlEl1fYUPZ+3jCP
qTL6qGm4VoHCPCaHS/Ga6YMrjzDXK7vvZ97lLX6n0Gsp/recS6LLQHHFAVDvzf+G86QJWgKk9QgF
vQJRgbkv9W8+nF2razcIVU6ItH5OA2t05vqCf9xqdOBZ01XUBYOjL+xB74HxBsMi4fizW4BfVLBq
AHEmgG2TAbTdqkQzkihRmiDxLPZmRcW8Rg974M4b8Ck7Ae7HZq3Nn1+G6a0wt9XEWHNNiInqBMiv
UMJiwnAbDzCtmWWdGIFdGWNNOWQU/li8iFqKLNi+RYdjqqqIprS3J8MkjJ0RLyob72OHHdTAt6ZG
50/nVSR/mNXESzQDlQpE5KCHKqdPg8xVx3syH+D1xhuBETtraiR0mHonwj4tbzZB0MWKm51XGUzu
LRrTsFIYGkgBZv2Arc2wEvTdx9pWLnHGl457Hq+OtMVoTNWI1yp4HsuMYTdGsRE/Hp92tQ/ZCZ4e
UJuAZaYA2L5W+Tt36khXfc6AriuFrdTOSncNlGJGAEer3sqM1jmhjaEKKiKP4e+4Y5q9NkXJ1Onz
pQJp3ygEmhh0PDT4OqlC+F/XtCdNURBBhqU4q2nNJdWYjDdamq/muA/u3u2zXWx/P4dx2TTNULB2
GImhGheQtoQYE6FiC1UKjzlyyBEkLuBAf/0gsTudcx7a7D/+JtzTeiiqdA7P0dPm6NrKVny5fIfx
Y1vTGzF1Pisxi23PKG8Ft9WY/w846otSInFf6IiYgJpzT+9o+6J26lcC6QuYwlbXkxxqdBAA5h9s
12TvKhYkvVPq7PzcraDIv0h10JuchMQ8QeJRFq5nZvwixkn3yeVtFKdLtzoXrh9ZuW2hh5+g6awh
lG8wa+LRAPQBJ/5b4Bb+3IF6Tqu5mY+NbVBEOfXatwgg7DZTibG8EDJ8WJYmT/K2+2MNOTLbOUVM
WIIayZl2/f+09kkg4pYhJQbi5R6Q3fIDServwmJf2YXuQeOyfPvfu1DwM2QajuC3gMM7ERkdwXI8
IZlIkvvfPmspLclOi5QFTmqbVNu0A3s2zLK7FLSe7NQa9///QAbkZNPNe6s3rmqYmxauHedYL2pQ
20LzHXrLB3djhDTm6Sy+o4REG3TPKtpCpTKcCH9F7NIqmoamWZ0xqTsgx5qcSH07lBE4Xf8xI+p6
FetrYGar86Foge4j3UEZy6iCWYQaX21c7gRjfm4Rjwr9TURdENG1rvsLjXUzQ+I/oNsN+Hc6BubZ
AfcBdOrDknBTG7U+UK0voSDK1FoJ7BWv6BMOhkPoLj+M/rHSgf90UiVXt0cdFucJeUPn3bddWZZh
PGu4/frMpRqxX48OkCrTMfgoPgRMshQFxB+tH2NWrcbA+ZVtvaj4DakeC7+PG15Ei5Ehksdwf1S8
yE5FvIJBMVU82LnIKoACUCqa+xiCVQiaiGnH7bgW9XNrW8RlFYp45NL6UB4WxWUA3ch6JgwxjYCc
9J1CwCCbz9DzlU1YwZHx5fcWVq0/aopGwfExVAZ2JU9PEMRZpeojwh4stIBzoD2n++5Pu4602C6M
oT36dRKzDp19qMROZTYTjT2wg1hgiGZZXNe4J57Cj4I8Sr6bAoK7gTOQ2rr+QM5LfLn6nr3oQR96
jkdYITIUSfG/qLdKYkDv3Olw8M1kMF4lz+oXD7fqyfeFPGNJ8Kn2mxQR1n+Ynz7+teT2cG30N1hC
4PobLns18phZRRfjX7896ox563Pfk6m6OxurasjHCsJNu8fjYjD5s3uM2nGt6Aj4vEmCVw2rUiO3
0REs5nh2QJ0x2r+/bL5xaU7w2DZoXgwCHwfwMssMXBLE33HenEBkpYPwMVtQK21rv5Aw9RAbxtdU
81GKa7OiodToVmn84GQ0dhIT94fHQRA7hs17sfswIvB9EY2CcjaI0ghHkNngp9ZwpPnkFYrsUdKa
CBfDKMVep/sY2NfJwIUOFB3DZBAzYxOI19UExp8tG0UlZofXJyhlXfx7owSc0yO4IG8Zl1iT4Kqn
anzvDxKV9GzqMjmc45l3deFVBva56PivPPPU4GfIYPCxQUT+mGIm7+JIvASS3OdanFVGoXQQDp0j
zntvJ98FEk03vBfCT8ikdQXph6Y6p77pLpPOMwJAhv+0BJlwMGEB1aFjsADjSajolHyofEoAioYq
WT2WS24L8zKNUKx02YBnT0KNZZ+TLcC7Zjurpyb96vp2XLOKrbkr3PC1+1MfwBHcpITyYnGz9XIN
CMvUVGowVSGXyn1BTHdUJ0nrFiJOHIEJyJxG35oEHHA2yA97DYTjM46/5o89HYm1kmSQJmRdJUQ5
JKNFv+h4TQu9gvs04dE7c3JD5gPkkYLi3syejufH2l1n8LQZK/QUgu7tk4XxkjshwoGvnoX+90Db
LlVhO1XmpJ0I6TY91D9m+ofRNZYbo72NslfrapN4SSshZgz34xOgZQeBQYaVEqwxGiGEjMIYzm/J
SuWh4ogjSnpQI9usTgovFHrw2EY9D0xZCIRkg1ECXnERhZNXrmXXNOs2B/PK1Ai3WMAZHbsOTIZf
NNxhvmWP0SvN6IHYr7C1DRv6gN/VfWMqppgf04jmMgYOmT8R7i429p74P89KuvLM+w0wYMZqJztK
CV/gBzoPaXosOTq60EmEAEJin6W8/sUGmg/QcFIm8tNcbuOVJ7jdzDHOy9a4kkol0Bemn2GlJxM2
LRK0hlqMYH7asrYrNDiOA+tchtmUZszR8I7s2k5VaX7rRtOY0YO09FqlLN8X73pUQnkjRACEzABK
XHOSSV49AwhSlwbsNcMQ2UPym4xnUyVKpXW2iczA+arYZOI7HhmUtszCFUdw1IFlNHH3FxV/a8EA
rXvRkuu+v+eS5B1uGCtiEQ9j/+hefyzb7EiH10Z79eSw61bjdDHaDs/enVWqMOR5ON1RrOoa5NLO
fONBrnDvnMqYTQaSBscFRyGptmNz5czn4okNRLYjITx7ACjWJmmk9fAQHd5wJKtShnenRyZHJvoF
ffV50lX7LmQ22+75jQywET1aAUGmqLyimAuxEk7u1Jo0fZhr85xsrgvrrx0gKNPab1F6wSRtLQBX
R+S4vBS+r6y95mh5H8RopNMXVoMDRMCnRZlCkuB9JDP25ITfjndeo+sdu0YnpPNtGpM/hsPutFqp
2S+ZwP3YmvqffVBiC3w+oR4IH39MyEJSGBy04EP4ybXTMROFn/YQjUBBtmvYpnods5p7g0PTI/UE
dBX2Km77zqcdq8lXQceNgR1s5F1bNtKga0RUJt5YliEfPVUVrUcOndbjts3w7oS6ZBirh6uJoEgJ
p7nnMqD6/cap819fSLUg6C55+Tduzc4kHcFA/vrROc8KaPgNfeeIFxRUm8TLaGF7dYwiGSiXYxUR
L9UK2zjucIfNN6TL6aLaefKfT5cmgrV3gZPPMSizwmBCbH0CEVS55MC+Nmy36M46poeP+aZtnv/q
zrc1ckP1S5Wj2USTQT14sKUqYds0EDCJKqu+ibhF4jld7g6RAfYQyRWgh9zH7AiiDGKhIp0O9ZtB
ZAbov/duBfeizh15lrwgsbKfT7RzFiKZX/lCQ+eOTLRKA+ORbFab1/oLlW5N7vBnDFWyl/XnvlVS
KhgsP1F2jFY/SNi8FEiL0BA9i3ofy4dSxHPTWuiDxTgLLo+0czvp1qqDFWx3yP/U/hKatejme+bb
9xdSyAx+FmtVEnLZ/sRU9wsiD+bJyKmzS7CLTJcj+bIFoDH0iNWZxAjKoFHiS9cozFbSMQ4wYhp7
+XMIoMCs7OwGIz17jqwYGR1Apuwt3DtqVACOBGnB7YQMVVNQyTfbk9MNdA4V0VZhC/KYYDZNDrp2
Cmlcg1J2wIRR6EEABpIJPsdSa4NdJjV4JGDMM6BL9Ab+85tPfAPIa1aKSHYUQvc/pmrRRJMzkD2p
AQAfDApcnbpDQ9Vzpr1j3XACrMnV9l44eDRqU5DXXTqdmp1kAkJ/ijcG7zQbvPB6F9GHpzgSTmI4
HsS2z5AL8G2n7WTWjKy4ZXwytAA3av6XdXqbUeBrOkTEd2z1XxmuoSOntxaLVJ3pwLgXASCF7ZRm
v5t4v6+IM+R2j9pwqTURl3Iuz72tCPXo0Np4pP0F41sPFzMLlNP7ivygZdjIqEZT7ahaVNaDdfbj
xZEoXOBDbXNPJees3aHqJiGOeRFnG/YnXdeM6LfEoHtxTQRUAPqPSyhoZZ5dLM5mw3I+rOh3S7T6
39ida2UlrwQC0pRt3/Rsxt7a3FVrJnsWz3IgKx2vF/rjNKo0CsZjqvOxP9QajMJF+X2koPbmOHdA
9398LF015fv041Ju4eCEw73Rd8sSI3w1H6e3hC/fdAQyPM+MBQaS70EMvpziaBV+nDYiBqHuOLW5
B0fAEtS/3x5D97rlHGPktej7vn5CwsefWOG11oZZV5Tm3yl3CevUJgRajpMwmp66r5kseNZTQzCf
1h9+S3YiP14kiHlOwj21sfYQDq3aalRRxKrdXrXpcI6u7fWl25l1EYxChoq+GdR/oOreZaZeMLL9
ZR0uTwoTyGxQvLa52YTG+qcfDCrw0U+vnGuzvs7IgjCFn6UzVceuH+zHH/gFvVubIZ8zgCRM0e7j
ycuwdV8pfsL9O5cfrybt2s3CS3E0GfqaAjB4VkSOyKR+JlkXRfMkejSWP//Hw4IrcLLZQEdietN/
qLJJGsJWmLQ8/5XUV4JWXCHX7BduIc4c8J/2soUT6uW+eUG+MU8INhEkhS0tOrqGdzejKYbuArJ1
u4qgoaqPtZpWN3L9u/AWLmHgDFwDQkBmwyb/i3HhywyRWN5JocmUrsgSqVfAWRZ2MCDGgZFfSQ7v
g9qhYKg6mqJ1MlaBxgHRB75De2L5TnBxrlwMY1/p2pTS+AQOA62DggPV/zwk3LDPHNHv54+J4L0T
OCzfSAAl5g6Rq/6ai8ErNmjoYSCWxUEmNqKJ2uGZ/UsQ6cDVHhFl74GEYvnXBZLuBubFVyueR8t+
mH4Ihmfv6gcX1h8oHAf0ydR/9+8KFU1/+MVHo/40P2uo6K3lLIICg9+N40OskhQkl1eCI67/NJPE
QbyJeEtTuLhM50KfmlFc8xsV6PZJeS8XBLG5DRmHmWayi6yNf/FBNVjpaAEeEllLIo1thDwbTA4O
QAmVfG18vs5/XIzReVLGH9oK9dA0dJhzzM/BRZm/cktDl78vAmeS0tv6w8rqNcyNXF32qwYOe0/F
zP+hsGnHOceE1Rz5gjmQCpc2w7uwa1CcsbnNob+XlN0y0EssXw6BEmTYFnBvDYrUI63enBdS2iV1
bUUDopVR7yw3MvjAIxBmHz0yVWogYRXPXX/s+Qphquy0oOlYAPn4h4/MuR8Ru/64J3UIwTy/21tS
f9v9fQZ3x+KJsr7asrqkI/rzeJtUTaXZmjPpOAg8x2JKDZ8hx5eQA/3mA+1Dn3CEzfegvwMYLa8N
lNmJxESq6AWFdWUsamawYvUH3GNaB/W8UGUVqaWdstg4p1cDJ1yon6LxW0F6NDNXchiVKUut7wMa
Xs1oUXhNdbpUGFbqweNWVdr0g3KJef1lCf/Yb2uScpMs9mzJSZHv6Uy9IL25t/Amm+9GC6Y+x4N+
YNkAEjwsgT9sL4Pombx54nU7NpjgKKjaS8JLhJyzedPjYG3X4aYBUdghiZOw541a0N4cUmM/tmw6
12TPhBbZpTJi8W2r1FSIogVcY/qSGV2VlXeeZYVZueoRa+J60EZUXwvbbGILUsquM+OWDEGdes6b
hKH7HbKPkUEIFpbV7jT/WE1kNP1Xz9BkDTgnDoamlVC643QjW/dm4QXH49SwH8I+2pO8q36A72ft
laRMlO5pdYsoJeIeMSNXCN1zMsmU5Fv7Ecn3/2G4BFArViDfXbLyt76bHp7lyUqg01xrTJHwbMrr
QrgOaHQqaD4b9zB0F7uMe5ltEJVHMTUqxDfR2CFmW7XNNS8dwMgTEsG6No3nJ5pV1/YlSrR0Qfrq
1STt+74s8NcKEm3mROK5tfiLur/PHoUUknEAeGSEK9YVpunqudiRGE3zGn3ya7vtcPmdktY9Qx2K
6hSSuTS+7LYVj1VCaBCjMbytEfxkTdjYjn/iinv4Fkiugp2Ru9X1dUZLZyUEBZscdYYyoEKa9zi8
BBQH/cDf2qhsZ+8YSH1hNnfLj7F9jEazooCznrKZF9iLbvfP2tSX5unVgf4JDBrX68aqIpzgvDgi
fJJLpaSsr547IBJJwuDmwmTizHKOP+1uq0a5kyj7NYCJl5jiL9G/WZCTpczFlpojsr8JwPOdVxD5
a4BydBchzG8MH4r4G5CHOkZ7vS3+Z6R+27QO49hiCPRBOCsdH2eDODhkV2eyIDNggEEBepwGq1pu
3i88FtfEi0AA+++BlyFl317VhHNj2OgdL5YmjlILOE9+uVO2nxltWXDuxPcLF43Lqb0OPKnXPCvn
1fkdDOGBDAkMoPAeh6R77qx61FaY/OYYcAPUDX9diyLTk9aT3SyhKAphfBj+SOCArBB+vlGr6Oz0
iLL3PTACyWp/gyYh1VPS9Yi/425qU/ejY3tl81fEgTmYRMBUJE1gPguYT67Y45JV4PtzRnVDKzE7
060awR14ke0dxuUbOdtDu5ArJ6JA3ZG86u7EaknkO0eqpCN2T0BKJ0E+blyP59DpdNeO1Hy3ZMp3
Kh/wizq0zyC/Mjljr/pbe5ss9EDm+bOKGwX/opWiB4CbKTUVg41jI5mhl+NXHgFFgnJFLcg/QJg3
QgiMvgnPqF7ThHnmWPhIxGdscjAZ6GWAJTt1pt3IM3nGT690CvNwxSl2czBpvDh7BBObkxPkutyg
y+6cXR8lNtBO2xSnyAUa07NR48HYDCNWFtc2+toDgTJWRj2UZqHr/NNricpZpufo8yw0CXWfvnH+
mESqmz1pVU2rvjSecVM/R79ppsRmxUB3eqp7ySbeaUsqIS3rAZEWL2D9za7Gd7mYpDnBaUgkZpdx
r5oAVnEgP0WhEkRc+0jIAtjykImpunSmGLIf877b/wdoH1FTuKn9eOtE+O8fWjrVTex075hn3yvT
+k94B1FvIig8/tS7AeMC6nbUw//emADdqGGIDVjwXPQvsbVATDsXuqoWCtC0dy/OSc0PeHkwOd8R
cR3sbefQts8ypFX3pF9QjnGmghDRE/eYXecrseL7vw4d3oSHOzATEwuRlJYBqYgVKa/aFeStdZRY
88qDogOtG95HpM2lGpa+d/0Z32qwF8r3GiLC/v7hiOvgZMMGcxsyEfDqBZLqvtev8EzmO4kGJ3l2
QG9IMUlUfXPSLWHMaW8POdUHaQpl75ld1cpiReJvQYDzRh8Y83qxa8bLWxCB1H9NU/pcf35OJWPi
7j0CqM9pOS1WlNhT+HQNWO4cTfGtyPM1VtrsEVmAaGCnSQ5wSP2T/tabRscIPh50hO06LiRDfX8o
6RLDj1JzYGtrrBch9G3HbPOM9yyUP4Lr31TIzDdBBaTohXD72XOFQA1ipJBl2KV307kvwMrfPmiC
WOcOecKWpuI3HZ1P7d6hrA6UAbqQVC7u7q1mWA7+L/4aXRIY2xK5mkdEcTBKG2jiV2O3HmTbA+dS
km4t2sSwgjZ9ceWZ7+1HBIzrh2x9Xoz+xocIx6A61Sgh+kAdO8uprjoSxH7aoJQPP9Bmrk6OePfh
foWwmKGSolIDKyso88HVzX/33f8BkSCoyD4mcTUdkjz/0wxkTMf+2BK8tjDMmnAu6rmwuKdiReGy
7JdUjGiR5WpT3ExzLq0XN49/o6Wr5mfPy9pevT4TdVrN0k1p10F5FSNYyD39Hd4TKH60QlWwD9Ad
9aBs8HTAM2f3Qsi+jKT23JGXdB1ShLe1b0Se8aFnsJPMbVJLnKQxzHJ5Zo4+Vij4I/kh47vrPyEy
omak4th0pcwPGSAudTgf2BPwHdbI5ySpY1Ah1H6asL5vT30DkfBa1cuTqPU6W+go6ZI3pEnYnAVl
pWCK62To2MP0SftOH3h2zu3lii/55qcAkZEKnZdcGAOLw5PLZgZFbicLKUP/0Wf7H4MQY+xbngID
aWHEok/P0xlLlvSRi5o/DJw9tMpgbZf9axPSXXHm1z6JGlXL+R9UhDYBsW0iBi5WGy8WTijx/M/y
ru3nojRiY7ASJRAmkDDYpf1/d++jvuKTegQrGZaZEfUpCAdbCL+AhaFHbY89QVE0TmFutQ76YB9c
pNe5Dw9IsDPBC9PRoUO+/CGjeXER8rICbOK7TbYZuneApUywdvbthsxzucnmY2TNHpQiiQbo8jK9
CyoNvebOoF8VYV9xvAab7pXwJAaUH9y300QM1ajF0QwhG1EXaGU2Hz33XB4BgLe0kjs8GxboB+Ez
N1qrrMzahzaqnJF4PxDmsRWA/oaDD3J3h2jQ2mrfXNlTMDrZNwAUYU+AeQ1QPecDBNYnBOQyvHV7
Kap9oMg9vzdnSIcxdniO5pS5QmG4wwsjc+kRlBm6Pb28d4OpRfxGLtdGhbaw2gcFeIcfelBvrkdO
G3HR7Mtfw5zrLQZIPRGw/xB5UapyCKmd/R0phg5i7WGnuQPetdZ8NP0kX99y61lDH5FJMreefxxp
SV4ls9vdqKPtj+ClECd/kGRTO2hC380iABJd4MMQInvG7owRYah507dKdQyWfk5SczlHjIXaG+hj
k08jlC6LGbUNE0MXeQ7y+7Q92To3Wnz/w6WuJaKuxpJo/BgJ/MyOWAmjlPm//2bIn32ACZtPRl3R
4tvFaj0NHZHyhwXOr1ixuHVPzyKNrgfdTv1ogXa9o4uGAFdEuaMZ9RXvzdFdVZ+nmycMxilP/wz3
fo1uQ6M7mkvoZbyHwQ2hwzEWRZGYSptveUmdiCTRFlzub8St2FbDB5/0ijjKXvhmLiIUgtLWOwmn
g80W8fFhCzD8kTvqaSmwCc4QIcnpjH+SUKKD3awxqlS5vg/UjblNo5P+4RD5sGWKwHD0j74Djbhr
9VXC9aTplXCLB4MCuOwtLwHuK/33hS+uTyEoOT5zqi+Qn3jfCSuExrgyiqfQ+L15nCQ88L8q4PLT
jJ6yI+Clfk9DzYCwoyOLgRUSMAYy3rZLtEkdP92U6kEmYGJ47UsqZVTDWAVM1z2l/f0SVpE78/sr
6GvddCxy18saDxl6gVYISchsZDQ01sWG6tP6nRPp81kYppF7ZKPWG8X27paa7ma3HkTPsTJXDjgR
Pbn82DqnPpbH8ClrCd+a4CHNXY8MyOsgrgjIxTJ9dvtyLuzlKSxRDGH2nNohwT6JM3lvC77Q0kZT
rVESPogm1blqwYJJEaHQYxkCNxKd88hos/bQpYOWF3OfRjalviVfPHtyOwcxE+En4EcotRTIyB1F
GV4r6A94CX9CPIVHYezRklxck2lU8KHbOgywNOVRLJrZnvjK8XGUziLXOWnSOim+Xh5mcL4N1jq5
97OSb35wFtk9PonZOF+fC2LSBYjvmwrH4A1psKMlDOBXc+HS8vqe/AbcmY+0NyEHy/+Czj40FFNc
LF9LXh5t0HamxuFgShM9ssp43/VGJWJR6yAHU8CJFu4p9UAnwq2uXhOf3bqC+H1H5cykEKr/XlV9
Dlmn2zQ1n70LM03/UMrVZGuNMNAjX2VXucxrbjZcUZEl1xKv1id9nplKo68EQ2SG5H7GBna3jreW
XWLg+cOigsyMvu42fgDUVmznyLdRPHLeyzJedU6FOVLGvYGHu4e77kj984/tiFmVwX/nvzR4u2yr
GG9w2UPtdMBVAibBKG1EnGii3gJ6fQJhisJDAzQWtYEtKns1CHiwqwsoBx/ofHAhgXGuIDOGNHAP
GnRVu12D+H9f0vSOFZ9Wz3L03F6G6KIhUW7bwbQfYfAiIMcvh1pIDOVrWjC7C+xxWo/9BwrRUwij
w5R/ZKGr1Gf31ZhuU4hN8e73l1vv8iVDGStLAf3AUU4ImLiMx0v1J3v9HTfe5NwYqDBx5nooNuCk
lvuJ2ZpOqnHqZcILxcoiHXu85xQh3jq8E8vhaZgpCmqab3394CE84tpRg2bB5CL22GRf27d/dLNN
WFcxSnC95ncRoMdvZs2h1FJ1hcVM3ouI0o/v8mdTxPUc4RB6EXBteACFG0QKBCCcJuoi3/pwWokw
G0ag495tmamx9oYU4/+t8wfIFZToFCUxQ/NBi2nfk9DLWi9pevS8betVMEkULwWTMhQXBePKXsia
Myuhm5B4L5r63dUzuRYnbJpE9S0BWhorXVpC3C0wIrnjqLJmEtPllvgnK/A8W+yqi7EqR0aeRzNf
oZZIjQF83AbePg85AFV/vYWIge9FjnLX+G9bKV6cAZVOFioL1Cs+N8F9OlUQzqbTgDWYVf2uyWHL
SnOfzWKUtnxCDQUaAMqEDvk9GHaE3/lnPTABke2Gxcm8QRN92BIjeWJj18WmlgR/J5RS4Vw67AHR
Va3AlSp0nz/PSi3fZ+Nhql6p5BU6NBXircOumCulad5xdvlNKt5J2NM3Hgcv8McRp2KZJ5CtFjwf
0EMMLvv1XEbYkYfVyxXY8uIHjis+cnSwK/gQGEt8eHL8QlANTNRqwuWxxYBbPEmlatDEt9j5tfC4
6AfeVLuBYDextJroaBgTmqh3L87l/t3t4CQgOEau0/HmA87jDvCpKRiDTDbgRw0grbWM7UxaPani
4TB5hEjlekHmBL9VhlFe1Hgrj8col2m9hHUU1SWCec6zcadwRFZ9qvtaLegWMNvXsSd+CQnkgvTv
/I8ZUXQT18S25928dmXZiFdaFodCq/CCaM7FFCM5Ry0ARfFlytarOYJEDv5PwnslH0viJYi5v4nU
a0Jirz1a7gtJNaCyd7ceC0lUqwHsb/NUvksQfIK/o/+yfUdb1lJCY7lRKVZZilN8dR5oHjPNwGmA
/xzI4LID7pt18jqaEzw/QB01l0CU0fOmWghI01n6JwycEEortzpoP9OdOz2sZYTwaDCi/COL62Mx
ghRlG7assO/U+KJafiAiFL+FJMqOgYP4z7lB2RhaWVbOJ9tBzMRAIhdZSn/7nmAfGaheAzamEfXK
l3yShxwFFuPc47JjIgQ8AkENrl7vmTEoBlgTTkfggjyzB/AyqXedFat0Xj5cSvL/w4S4YjorUNW/
0QP9OTKFIxgqUfug7nbuLInkL9mJLcLG2YmfWmUVRAprYcTzI0i64iIlwUsECBbbDhKQxtl7cBqz
KOYRASgs4JdeZ5GePNd2Igdx4c0JkTI90iKGTE8r3Y8YJJjT+9F4UKVS9hwY78ZVrTPeTo5JDo2q
9YPGvQdeiiqTegZHU10CVGqbAaftRcvNpq6LJX/+HXG1Zdj4D4UNQFlO3vFtTXtY7mbSUqYHi4LO
BBLZsTNLvGNUPK3AoUCpVBS8Z9B7GFIAICcGYbrihq1+Kdxp8tuJ2v3tSb2NPQNdAEa5cScPArAH
M8bZMhcPBgXm1eOHTS/iuyG4xUe7WuyyEBp8m+8hOIoLcWQgrW1tVc9+C2LFF55oGcfMar+kyQh8
gShSFEnlrAX8juuzuHZf7l2eFIK9phsSso4nCU81bDD7VBiYoLYLDmgc/Gmf2tQUJj5awP3zgGb8
zKecXCSM3H3ej2a1l851qLf7IoO4ud8TQ1BOvoacngAehaB9hQ3uVkUl29ZWlRF3bE6y1GyI10MO
m6m4hJ+frgOx1mUbv3k+s7r2x8+z6G0ycQwhAsBymdJqy0xV7aH5qkuJCOXfmfQRJpN/hLYphL8k
J0KdKtwGW6fNRNend3e/6L2iazN8lKh5iUPVD2+4u1DOK3RdRiG4oENfTcGTB3QrURNasPzPuVr4
8yU+foWTAkQDkwk9ghuI32TfS591tXGY8IDd0Zqo1EqLBVJJHu3dWPD56WfO0q6OevlMu1mr7Umw
3BjH9mBQrlmjIzbXaBIiuLvc0ArVjg7XLCtOExoHAdbTCBVHwxQMWWvR1C3AOMUUTHUNl1kZK9KE
IrHUPIJSya6aQLzTAxQTdy9mCFc/Gbxyxjlb0VZvgcaSlcNsl7XzLQwYz475R7XO3VdqJYmq0Mfy
zqN2gmj/T5tvSyjIqd3T3AHSfKtNmS4n07hwqnWhQy0XR6JhtB8CYHjJZ3xWApZD2AQ5L56XlT8v
L61HNXGJx1ExxsoNjLyanhHic2/QRcxCASt6QlGkfAdHRdXrr1u7eO3A9ir0jj9sdQUJiZ0iPmGR
0X5Lg+/kIR1wBp/lzkMp1qYKT2EP+zfv9HAv5SkSs03LWu2zk4z6Z9+a6fkPR/c99I5ZiRoSbk3m
A1LxtTZ2bCmj3L2zcdb4XvETXC7VTQi+u0FG/1ML9d+u2zQyCPUx528dlgs8bbJ/TAnSfPb6TsbK
df4Qec6jXD7ZKEIVgt39PL9DPNwYEJEw3DHfRqqn2ipRfiSbVxtForydKfYXhbBzslzVXeOzQ6zs
+y+xKSqI9lxFJejlFoR6FgPgJa+wT77H7Gmde7fG0x/EvxbOmSqroGgn8VX8QwZihie8aw8jaj1+
OHFDgRrkEJrcMfB7od1wuccOla63mKeIY/aa9ywHrbAZPX/sC8p8yyM5wO2Zwy2tFEncoqncd0/W
/D8BZT1lU+G6d62uai58Ya9DDZkeuyQwDGM5kDhRRZs1U4QXaz4ntbpubSe+p04/Dl9Dv4vKlf7Y
oRO7lvCwmHLxhgdKpW57kf0b3SmuITDwHqPE1t6ByxSX4X++DlNNenRhGdIKlGoJ1Ad7+xJEILyg
xQWsxhAo0vLpo0vUyg/Y1dFMwgQJcHwW1+HxWfm1/s52KXr+hKP8A/rdAuTcwSK5a6nCZii8Apie
AqI4QYlpiYiToaXZNv1/hEzLNOESh7lY9X5j8GwdZME0DUt3PZNiJNXgF4LWvoMdTdne0iyV5Cbf
mP0BwV3pTugfhTDMUPz8NepbI0KWQjk05vZYSNhIxSC+xQsEYMCap1SptHzX23vGfmDRmoMebJth
UQIz15Eeq5Zrxs5zxU7skW6RH1MIQrbtAVzXj1ljR+0IRctB9HQIUxMAkwxklQXvtCBxkr5zT6TX
sy2UICbYXBGQCdWZE7XnIxjXNexlejNEfdMdczEYMPN01bFgip26lDBqog2jOaZFlrQQ74yxiVTP
PwIAUNvG7VaCSA/MchmpaohIy9gkzAUXUyXzC+zgM7+6z2ba1t56tjIdsJW3k/as+1t2BgQjUCGZ
U/q0SavsrEVKVv6mOLTeUJBDb52k6ON34SUrDhBUrFso/qwBYG/Z/LjPbuFOgTXDjK5Z/tgMjkeY
STRAuA1XbnTzxMtuAvNvhsPEFG44tZSOdzFNvLgElwrslORWfbkm3aPKLSXsKkPFCb/gBMjxwr0U
dXBBbvxOgvpBs4GWWC2lRCzzYBxzy4OKSUUS6caRxiVzV9Fs46mMfURco4qUt02pLcIrpcejv3U/
7s1XMNF77/uwSR5vgeAhZSBN8GS7ps2FfulFI8kXezBp41rf4LiM7C/mihjj3AV7ZxGtsgCt0BUU
mHAz/q9vjp1+25kYA9zwWQl00jsJWO3m+/OKW95cJUYGW+pzwCfPB69wwC0zGuBhbInBjUHOJUGm
tkbOrpvfBJbxx50Cla8XX3qLJgC2Gq6s1Oh19Ij1vgNhC4Cmoj6ii/U8BhaJcS05llw6Xjvh/eI/
7Ey3XVAmmroPKQZFWvYwsw8Uv32opBlfc/wmYQN2FzAqOwqqFiggifehR9QnKT4X7PqjF6wNZo6k
oy1OtZ+HWHMWEyWdEI733bBUxTIzTKGPu+I9pU2W7qdNZIfrkC3zok0yTdgyZ7rDGPtM8yVRiuv/
E9go54/WNffgUARY9nhqhVcdo2VpQYUT9dkBgCVLZLUVO/1PCuAMwUgCEzfSDA8qOB/cKYJnY+MT
ICh0SXcKieUEWEz2U8UtL8B8wutGlJAAJqkTSQPKRnXAWzeULDhwDH/0Lg+roUXCPi1QOYhzJZBW
O4DgMrubF7UhvU8pi6X9QpxMZba8Gy4BXOKigjk5EXr2Ty4ilZTFa9WGbGyTncZVYSfNk0mQ6AwK
0VjNvomXbwr/EsDegEjNaSkFfLZ77JBdS3akPs/8BAoVQsyXSTaTVEg6D4pHToedFVx1DYsBbdrH
oGvmiLUT3ayG9jxMPrYgbAqZRUgPybA4SbK1CEUJqWj/zCOdstvnf+pSH3/m+/AE50fbUVHaMdyl
Tc1A4GmhnDGvx2vflJ0ebzt8zwZarfw8YrbZb/sRPiGtbNzt6+ya21FXm0dSo9y2AOP6R5ylLBmz
NPBFYmaJeB68PEcOWLHQxLlKAMaf+2pbidZahhmNUX+iaRp49IX4cxE4elbk/WCO/COMnKAwxc+1
H0mf23xAeENmm/n9b5FA8NHKf04kQIyD1vHbZbWcCvr6lL/2mtQGO8bqIEbnj3bf+JqAvmGbEg/f
Kpz/4k3VyrWAEfIr+nBMatTx4Yj+4w/8TOe1/Gt/u0n6QFaseAka2joXDUalOORRxNaAvr6D/fMm
uINc+17W6u39HpFhP7aSqZn7LRtkMaHDtPeApplzOiHEq7MqYAoFzAM+WysvFwi1jrTPOTManEb/
05S3H2CFcl2M6kCx3n2pstD9AKrO405JlaZvbyONi31LosUoakvW+5GRxzDdrQSctuGZhmGIUldQ
F012vCN1znYoZbofV7zaM+3j9QecUsJVQqLd+NkMp/9NnQaVG7+8i+vL5DVi7Z5KQN/mkVheT/eW
ly1WUS/sF0oiyJDkhevCQ5i6/mrGEbZhoPvm4zMsNUp7KyP8VSGkIve+jPCdpmuOZPdQFT9NLAW0
sAGTkRyFz+xxfHG0bKOs1yceLw8OIAwxjW6lInShWO/bjtYkCgwR0o4K1xm7QHkeAIdoCrd1C0+k
LLNRn68w2JjdMyEBqcz6k92NtHUU6u3eSCjGJ3l7v0m0f06HOWXAfu/ZKR7X07FAqtEWTT/HJ7Fm
CbtnZBiES6PqVc5x2xtukhEArtpAO/BPPGsed1qEbhwPzuYoU2LKirAerWho/wKubaaesnSzx1mk
FsykbMl7UMygaYwyl/iYmknUHpPFo4o6Wezl52u9e4PYr3A7v8rPSIZ5UhXj8GEu6Mqsg5AIExxD
NAiOx4Sjthpu/9g9yPW/Nc/SPgWEwVy/3xNHY12STwtv42rcbsOXsZy31PdZCUhqpvWRNkefuLx4
K68XjusjbdsmjQJe0rAoFAA+CY+i7SM+KFsNspbctL/UuCCnFtWxtiH43jtXrMNgJQGRAgrhGDat
8DrbQInMbl3z2MayY18VTXNc1k2V6HU00jigAO4NuQK8f9JeU9lxPVj6SOL+7GZRUzfSpZtlCQgH
tjhg9O4xj92tOBBKxXryCK2QkQ0Bj1eOBNJZrWeWxWJCMLIZfBRdZYZ18QTM+0sqk01L9nuNI7AG
WbFLKc6ByCGw0BYz2wUEPoRY/gRZcD6IHme2Js1yydgJZ2TWV5P1zKTAUBjaesL5/NefxBjG3Bb5
hqrzM6A6sosmC0g34PIPrb+vmqHpeHkG8H/HLPBn471xw+rYLEF04tHInB5lTCDKJemVb+vfLJXi
rdi3GeHq3Athkm0EZ0YdB1Yg4rZCsC66AmWy9Wir/BEz40Kil4riwbZJtOtwMNaaSklGPFZL+kTc
JKMLajycOsxw7WCtg6KjN7yqftTrghwm8VaSfaD4VUsI28SyVFV2P1vsaSWDT+K1nmu5pgi6dbMK
R1BqbJoqtYhq4P8jqKMKaBDQPbsvMdBxaE9Wp7ee6xfcmzIuWLV3obqHjsXkEo3letpO4KSTtlUO
nhQ5GOj/gUj5N5+DXaoMKpWDuekLPzrJsfo6aIQhviakrowoxbxhdHvDezOJcWI6wtxBCyLhn2MO
+HmnE+nz15ZMiB8iPGGVI9mhwhF56x8HcMeJGfhbb6Ge8RnG1/7fZnv4dA/kPCnTvFQYwKrs4i2d
CbSjyC43CLlb1tRjgcjyHSlO36VZv4ZupCKh6e+fSNkOK35d8uR0LULZKCie5o4Y1GOkpwmV+VhS
Pxc/bHGekyHLkrFGhNccZEg8KAuIZRY0bKDdjF9TF19p4q27GJUNL6DO2KuvaTXPAlDLGGIT0/2C
cbRhUQ7EgYNoVP93C1wSv+dZs8DThZU5Tt556Vji8PY//OsMC7eEXoseruCU3rzxUankkyCqROzd
QzIti170z2DLS6fZCgk2RO5U1+7IsmPd/mLa+as5izjwNAGpTET3w89nl/QZEwnaHDYFxcfp1SOW
sLpH9l/DdtNFfzj59elSQNEXSe9uaZTH13uZRyyQ48OwZaIB3OiXdPynAqKZt7fAi0MIC5f5NvL0
fSKqyhAZc+K8MkO4DMvGkbTigIBIi3RiXz85rYg2iWCUG/UmLk/0EpHu7ernGB/qGb/pAF4JaPaM
gp0RthdXDUY4SXxpjc9HO6tIrNkn31YIXKKFzO0UDTQk8WolHOnp+vnW3MDm5v9A6NYLx9ADcLGf
NiMOFcRmg5NlHjSJc4fc3eNsV0+6zH1ZtUJuZFJ7Re+FpnNC7U9DNF4Ms8yXZH8pawk6yPtlbGbW
S9t+rOZGJr9t3pi3bqD7T8vOCwvUvVkR9V6cCPMtKGs//0jBCQimj3MXvsJ5fdGPLw+nlF3Oguw8
ntY3ZPQ+zl61SYSskf4Dv0Xu5o/JUZKEcPL13BkU958VHZq0CUEeL5IirzGEENt3S5vMVlfih3eX
9H/1KsKLc62XhjRytyEYbDt9QKUMmurTvWTY8mPwzixrnSmkymyrDm6mU+79yI7I6WrOD7S6Fe7L
ct5+mW3WDqEZaFAplMrLuzoQb8M/PIskDtXTGdpwGFiVwDjsBiTcKPeqx+4hUhs/9lPSxQc0GSli
04xblWOrKaEkJt4UyIlzGiVA5Ty7h99I8DCxCa8rnPiWPEe4nIsCAOi5H3oi51iDV2yuE1R5Ki3S
+btJEgfOAGcDCPcG39qmeWl5MfA6gQ2izfdZuPAmrriY1OQDbHkzc5F8DjzSWtum6pIBf37y1yrL
ySXgzYx+dsjIxa7OcS4IDuaO2A48fJ0JpBdNseXECi92rRJD9DumLfbo2o1PtnC7lwH7n0Wp/coR
UqojFwXv9I1Q9x3lIqgVP2UFHohMeOtsdBNeMfILsT5sIBi+4Q4h74jhAVL0h2jtxPGpgQ7EHZIc
tc5h6pl0jja12qCYEVlNsgyglwXeXfo44usao5crQz/wS6xBMqgG8LXBP47fBjnaUXPrSYRHwkVT
kuc8fVJz0iLxRNvlgEVr3gKjkFUZfn3WKdjCA64/wzBTr07ftvvDfAiAtbEVB3tTZS1hBtHuzOQb
Ly5NDtq0HfRsLDR1RiYD1USFNpn4vziJxe0ACjnG6XIBIrodN0JxNHZMwVfWsX3+3Iu3RIp8txT5
Bag5R29X31dhc1z87CT1awetZ5Kedy9DX5WUuiza4+0v2ok9zy5b89z1Ed9u9CL7OXuKEnKXQD2D
QmANTaUXesMqD5z+70UtKbjVR190mgIQmjM2JlECGkQMEsE+0PQbmszEiNsKEhlpoTnBl0C2IPSl
TLFZr7patARmf5lizdB1mkc+VAnKOTzF/ow5sNuVfYD5oKYlaxF4IT75azmX9XNeRm8VDpf0xAa1
YCtsT3BdipSIWSwIzr3OlpRPUHXl1bmkeGqS4g/PwzzHBIwa4yqZ+ggFe2r2iEUX5+OXUEpaaH+7
1hvZJEgHbtv6bllJJENNwSQZJNJPSPtwADImkOKZN1on2LgbMhhUNl9XZUxgQm77v1+1s7A74WiD
9sOqc2p3o/4OsPxZejuu2Ve4uDsn1D/cThHQjq9rWzQFrSyM5XGW4OboUVUd/3glyZCl/T5h0Fr8
vUr36NljHH+sBB/BRdcOV7FSKSyYf2PN1a/IVN8zgG6iGL19U8lYtizZv6ZTZU20A9WbBF0KSDJe
+ry+oR+D8BttpLguDAm5hbhtHQgitP/dcxM3ReEEmB4jezV485NWpU8jEObg+lMLkiVdPKzCXqib
B+d7c5bAvNZMHt2lRKMjmToC2/dg+oBgyb/mCGpj+byW3pikCzDGbXFeATk8QuyL9CyvtJCSqHVw
hk/MWHIjE6m9sxk7xDcljSvnLKndjDBnywMo7OqYnxxy0uLE7CQVC8dfwjoUtRr0TUUyEF9XlcGA
iRCxFNU4F6eLCYCLL7gbjN49XDPSvtD0L4efCAUUuevOzmtFnbqlkZzIbwZx0lVwq4+7qsPQQzE7
eqd7g5GXMhFYz8ogyfJTKRPs4lDaAgJPdT5xmGnu8xvj5o0yuq7h/abWfFUXIIRY565vv6iaIbBh
XYaAaNmFq1n6BuhipcREN2axTZ/MBP6nBZmoupB45OQrhePsjMuACZKtZekAHeqvdfLs2ZUXhAs2
6Fa0cL7QrS2jCcG8vAqjS1VFVBxXBCR5IEEEYC+L1UJbBk7Q8xB7PeeNLxQz6KaeC7nJsrwF6v94
KW2c3fEqRz7KcG7kr8C0XU5W4NB+6cx5ojJ1sKwuYnVL8SaLIvNIVRga6iWdU1tFdB4xxITCXvZX
wZPrZZVGtj6zH7Wsig69lboJB3nhVChRTLg4fZfQ+9Wg3LbUwOOPqFCBx8wpvfG5zcAGQaCz99KS
/A2zRAZezPcCQMOL6Ock8O6XyiXzMHelGk63BORzZgcBG7IKxFAqlLM2M52XaZTF97a/Yo5IPEmw
JyWQqsnQPxr8PDuUH9CCFy5RxbPfx0KTuQEpXOzwN5M3I7APlO85ZjxZvBaoQ1bT/yEPA2fXHvx8
kROSSrqu0h8Cch7iZmXSOF3tGOsm8kanJeVQDd9qB77gZ5Y5Od1/W0UJB6c3uJPNufnmv/PlrSfq
zkm31kWw2mbDWemuNssQ5XPoxguPlGw4dMfCf6MdRFRgPzOQC8Dwzbm4VAnqrpiVnePxcBJVDxZx
VJwe330xMAMPLjn40Gn/oHE2+gFHwVwYvCUj1Nvc19BDCp9pPk4ii0ACidT7N3i2yKqzbsBd0wrG
KOH4ScCE+fEWX8a+nfIL4Vse7DnFx1y031sByOeLzTBG8ZQc+HQmaj9iQoRbBgRS7hCtK3oJ1Y5C
K3wTA1bdMlnQr8gcqMc9xnm1A4Op/onQjUyavjaOv62npqsSN+i9VNQ5aOIlVSPfJyoWuYlJSMS2
u9VV28l10sJgQqaVopSQ9uoEQMTn9z3w/gcKmVjyN5Gl/M+b9U0mlQasY/zXhCjhz6InrFqp9DT2
+J6wl5OO0atOXvNxnHjVXsQxrlsPP+E0AgjOWjRxrOgDs9+8D1mYIwUQP6SykauRGAVzIu+Sdlo3
MHzcJSoDoJMuPH0fhVn4/ApejiTvq9YRGRfpnvugRUP5QaXtdWmGRnxQSO39jD1mMlSm0KGOtYxU
mFbgFMrLpuhnwhKvx72i0PF7lcna+EYlr/I8SX+tuqQZObg0NO6O/FNIn7eyndpjjYiVdkZ4zmdX
7XXD/ZO4yL1PgxLP6xllM1wcrvcgeyInEQbPMUgIsU5KigXXjcUE+0nt9maG3QlyJoC5CR1SdKQF
uylXO7TBynTS4s5fc1A7m3pzVZ9IZ9DilpIn9QyU2myvHB7We8tgzrLPu8ahOGytzPVK0l72Q8MO
yEMon6fTHkTD7+qMC70b+NePb3HPPZR1cpAcHTqwzNJ1JUafsWlH9wmuNVJzw8VP0JjaqjXbq2jl
rifLTeBZEb3/kwHAIutflM/3p8/B6kkaET8uqVBaDe1t4p0hq/w4vKUtSwE+Rc27L+bixO/t46wH
DDrhU7X7WBVfy9W6z8Qsx7u22BkAs9a7WPaFeH5mjb3vQQWrGdIS4D97DnV11FnnLHN2xlYCmNY8
KhcyLnEMZaHtC8URDC96nSWmIwHWoxYxRBaFnqjv5YqrAfTZAvgcaFDqe6Xu85tGVko6CoBmFV4o
mPbWF9Nch8S1kOT+ZEwJPgFtQ3iT0+cCwYNOmzfQHZgXzLZdk64VLzBuyBno+2trGZH6cbYwOrco
4kGJot2LkQsf3DNpusvMRbjCJzossDRLZyydkoC0eIlTwh7DkUoJupPlONzOKn4XVyyt3NcIbiqu
V04K4/4nra1jJRgKcyHk6ITuAn5q08n5I9pXQYYmTxzgl2vW0JwmACJ+i4gcBaubPQboK+RmStbO
dh8k8ZgLKB4V0F0358utWJsdRu9fOLio2HFqBKBi8Rbl4mqbwVUrdKR7W/baY3h7HabcctBz3zJc
5WrXk+WWvtiVPDDv11f32EZF5wr3OFLOTbakZXEr42mLO8yqFauEzuDwnLzu4dCs/1qI4OlJ0+Nk
QFe3S2QKRnicijZXVUsW8R8sCC6kcgQD49jTDWdFHx5xTHNZxcZW8CIqFPx2wRL+euM3xLe2dUYa
fUFhMQEOAdmxNxVyrYQgC+9mOj3PEYJKcTfer1P5QJiM101by+7TPOofDFB4YNAMaqGSlYHOhXaO
U1UpRDsXiYUXqDwf318WJT6Q2Vy2bgXRSmyVxM2tJgVS+WDElNh3HINhqASNApEP4dAwpaTZs4YC
DoP1D8Of4G+U3cJCKSZzRzeAxUm5gYPXeL7Devon+fHr6kS34BCrxTH0PuV7SBs8OqG3iPO1mXbk
BwN5KKxGqGUa1OXzZkij8RcNesJi45p6G9yPbbXyB5o8lfS9D5bSuE+e8WYka9Av9tAQjjysUNin
XEz6XjrRs+TJhll7N1G5bOFu9HjQw1n053FEKOwsBsPDmpVMwbrAKBQQvB2wFx8QLkvNBJY4AHyR
86fwVmVbp53xfrHLhZseGVYHj4rWzh6Qr6f1bOzDsWmKq9m4KIhcyhyv546+jrF5LOmMV+u1uc7i
SkekUX2GFRv9FEMQxW4uH4qUJ6Dqpv3AgCnptTdfWAxQYYkUm2fZI0g2rjfeRH4NzLmfdTnqhQV2
ymlqmZdMa9jcWlA044Kbat9zwrJoXYpuASZytpkOKVDUyCt0tTQe/lrAD8zpjiJI8NihY3RasEct
fIFBj4Lb1X41gG9u6VO90dTBXfrT9HbRiuIdsg+PELzWx49MmYURzLesYkmw46yAt3nVj9MUSOqA
DrxxEhek1qTKdslphutb0+IgEHaQNV9xIX7CUGsd4iZykQjnw8DtQgjU8Oztyml1zfbPi9zEjWOM
hgqGJNtZV4OtXGRNUhqtoNxx/quuXIIHLwnZBZ74PjsUD3N+D2x9eRScdXpEW1d5MnUx16QsLQ9u
b+u53QFH+5s1+8jRVtBfOpLsbEVVFp3tstNZSlvDjCayvAVmn7+K91PHQw13IMguG8DWTnIRgreC
bHD64/4JY2duEf0FypsOyoEDXZBnCVamrofGV2CzmBMtrBLSs94ozx0GOCHv9P6Gl+hca8CaGzRa
f5yG1iGd3No0VOjpYAM/9sPPwlkbJrZwITR5Bn8jNpsJEW7a8FwuSs0dt+4XpEJtt2BrZsbWs53g
oY4SngqkJvM1+Ya/xmIgf9pzTZL+4pZfBlGhsgf1LGozsPG9QZI2H8PWTODOQnu0og7uuuEs9vqt
P5O3q8PcPZ2b704PuhVc8GtMef8fQZYnzPu8VWyVwyqjLLSM6ChUQx4znUAZffOxqXM2xTc/baNV
SEmWsL7gsQJLBvA+7dwZicuS4O8DzhQ8dn7XzA1T2nMPCFhdu8h/SxwjIH1fYXRiIaD/572QGlvc
wC8LXpytiqJ78PvzqhNFtZxLVUETW+jeB8lWBS0/mhnToP6aJIadao8DYXQXwrffhaUeGqrtTPM3
SdJ+1bL0HBy+SnQgc3KoUn1yL32nXhcY3M6eKvX6QeZibzo2Gu6dPYy6DFmHs2HeQsb/vwFaYa4x
Xj4JX+0Kueq4N3BiUB6R7ngh1/o2tg+KdYPmK96sCIaOzXIKSDMhT/4Y7IILGuRF9Fx0Nyqfd/ny
uaRl+YIaVvbgLklaOUqESdQ2p8n21erWoaMDOAfRAWPSprLlCYyrsd2Up9XI+YsIA1oSNI0AJgX+
lfIwPU32ZjeuNcB5+1P7qi2VsVluAzgfrW3WNmu5ciI2kIw5EyIF4ARYrzUPfdFhTgU9jkcC9xR7
1Td1xzKQ7oqNbAuB4bmSAB0W9LHu5l7Gsw+ixhP997PllOKBPZKx3h1BZonr7SsDXiv77G99d97G
u4lLyZQqyzvVu7k7GCf9Hlw7e0tQNfBaaqIFr9VbS3Wj/opviAP+5xq4NtFEFKQqBEMWI1Wl81do
x4spJ0LekzILu4JL+8WNgXTCJDSnBB61KfZm5GOie6Ks6IXSKUbof0uAw1QIjoyG3fbylE/WSZhC
oH3mcRKDNWWxHumM245A0jVK6Se2UlGp4XLwcQp+Q9TvCv43ytLA6YjoTxUwTpyZ7Xu8XHRC8xYb
bvFPI5+D1lWwSv9vgvK4J8dR+VPxHli6cOvM3x3jzTqYLIJQms5ot9nqcBWSoPIDEEmQid/GS1vc
8/fZS75FOoqclWlA5sH8OjmdzJB/Tg1OlZPN+BluMTjDdezX6CRnZa3zAij+urOjUAm16vYJPa2F
auCIBSrMl3DLxJM38fFGj12EzHUgfW2mQLu3Pat0hYtXPBBQYpCjA1nTIam/wi7kGrGTRsHSn3B5
Ts96q/Ug33BdaB+Y+0CSFQrhazMKW+BO8HTcGnHUcxve/6ajAFXqgDZ32suIuuPjzRTX/12SrjXQ
fQbCArCwk+b6pHSTso6jThZWb2onDj1TkUQMVN8Fy1MysizB0eHxoGrRiZZkjFhvI8g9iJwDLlJh
68qc/OvBC0Re4AUIDm+89/dx1kcXt27qsOUhTYEK3GDgk+XI/dNld+roPenNmOgj6YY23vxMw7i2
JbI6LJFy4rHSpMxzea5XeoSSJewAoMlwv4uZ10jNK1hTmsadAoMMr+/89qRUeoChkREc4L5MYYQ6
WxtDqrIXA2vlxjgvODazwKgV+1vqyaTAjOWWuxFdcKxD+A5rHOI8pUDJu3FCLimQP5+60LugHaZd
IAllgGtEBIfEODY3MQ6aI1WAwxKd7j8KDUJfXOrTwp8F5EEV9NFoI7jr/ad7Entbl8FZwBtuvoOy
GZKrrjmYCt+JNy0Yv9AU2NbC+Jpp2Vu5zkScHzPqNEELvPBPt+qgD7GXfQ4bx70slrMNVVlLMnB2
w4R3LGh2nPDwu/92sGs/6Alq/ZXY8Qr5wmETDPdq8pwNTtmQYfKxei0WPerNRs6crHw/A8bOqzD7
dypgrBYdNbgZDg4tAP7XKynbQV3VvRWqzloDCmQqWgcW59DoCPwlSZpCEvbrNj5CVOZ8G1zLvrT1
tySMpU3uOekFzlRZ+C+ubiPU6pvQIrG/gg1HWl45//npUsHkRQ94+KWAbKBrdlC0UIy5wOZZPZSL
gy4KWBjeKS7KBhSXH5bLmjzwX8JIkrJ46WLYZv/Kxt9V3Ur5NP8rjQjGWLVSGN7CfRJDy9EivxYB
7Q+36HG3I/oNjlWqP8ojjwl6H5CxjgePLBp30nEVTWZyP87km8dbe1swQLe2W6hm/6p8ANzxgsM2
5B2sNaDzmrwgREUqYh2rDL+LXtjslch9TWOGmzHDcB0nxOJtSo+7VMWQQOyYUc1R4XSrckMpcBSL
d9ZfFQlTcwxm5N8L3AMQ0WFD92wd9RrwVPdk9X5QzzZlIYJe9YqbenhxKbKt8lNAKo7C9MInW+Vf
rPfPKsDRcVSOXvHOLwhl3PFHp85LIuo+fOf9t1Npu+XarvQfm3NkButVA3zB6br9DZZ1P3qx8x/k
eT1x6XBbN5u0D0oQWgwqb9zddUwDHLKlAalOrLj3TqAzI1eETURDmFBX/UpuNyLrPgVceiHSQGCB
zDqM/TFsr3nxMMgpoUX/IKufxCfVjeLbAoXnV2vNp1RjmneBIMk/0JAExqtStXeuscQlVwoe71rK
wCrd9PlV6PsHCdUnqDtIpdTKqZMgGPoyx/7skk9gytxFFRCfv0Htc0gA8HLHHoXzxtgZS3Oj3mBL
wYZSZwHA8r11kCwwWZ5+WiO0eebsDFVpEymr4EQ/G8VcYC/LM07ieZ4FHGmExuLI0beSqP9P2tlB
B65H+ZKLsNSpzLDXLbQaaUZPdfR4nM/5Ji8vJEtxE8xBxzQ1lNEkL2++PVAhhge8A2ODe5SkqfxA
bJyYpEM6EckRVUbO3k3yMka/S3QXk5yoGaad1uYBWBQrE2beoyGp1CP4ZA978EqaOyZMDV7eyk4B
pOHN5mjGyQ4GvOqXVf/klSs5kNn14ye2ttJqsRofi0qhBHLzhmmompyzxdMvSSuUSwKLjI12jcu3
LcoJs8QC6bPIV3Lxy4Y4tphHLh1dyOwU2M2yhKaMzirkmbJMBfCX2nJCEGM/WhsNxt3x94Bgnrwr
ksWTchAyaILfuYBGJk0VXppdoXtbKdE9Tz5Oc5+2UOxJPYeG3ZPXRYWp0jwXXaZsJpHrAnf4m174
mmP2LI1hGeOLG+hsIT2QTjQmlx5nYX8C1uUijEuQwLmk8fgv6VHQWusb8tv/iAbnoGsjr5Km0r7s
A58rimI5mjfa3FisMWrgOxmzPHpRkpOXTAMaRlGdkG7eoauJK4SALXCb4IaY6ggzQABhKlq5+jCv
q+j89nCPpld6pSdi0T+rReqmAa4mODtH1Pn3gcAAqLjpw1ztkMlLpqdMG06KRQkjz8J2vob7TAQO
wIcZMQgj3u7TMLDe7iURQBWjM4GcC94lXR0ZeLfkNSIymdQcbV++CvStPE+2rt4zHU+KvktrollW
NKwqvx+ElHi2P30hfmiC2SGOQNSqMTUVmCNHXePMQWbUfhL/nBd1tmUv4Xv9OEdAQDiGdIVdf92R
L1lWxIoMdeA3/M/iuQfcre6XyHUUZzr1G9qvRvESLKJnx5wpyEcm4y3jauecaQvNNKJgGGe7ao42
0vx0egfUdMBJM8LB2284UbOET/SjTAAXBAvO56uCbXvBfEiX1u8FbW2dIePnkWopwgTELQ9Ytzb9
Fbku4clm314RHxjmzr6xv97RgC5NpD327pqEEGJd0Ag1lHj9QRMdizHevnrJHtz446OLUWZvrNP/
BR+V65EDF6TrOHWTwxgvZDFAqzh3bJ8dabbpZC9u4edoGzYFswjaTVNm8eZp8JsJfFT47bNQmTy+
arHHHY6Xyg8A9UvQZdUy3YqlRyLKH2XMHeecbgViRTssZFy20d6o9FGpgQS1RgXqISf5r5Bj3eJR
5Kjymre7zIPmLV64NtD2wjSGZBOeeyoo2VU1bVAS5KESj+6t73irWQ+Y9inXZbHhwsdecVu03EmG
gdqwnQGHtVvZvWtI0cehkfS3R50WRtt8AeRtM0lQetu+4M756YQ6mFdKOqyvJjKvRwzCcXd2voKL
ewKzjz5LFLkZquaGKed/vp9iCkXFWI86T0KelatMaUvbIq7zSnVrzC3GJKCXV06hKXMTEj5z+m6p
d1K4Ga2ymEoh/tx2dPodKodVUsxfZqPS+wdVC9cyuBYgALeFYjToNoHqu/5htDizO5gSfXuRWCWa
E55MUYSfJb7SO6YwhJgWUxI0+enZcdRodTiNskFMJfV4TF1HzfiIMB7yIP5TH0sHfi5fq9oom+Ti
rh/dfqHWijxiBaEkLZsUDQTUBtJahYX0qKjH22WlEP6qxy1HzKYGUvyiOAbLlrVjT+6cBvJH2QYW
k1gK/l+I9tKTQwnMEtQxbQSHbCWKaTwAMenesURigxMhiALnoWLSQeOIEYNnLHbNZXTWCE0QeDBd
YT/mL9aZlcXusMgrY5tiskloaQbKaMTUY4NJMdZQfLsFVE9Mbq0+p6L/jNlk7Z8DxnX4rC6XTfSq
KtSS2BuoPe6Y8XKJ+ho6AatzJT/knFpHYzQ9a/dRv7Jgm6YGHNYCO053bgw0l57LT0OL8/l/Dc49
bMeinIkqSLQFR64g/wUSxRwD06ajC5NibMzEeB7Aq71saa5KOB/GkrI+/dWcJnOzInfcDKUb/O85
XFFDi6HoWY92Lv2ugFKinZNUrjezGPUHZrT6gmUsCWgTVGMFJra0YbiptThcLIol0QggaP/ihmSu
rhYvnMN8tztY0etkhuD6qeJOOduq5vmBIPRPCyWenW6J6VxUsAyECMeXe9l+jqw+8uOB8YpIYskw
AmJJZkLVkzX5hr5r5OmccntjUDa+4+1jv6QTUFg4KwUlrh6iVZZzqmt+EpLT+UWZb8JEx8sJ73Gw
dPKwdTUeaIVDCmAdc8lwC3JXzsCemeFrJX4R+swI0eDWw2mXaOsGfIRoV8WXy2bET3v4YVvjvdDx
pmRLrpjjjmX38WIqhKUH89Tl9oMBcpHsvNPTFUeGI8qoDES8cXtZJV3rC1aacfg5D1EnJMJi/Pcc
RELTWidquA+tX2CFlcDCfZs/d5+VgUkoeo94iFaHZibqubIV2yUY0tUnv7p4bHVZhKVAKtGOVzQw
9ADjITfa0ernazSnrY6Yrdo8LrLM2ZSBx5EQurVbRo3Sn84yIIFOL5NPhCk0IBT9wRI/ib0GVLaZ
h+rasnh+xa3ErmZc9eYDZSuGEfoAswouDQamV6IRu6tayYI8DFE3Agoorf9t2cm2w24cMG3OZN5T
cDRU8e0RgoE2K8gqovNlb2mq2PUtlFnQ9tHpqxeezJofjJkmfreAIV/ugGvoWDjTzY2mg7LkYmdo
Aw+Ho7/1Bh0rm7KV5jYLOroP18DaWSEJ3n6Vcd9Hh13DKZXcMuotayKxlEB60JT3iwjWBI+VVZ08
tDdTzhRiBNflSG2ADVdwcC7EP4Ee/R2wOqhr7IjwQ65cvV7a9WhUAO6G5Mb417+zP0VnpAh4oisT
4Tls76ae4kGlYZ/bi8yzPZpQ1Sx4y+rX9Uwyf2SnPjqWIErvzrhZ26EF1z0QknMyPB8kgufTlqUl
N3rldvtPMKf4WPeRa6eJCicvbMTfS+/gVObEoJGcQ3/Elgu5CLU9cLED74CDZ8dTH1c/rpSkE0zS
8j8bqjhdVdg1AWl2yWZqjiMugMSTJKkKE/3t8k2dy0AtTC3B5W/KPy0a/kpA9ijV+C0JtRCcaYdD
t53OuSvzQRc+7sh5W3o33ZCrhU8HyhbO0LAAfBMh9aspmLUCHsdDRnbZn+ZmXIwAf+kGvOgXKSqx
eYNd8JHo7W/A5pirNV28AxJUanmjrz1buw18re5CJzoPCerksiyplPyLg6fFM8QiF4W+2XqixXUH
7sR26C2IIT4gf1ea5moI1POKCZ7lIjtitXvSDC1uEHmkoFmNPcFkl8gU58YIqeLSkHbgYtauTst5
iz+kqA9vfyhaX6JnKhVsEp4IkmPgUyUXr0DYglS79/FILXVjJDrmruQAE/1WTiHmYXsp04L4Qn9r
ipTc0NifOPSlmLulEiqmxqQKtBFt9NFPtqqvTWtR8jI3H68oLfFRGTasCxQm+lZHpRayWcxRslLc
THx8YFWcaD71QdqIR6exV3CyGutFUFe+Z0YGTRM6IAhI9E+lhBVayDf091ORFIDfb0aBl3JBmUDa
ocSi36AfAlownwt+be3kLscL5HLJZjndl7tiuBJlIROAK11dfUneXr+B86upI5DyjzHLXJ1kLKEo
hIsF3HHHwNonvDBDdfACa73tJnB4gtwkjZijxxs5rbQG1g/ipSoufNpaq1hS1v0DvRX3hU2xNzBN
/ZPL2QON4F7ISC3nPDSqogW61BL6Hw11FOE7n7D4pDUZSsHwOiRSk4iSirrwEbRKhkKI+XEMchB1
ynYP5nJCO7osfXUWLW4COSQAHV/pNqsoEDlpOzae0/yA8TL/gBxdfjw/onmxezMSmslmpkCaPNl5
gJ3hVFIj4Ve1FL3her0nrd6wgMujiPYlExUb+Y6+2ACn+EaID+kSnXyfw/ZanTzGB5fRFAROdfAh
xaaXD/DHXgT/sxDv52tYB6T+AoqAmmqmfwLn6J+YhzwGcLgRCAPNP3a7ojFKEyGB/vpgAywZqYJ6
zIbwt9yIQ5IhKikoYXDSQOhAd5ahZi4XbT2HprnwcjhRU7Fn3mJLuW4u0R7rAjXArFSXB9TYRy/3
ozdpghHAzKZvFVVUP/PwrLTYqQ48nZyDv5XIXiZXZuFS9dYk4ky6r+1XxX3p7KGYpVUTT+qZhDUq
N+DETtJMW+JxWLEsloENKXUlz9ERabH7nL2G5tMhvB1HlFNu2y+Qn3SpCKHGJs88hAI3sJeR+Dq8
8WU8QFKvfPjzcFYew5qHMQYl+U8RNWhXERQfLhwM2nuR7DTl+VVuTRLr91UprEmSKkdIno1NyQul
1ftnHv8FEg4tSoizIWRzckK+uBe2FjJfGj4wG743LxY7LBMRroHe/msjrwVs4go0hKPG8zG0P8gn
pH/9m0tmPQc9XV8GlX445Jfn/7wVnuaibQ8nqqJ1X01QwjT3JYkf7BY9QE9v+TLUvFikJ7zecDib
R9Nuq+2PsxvMPCwGgPPnsaDLZe916/HbET+Qejohu8BWZwSeDsNNDWNN/7LpaUu5K+mr3/kHG0bI
VhuVflwk13z15JjIdUB11vFftXQDZTL/7E7ZhHWCsnAbTqYnBju/NrjRItnu0qpVka+QiqOnhakV
RsO2Zce93ol9HrLV22HZZD+sRBp8ynWhqU7I+r3zu4d+GQvu7d7bBPUHJH/yrnse+EtmXQ6DXGRe
GLV/xGrmGilvpwlsC1vpJOsb1LH66FoH21AfCCdKW9RfO+DF4BjZU6TGRVD1CCCXc/hyBIFYwC2V
VC4OLeXBJt8y+plNwVBILqlCZoVOafQQZncUz5YepFWxZ239N6Xw0m3Dwed4TzHrWGY4MMXdUMQq
2Of75O7Lb89G2Xs6VinVahzjhn8QvJ9Yu0xVnbh2J3eQbmCj3kZVyuVj5Z+QtvLoREy2JuCGyvv+
JBrYgm3WX/iJpEzaQI8/3kqSDEWgHxZN+m9fRdQANLTmXH88nQYJsp9Ct/sntPSAGIHF/ZEwCVgy
ySEl6GlgweNrM0OzaAFQKHDXe0SG4sm63oqpOgvOKWZgLiSSgXlvzj86keraG7Xly4lhxXraLxya
0VkxuqUdgQrSVcg/ID3OvisEOEg2oymvR4ccnUviPPKGKEVYKkl27UfVHfQXLmpIiK/Com5+vJ34
FzjLozyy0zgJgYouZL/XRtK0+Q0fUSKjVk9o/RIaRdWrAf5cWub3wWReBhqz3Asm0HKgFURTYb2Y
54fpQ0AT8pOsG2tv/hHSVNy+0EDfJaq77Pq58XfGv6giSecfV+eYXKixsZgjdVdUvIEVjcX58Sdq
KIl5i1zu/v16phwKFjyPuEe4f1YGzP7L/6Mf4v0JKoO3ol+s/lv7ucAaqvSXK0MZ9OdyoLFdLXrU
SzCmwC5m86+mYeGTPL996hqdalhoPtGbw+ieJdSwjM7V5uU3BEZhFNVI/+CIdPzXZz0ztMg7/SdP
P2/Q27GNE26it0VfDbMSxY/nL3UtMKZ0ESGUFD/aCDq+qVDv5MD23e+G6ZHOzxZoL+3gQSNnCsPq
dMLLGxT8o7bsKBhFNv0nadkD2u9RM2lUOHO9IqHHhRkuy5u2xZe7qsjx0r0yHRjn8xBzYtAa4l17
FOXHg62tQx8T91PRS6N+v2yPo7sl5Ea6nol7qF+F4MtLO8h83jo8dfb2RKYRP7PZqfdnvy9oxaRQ
9DU5MsGT+D+D7npw2ZY/UsY/hs6CcOUjp0GipqRNMZkcR2qQxXWBGEg/FeCPxkZOc/wOwA2EbQGZ
6l4EZ9h9umKwKW8l6r+MZuagU2f5xDQozxjEe9i3GOhSYhCUvN1G2zgbdx9dLt/BrlTQlwX6iGbP
P7y5HU0VbxOxMdbBpBfetjOEUzGKV+yYBbB+kwYTW6WlDqSrl5o2CHrwlawhuHFvFLrvhvExa1Pu
8LoD0FutoqZ7GJ2uG+m4HIJgnNVVd2IuQKmBTWA2yYwBkyEX3GOWYXGLv9wGbW4LRuThL2CfKGBm
uSCGaCJ7ErsMofxKVwGXL/00hW00J1sqbr/8HgIAml56AScsDiYrIE/UwUdd5jHWndl5dyMNUnZ5
vn0BLkubRZ2FwwNJ9KKewM/Xii3lTpqKLg72ZlBhvoFJnsDbnV753FJIZghnFm9wW03fovW0vyt5
phopKcpCmin9MNRr5S4n/vwnFDi7GhfrPMWxrwDnpVYXZJT/5fz0NctvwYooTbJZp/Jn1kKQk2Yv
LX146Ow/0pnxq6xWSqj3vXYiTZnDrMr4oSwjbw7yn9vtm+OElQkH2N+XdzJB2yFy4pkPyWTLdsT+
iyvSRoXoVmaYYUBWodvv1uqccQSlQ6xmc3bjP4ExrMiOZD5RQ+v2YxMRDSsrAcGaS0vMDYN3gPH3
EV0hp2MD5hocVblxADOVbUAK3eCL9Su4FbzoQa9oyDRddyJzNy29sVXS/gwEMnlkN2wP1KEI85pH
pWF+g6bNOXI+wPI+ys864PalgRGkAZTnO86HgfysxkETtE1qV0AHFyG5h94rGYgBgHBqoBu1Bepx
JD6xRY3MlMe2kwxTw/8WAvIk73LJXl8yWzO8XSAPlODOTvhe3KaWW0PniEKBWjNiKsJYWi8ZwARF
2CX1T2mlqQB/VAOTqkB9sswIV7kEoUI67SCtzEnhBvv+dajTHWsmwxIVbcfAowUZwOpTHNgck39s
q2rsF1OGWKi1dsm5iviMu1MB+/k1+Y1AOGbyfAUE4wC1jSXoPJd3FP16tf4FajNg9TffSZlcGJ3A
tkHkxB+1lUtpKMSCfu6EADVP5KUoqzBqBClohKykHiddU5zrnP8xZnCIKVXlwSWIk6No+hd+NmYB
YxwmJD0AAym+kxcmPzRUz9vyf/LlqWo31aGz6bIIep/d7xLoCXxf3vco3C6/uqJWXqYht1uGGa0t
JyrDvJkwwr8+iWCQRvFj6dqO4DRP61EEQoXEUOnFZyLVb4wT3hOg7yiVZ+8bqpPuwA4Lt0WRWPJL
h3BWi4bXORcLaDj5jO23xyO0+zCcsg4Z1OmhlehJ50IPn8OyG35Ctn1//ln8uf+IPZvds2zNM7pO
zh9xfXNSLDiVuMzmnvQxe3ZD1971keGdfF+NoLJahrK0+lTqq3U3LAQcJxVMnORbzYEoJh2bEz9I
Z5LYR2IcvXdaZFjunubvMIrAxQLIFOiCUJpezS/PMIsrDRdT64dUoozADHa6a212SuZjySgwW8oc
RBWsjTyhdDqxIOIGxPtYs0Ggo0piy5KR7Q3gs+95QbPY5kZLdlkWYor0P82XzyTQ5Gd96DDYGCN1
K5Tzj4g9MJeRb7aiPgL9MTTVUAT0ZYfoPLYyz5snhLHQks4o1HIWhZGs3QP2ZBiAa6Z+VJFdvgQw
mLKVM4AGPd7JrPhh6hEiZpBuwoqX7ptiRcHhXy0m+6ggTfvpxEpLlKehDE/9FKF3BRjZwR2eSKsE
+UuVb2ptQDildkUfYlvolUjA31R3IbMIg7tsYGGahML76DCSkJQWViD2EXfbBZWMBI9gJmOrG9GN
dx6g5GmqUDG3a5Jt9klUremDpiQuQ3kvuGVL2AFO+1xfd0reXfWWiwZep2DjKZLJo1a7ma36MP7s
ITq5lcCHcRMAbXOXFQqIkGLANsOLrybKwmw+lAnIJpEzhGu8S+d8AZAncyKwxHR7at4SwJ0Mt1oj
hJm9ij2pu8jA9Vm4iKsG6k91XLgl2cVHYX/uqhmGitYmodrp9ingwEsJ9CfuPw3N2VArdwB+u+HM
nlYe/cbmA4zTysWS7qOiJziUj5PGzHrvgIGcKjXfbr/Q5wrAm6NWJvEFNMWjPLTiePGBCSZOZxlS
No6vbp5PqFlGq3mzJ/DTFJGb+0sJFn929X3OJR3ZeD57bFK5Wp3IjaVeBb5sqFRShWoVI0vNIK0m
t9h+fSlElGeSt2jfho5MyObXkLCaXhkGNg8wDejDo+1iPGtSScuuNEfVz2WhG43rwWw03+nPBmkb
oC2VcA4wLJM+Axg+N5KMZFpLFhD/C5GI1xsNlxOteifGMFqOhDIVDljE9DNCyEz0hNmGzl8++o+a
smslA/Ug5RjMEcTJxnFsk3uKVdKP7cIITdJ4fi8RJHKDXjUf22hbz/cIvsQYITdj+1O6mPt0DXwI
3zNlrxUUm/XnpmYkfSK5zdVFdufndY6H4Fkr1fW9Imuc5zlHTU2yVj/mY+3wxSscvWA5GHfW3UfN
SfKoJ5H6gWEdae4/mEMpukwY4OMCYzLEzTxkcyw/Mza9mDJR2hrh1N8G04HsCkbPl3eFkLxdPZrt
irpS9ru9Id5vB/J+i6ecDyTNG4mTa5dJ7drC8jH1TE4Hez57luV+3GDsSj/3tDaR0I5vfYqA8+00
W2UgxDR/Dil3oES0W7x2eCBQg/1Dn88HOcLmPXreh2v/3CtBeuWULw5dPueap+4zmKzVBcWCBQI1
ZPJl860WXjzbMN2XaL5fWAHXYF5EVnYz/qnkKBDaGe+HHNBkFfT2mnOSXPgqjuRNZj8t/8g499Zx
8zHmhKah7kcec7AEOBA1ZXN0182iX418gxRaHp8GCa2p7aB5yZTt2rpCwJRlmrfaQtqidUvLB8YN
iuuspOq6C0iafbHUmpyse36DgoL8nkg/01PN8QjuO/icUD8WU9B+asTV2YkkkEyWYxtYWGQ49rpP
kfpPg0QHN19TrZl4ALISjMKHU2mqwYhcrhw98a8mOktUk4DVEWRtvQiilzJZXm0Y0cbNWWpfojBT
eB+ZcfboCogTKKMNhHE2jYTD5CGob0lXt85MBAOFGV3a3CSplD8gRKmGBxUxJnmCsWMbQDRCB/hO
u1aSip8mJ1UKPAjMCdADnUMHotLkwVFSHXqnzIn9L4tsyDImyr2eXwyJxHDnLT4HRaCdBaDaprJL
gzOUBdevTBvYXuSFQYN8l30uW5NF0CLern2IOzoFgq5UllfMvx5q0blCqpFjLtLsjcGwSNXCWLGm
TKW4LKjyXnM73uzx6gY+83VJR75o5AX8CJhFjbg95vu5Ks9mAo91Z2kV9LYt6w0awEXutcKC5Yq8
D/0lQNY9VkHmT7geSqkZNj1Hu8VXCDi7DlMSpxAXqzFD1lX36D5Glict3mbB2fYSKcEdy0Gy0LPc
fXmxxWsJupQ8oXWFOSezJpUh4bll5Sn1u5o32tnTa29vs26zMtKmNIZD+JBI2hP0WbmAStUoBD3M
BZlTe5H6n9ijw4R0TL+8nu/dT1rwP6i3bCIK8su2cFo0wcDiZnDUtorBZ6R4MxHEtEzCMzBhxWnT
TPz6jfFu7Hf4gVLpIHRlFFW/kp0fnh5Lq2RmZOqX2ixv9zBalZ6DuskqKeUz9x75kQXxKgIoptEk
RDvEP2de5QJ85AWwRtx2ya36yPlfHOPCQXprPMtD9b9diA68Gh2AuW3ltEmTrGsQWAgYpWLsR6Tn
3id5vfGdKPzHK28fJWAiDS+MQL+7EcSOgPiDcf8YOE2cMP8/GltPtaK8VCAZZPdIt0ovLJAFKj80
MNOSJK2qvPX0f14DCSBbPjlQBdFNFfAlCneUYEqbMnJACLC1AZXdKHSs8OFgRlV/q+wcZqE2UW8m
G7lun2lRtTZqKexSLtIW2kR/IDoTlpm4ty/4gxjFCEqtEC239udHMnZ8yK/qZGGqcqEc70RVqG/v
1RC/ayq8lAW3nuUM3kRTH2zcJnxPbBnCm7EKglH23S66uGfNPT/pqLpsjPHt5nAYge4U0YXa55Vt
S3BASfaKyD9mD1WkN44tlU6mvE9LwWuk3vNxnwuu6Rho178v0nmHpzeJpRnns1/1mBMADB3kCJjj
fNdClvNei0GsouSbYfVXYMf7MLZgi4Z5twh/5s50hhiVOlfUT+v3yqFIOOSsjNDFplJ2rmJQrHfM
UGm9SHpL4wkG3F4DYoUStiLQTr2sX9oHNEB958BwJ2sFG/EIFEL6XjQbwsGvWpHIOkiyJAdpuJ2z
agKt9Jx6lY1mVz0OqtEMc4QYfL6sRlZl2saZwB/lnIYcc1wkzpFuuxMtQpyt1z56nkeGfPmPyDZ1
js6TtOtkWm6LRxUTigDQ97hQ8trJb/Fal3BnJZ+S1jYwezTPRMlZI6kBQe9fdw6ro/nyjDRAblE8
BpoBp47iXyqXw880k4rA5XtmAPNrDaAChAJQfXv69f5qS28NhHsM5xZiBdFqfOpvryJXD1118qXj
wmcMu/MWPhYkqU3vFIioE89Akz1O/59iy92FQdGFMf9k9W+lkWMNE8YEHrDaT+TzgiWeOqBold4Q
cl1ntexFwtVXgIcfc1KwKzf0CmhrOxfzjEKssQiy56igmebqEdn2A/FN+d1WvLMxxVDYPzsITid2
7C7ILYe7C8J9IUUj7X3JFL9CJClS5NHgxAF+6ndcr9yX2GZVSwIZWzrETGNRA6XGld1t6rG2kU4I
CiooVmPRI1VJQJ/IX3wnD8rY7U21Z8Sk50PYTX46hnBS5Lpy8MciKoq6FI3ohaUDxcvLm3aqCSU7
7ii8ij38Go41JrLv7VDroOpmciu2ucved7BfkZS05rPzlh5eayct7PaYeBWkqYwTtjnE+ezgr2RH
PFKdy7020TovW0RyoGhfubcP2sgaoDnMsCrw3VDdt2MGGu2I/Q/w8W3TzMdvNZfblfi5ruKH0IOl
/WQXAmWPEyuh8HJBRMglMzmmmENJr6g0jxgXODoKSt5IY81sJ5uI3EKFGsQ5wL7NbJHTD6Z+eTEH
fCXs6YBWcvbGvLdhuBsPN/8WMcbFwB9f8yzBqXXeqwKbmAxDC7zYSU6Ogf+135+mz0XbeFo+P4z6
qkQy7pTUuKGyKYISmp4RvlkTvd+Kh+Of3uOJ0fJUkPpzZv7pP+Ph1Yf8BOPzd5so57iUkQtC9sFd
cDvWbWswsAt0nbxjClEtg1OdCb2k0Y+Q6kEljdkPbVb2Uqvth4aP2dCQLHFUhN8wVhhy3l7jHUox
0li0c5MRsRtXwc7O9VYn7+dLaMN73I94KWBE8Sqohk2MHTgHtZrtBgVfGZ3MKOXjqpa30wxBjfzP
CDv34dGnR9QuF+0PAwd5fxx8ZgIMCLudMupyZTUblDTavHjrbXN6O0xrPFBfABbsuHht3RmuR8hp
8viDFiNll7O+DUvqN9Y6AKMYthnAvM/4Q8qJaOX4MBLProOkCEc2yVjJtyf5jIRxabNcsh82N7G5
Jv06QSp64lmQKCHJd+npV15jAOu1jri8MEM5N86ja8/Sns+G5RUCsr+5hfDyJY06A3nGzZNIE3Mw
h+P9wiYo2zFUREa54J9VRvlVSUvur+SFKtBVLDYyrnpE8vZN6piqR/z5Z24aw/NNZi3iVTJWcXbI
BLOwrEMU8+uvxuSlZSPpojNl6iOSMXjnYd2L/rGqZjs1dWRSI/60TiyMINbaWJsytlMpgdaSJsDw
oISa0EHH1m8l2BlQ3s11odqzbfQ15TQjHja4xl3zGC0JmaTJgt7/+qFwXfGKQrgQwjI33+15yyyE
9OTIQgpHFF7Q7CY7oLf+EtCniOdo9J4tMv7GLKw/wZ/Vd8xVzZ8WFuJd3jcjy8WGpr/ZS4+T1QNd
uBwlCpzEqtXG1JJveRyjcSRvubDgKlwTmgMew9fup6bZcXubBUZZgM8Hhk/AwSmm2y9ycrBqPWLs
DPfQ1MoKOIJs7OJOfxGK7yJOppsniXxS7bRWX2lI9q8eV0iJSfNTP3Bt0q6z44rLiEydPs53rHv7
AnG/y2htBPm72Z6SLBcHj0m2PIBO04uHsmbGGz83vxzETJ4qAvEFoLhLfSx9JGNxiWXOy/IPQs/M
qu049nqxdFXVLF3Z6MQ1kLydoF3gAqDgx/XHhvimNE8Mue3s3P+n5HKJWVitxL/gOQuh+pTN7SIg
5pgj+AjjT+CtUaDiojilNpcRjir6G5nyBOyWWCjZMrUXcXm8OHY3VyC8SI0u8rkd6GTL1bchaSdM
kxPf3SA44bwBcMH2Hh/hrQODK2iAo97ZjOAo6Hm1RMfXP5uc8/aIyMbjenRyFLv8VEVC7Hbyu2Oh
5RPyQpcWsgcyvuVPIwlL5C9inWtNtLr55rh57X0zDOsRpQLX7hwzJUV+XvBaH22kkA3XTMP2Vg6q
fBMuPax2gawGlH9PG7DkSGiIyKLGXBAD81cwtaCF4PLbg5IzPB4qx6av4srhaHQ7NOdBeqJcAroV
NCSm78rcKMZXq90Yg65ZO/Ks46yEm7PkxEPk20jLrnIDUa31QkIBGnCT3U7e0PX10QHgdSFFZMfJ
faqFSWTXwRoIlldotCorO8X3maBy/ld60tpvJX2vQBFfhgH1Q4Y/EeM8M3XXLXReddEuIteY8nnu
Ek+p8tdKZjtpG0G5SESK0Zpp7Z5rSbZN4O1BIbxXUg0YO2dBFfjodlzdh4OOSyfuEBGxjhH1vJXR
KsRLopFSRXagjLaygTjaDIovWzEoGrCHU9Vjjbf6dcZmk6nkS0pecTe1siYnVeBOAlLj5swSd+jm
5oA04hKO/CJZm5st1FMr6F0XnS9562skRXLPSr+8gvOu6PZeYLxbH/AbBgMh4tZ7yShICtUjG9pW
B8ghiOLwXSp7iiSmvHDgJhEHexHuawr6t8LGvummLJTCsJ7Fn2OXaKFzYRgmP2JVIxi+oTbh/m7R
PJKAj1TXJouCP4en3aWwdWvR52XHnFysqiVwYG2cQvERWAnZsKCkks/BwZiDb3XM0Ug8qP0dfWau
WOAZbVgKslbkmW8HgJTqMfMDTuRtds8w5lOJSPoteFU6sTk2O+W5tkbFe1ikg4f8ojqi9N6wm7ld
4rT8yw86nprmaGyU5BKv9eqhka75N4APaJPm0AUfH5QXLxoBCpt0jNqYz9K3OQyyLkplIU5Mrkzd
LVXc4PeyFLYS5UAeGy5A4AsgaheJhFBkIMHgLZykXnEBA3yRHnVmZDpZVgy+blf1lPxKRTmBdlK4
WpUzUmII5Hwe9xi/gCZ90ubgW+bAyNaCUJ3ciEhIhI6R4fuqN6mcEQbUqIM5DZ0w1pJnShWCCgvA
aOZEPZGxQkcGjTEToPz4h9R4SL2RFCj1yWydcFKejWQ8S/IZeIwd5iPWgu4AJHONCNZeA9WetSe0
ev6h/Bli+G+Qj9RtebYJBae4Rd3D1wXyWU6MY7HNz0CTFGa9oQjMA2xxdkikcrJSfr+dROg4DQm+
f5jDGi6ugbAKv8kTpNWU146/9puzrG+luB3qYIGFFg7Fl615CQGnWL7U9XK9Aq2Z0P1JsJyHWcTN
MhzhyKPY73TFuVl8PTnRqn9nLpNP37/mRshVePY4l7WpFGyqwPqrzfkBwT9S1V/dgP8UL2xaexQR
v8BHTlp7Z9eKJbssVGQ4+QdgyfeUIh9gfOiqRwOQzaFoHq4ymVWHgdFv2GMJoBO8foe2LT/NbACL
OS90gDoPx9TFMnFsTJy1M/p1AHtmSvFfiOJIXfVjM3GzLMwY8JQINuTYX+tnR1E932QEfuaCeiZm
aG7m/d5UQlFu81iiDmdh1+yKlN9MUcKzgh5mUA9h/hxSEwBdd2YLdYZuqMbFLJ0yvvPERqFlJ6Co
nHjybrdC3mBaKaFANvPS5VQs/SE32sEMwDQJtHRglnugkrYCPgu9n9pMtG5oCdvH9/xup4SyWw4o
dBuJpfZVXU3rO/YoS4wX0MuQfrRfIKwh7+iFgW9JBg9ZjMWnEiSivJTJR33Bcyg4CFJUqGHFnD/E
QXL3wA80SBZ4cunxhU2pROslECqOwTcBdyVC4mMMrE9y97c2jpFbVU6Xy2wwNSsXlwVny5GiPNWA
u+tN+xQLTHxYz4HEV9hDgEalu0xKclDjyhjdVjBbKZhNjVCYNkpmDAPD561WS4TMKFJqyCIRuVk+
bdiW8zW59CY1i/w6SvYvk/TCkguNhK5Z4dL2rIqzb9o/ZMpySfVplUCgHRlF2uPodrt3vMnrCc7n
PMVze07kdyfR1m+zqCxG5S1A1JqoH19PaPj+hSTCRRI+oMPb1Lzl4UfESnc3M4lTWJwMWaDVQ7hE
yMYNp8kKLb+eMCEceKa7vVWXb1y0de0B8nKIHsIbN74EIvAKVUEYgL5m1bMHdn/BOuB6BKSyTH+u
oq5n1iJJYh2vbLLbuRHJk28rtN8twjHtWUTq69GxmsZ+Cf2hR2Xk0PapnvCTYQOZVnmEXIDVbSdX
OphYQEFYN7MWiv61k/ZxTXmFGtOrtNhe/nzktcqRfDXaRNpkHSraifehJzw+Gbf/rA4E8B0h68w0
pq0K6XSjKY/IgYaXeaDAbuDt42Fx3poRUIJc4OkL6RXWdCxR3MyErjFHe+0QP14yTzBnbIt+Z4dL
jlWBjStmNwZ/EuoapKdomDLmExtF52Z3mmE+u5sYaZysA0MNaOMOCi11JB5KZdH8w+3pXvq2rJq2
S4QzKUN7/HhFywWzbV2Q7jxiUgXDailDhxTxOKzTyGBkE67mnsval+7M32LMh2ZdNHkwb54pWTw0
ZnyexrO13MF6fsKZSeRbSZi/1QfJjYz6DC8vpxF6/njH1DUAEMweFHsEvyGcf2gEstHX2PLmCgOS
EUClsM9xeyNj0n/G2g9C46DDjeUWEQb0cIkX+VffHiB7ZV9PxP0kXspYWvGZJHxxVSD4AZmfVRoa
FYaIgFmRQTl6hl2GrzlgERvMQtlGFF9J84yNcOQnk/DVERDv7ADmurn9lriujqYfJGbR5kUmSdEc
xJ2hC9nWcCeaZV0qRl681eL6FfP++tkIzvgPcjoXmRPxHqWk8ZtBds5FkFyRLCJDqDXjNXXvW4nT
7gZpkM9MDt1Cl24InL1uMVR8lJhhfM09FRdl2TtyDPffhnV17qz4bluAyaeXQhAtijO7vyjs8yKs
cs+r9RS2eeAAi/mggCqJW8dLHzTSndHuSzhF8JfjS0vc9Dte/NqyteJZucMvRw9nrn+zogMo2xio
R7XvyC+X16xyx6kelmcWfyL380PXXIUcPhIDznEDlxUxl1xA8b+81OXHrnisxgU+r3apFYWEPtOT
ZG39HzzyiBqTXzc2xY1jkQJMazaOxBTqsZG0nwyZYX1nffSr0hNjFTnEaY02aXory03wsZWUVWL2
wr/KwsGt0HKiYYuu6PMXfH6MA4gXfsPOSgs1F2/u8aUTp5bGaEriZ5MeAgkC2KXxGJ0q5tCXUmJm
qPDDlLhnbS4TnoMf1EnDkWQyYOaPPmLPF94hPAzVpXlaelNfUqcoyd/2gFoLDHa0SLSfUbSj9D7M
JEPWwYJvA/qsecekzPtpjmPNTEgF5wk+f9C72eh3KTZIBfiqm3DYp2wS0nFW1djo6e8e5D1IdEJd
EAdgZJnDRy3y2WBKn2UEwPjSBDEvhyBC0bCoWcPj+8xusNkmaaYFAPzuT7K+eeX3x4mi0lEK7BfO
v5fgwlvChljG6k26qb0FZ8DnqcRf75BqivKeBbkm4yv+vE56wB4wBfiRXMXBDl/pHzMA9tb8Ta2+
Ad0Bn0B1W1AtBBWcnkKYF3l4wujOnRF/ok4oMalTBXPPtjZYrnD2IzG6DUt4RlGX0kyQvcJeW81/
TXg+C661vGQu+6HwaoeN+IqzTvt5rx2GPhrbWPZE7IUmj7Nz+rtBSc7OFoXPs/A9IktvoeS1C8Cy
sdJ/21grO5fKHQoHgy5yAFhA4mtsqdTH3hzc2ZFosn42SUVwn0wIU27h9MACXAUHYNUDlI5LZYh1
4zxI7c+9zGL4rvhagzTlMim+UySretlY/rcF1DHayBBBbpuJ6CcnzZzuNsiFFBNu7c/Wdt/2CPoE
NMBFCO1jq4ceBZwPa+mpFU9GPwIeJtuh5WGDruA4zjD53Cf7A1k+WbGeqKjEK3DvHI5UXUbxNMlo
2yy7ohtpmN1/IZjqgVIdu3qFKHtImSVbkjACOvkgZEtOGG3/Te3u0YDdPLlE/DkAShgHiQX9ckBZ
gpjgHtDcMWI0I7BiT6C05aWKQ2835DCIfWuCpaLhsXyXf3SQUguTIC4QWGn2PZYwIZhq4upBWxM8
tF1JCI4ckuRJSgInGcd5yFCtNWGU/mnnulJZ4OKCJVAY3sz43kKD35xTW6HLxN+Pn3agowQCDioV
MhBnDoitr01WMN5nk2sTdMTbEfHkgct1+RwossDaFejtOei9Hy2BeW6ERtWnlrVbq8Kb+Jl+uNWl
KHLcLeGHKbtooQDkymMhho5Mr0NrfhbE29mf2b2OLXp2KrafV+rALIRnKWP8zg5dJDcne26aR7u8
1/KFB0s1WFKOfivp1z32enXbPaPcGt1aft7sy9aipayeYCtRbtvrorOfhFGP7dLY39uHbyKoGKVx
xGIf5vyJ+yzEkqI7VQIu5zNpyO35F2iRcU6kyLVH+oZBkcGJ09BzZc/MFf0HdHWAFSXcP6W+3lsY
7ksTqppXUfVFKNBJRjGhGYebN3Abl11HV45ZRMTuIpWSOiLlGbdidWbqhAw4kV/l1/1VRnXLbPhn
lvRzoWR9/A2U6ML1qpwOWRYjMA2vKiuGObijjvRyiYrKpj9SHgAI0K9VdTkh29Vo0XqD96BLGOuO
GLCslqe1elor2vIXfWzfU8PnMyptVbluo/jhowNDu+tJtkjYP3f6PdsCecA7k27geSvbmNVFsXpH
pxUTCETTrfN+s7A3BS9BdUlrznpdckNaiT7GwI10ixWCk5DDNrR8TKAXmByLG85SAJr3qHvixc/q
DXlP5nd09Zb+wEs7WhhR9E6CA9PTObGKOcA1M/O9hhB7x+vwE/5t55KZiLTumy+8hpFblBEBJ1jI
vZU7dHSXo091zpGznj+Len1Mlrr6MfIXrgLdkoZ4fcYpe9pl0nZV7K53VxW5WeQzuHpDcPPQiBYu
icD+uuQrgwvoyir3bOICQNPrmpk6/III2tBzsfJ8a48XEcXcIgNgeYcdL9A3m6JvCE284+Wa6sZ+
O0JnhDlWkR8Pt+3RGCs5x9rLF8xImIUdgIUvx2DRu9DMpr1u4CT2+BxSPy1q1E5nKsoGhggGAqEy
LIT8gkMFaTKUgV7+Btsp7NJjz1IATiN2YJ/2iiweCc0PdM5rl4xY2enfxRTzDyXdSbMXCRUnWmT8
aWhDIfku9j6NbpH8A9vkEedG07MeD29XBJuc11XQrclcDAjaGjwlwWPPX8XWgvCL/aqHiWSmp++u
Mr3w12daYV95gYCTxImWvHMCY432gkjBeU/MX+UL4K2vAKHPqnARRoivnHNhPmqW9eEDQWjy88fl
w3VseZjq0vay99QCY5/lQFIyRzznytpuwZSSgr/PAPUIxMyWefiPwc1tlQh9NryT8l+WrDQYVcln
2CL7rMY3B8JGhOLyiXwophDqOAEnhiJEHnP+m+GZjCWyqp9KFKhzJrjUkxJ6GqSP5j9lvvmNiX3N
wRzqPowrVOVBXBzW6MyhNLUyddhB2XB4xrG+RFFhVNpMxzLLr66CUupVIpRlvK6yNUc+gvmJECoD
jd+C7uMFcHS+94hrnz617tWDX1g0V2cxZhPLQPRmMCv9QQiGT7Tpi2UodzBX0AzcPQNrYLWKWbvu
Fugeg71OTgTN0CXCKKhgIT34fV4iZvP3iU448vQGXFBKUlNUTJuz5rt5xHsrAt5MBoBVgkrWAXWp
7it7B2+NtqScj0fRdxGuzgfXE8kiG0gZfbIDgAN4ZaWqmX65KB5AF8Qp9iTbGIAh+Sd/p1tUWD+j
BxPpCjFAww4oxfjfFgqP/FHgkic/4pr1pwgNEE/ZldRSeiMmm5agjjdn/bX+k7wyOEIUkT68VJ8X
BAc7PKEvRiSRHVcF+emk38wXqPV1NY6mEHt7lzzNAeSxkiMn01+8S2AWBx2VVKlnR2+FtsOECKFE
3tlHvHf+oyv+Wa7PEGVYx53dXrlW9U3Azq6QtxmO0pjK3nNKi+bdt3g/XaGrf8MAIFpyyDgCsoh1
aogEaCSEUs0QbUfA+7y3+X7uAmGpmZW80ig7YKDK1KpOGYsvQzoIcvchVfWFCkkqusZRWpnVR8n3
eNJn4quL6YaRo1ewR5x3EwjRYv4rEHVWx3y9YeofZ9tF/1slK6Nh+0wKJsX82iXakIcxZlcTay/G
6BnGRyn/X+r60xq4c+TGuTMYSBlVTZsjftfFg5c9Mw0TegD5lRgrEoOWllJQ1Q2f56KEIuDgGWPI
1e/faAG9r1zmYJIlFwOO1+TEXcfphDYo1QwA+V1+2ip4JM5dynF5v/9+de4qNKw76Bj5d5ExLIQp
OA6lUh3mxhtpOWI9xdVTIhacZzkHkrZGYMuru14T0mDaxAezXBq27eIq+J++VksE8/KEYj0nZHsy
shp/Tp3vhjZX4VcXVTPyN2HcwbEhsdCga1/+OefEqejgGo4kfsIYnGVSOr5R+biPhuFpw6PPUEXk
pKlUgBwa3IaexaJM/fSboF/gf6P7caMr7WmUwQ1J/1aRsZAZlsMlk4Ld2qFbyjxGcgKtrtf8/TZp
/oclH30UDW2nxS7mZCkH5ZRrHxuYMBKFof+Nnq9c/7YS/FphHjLbgFCCljcHR6K+zSNeagy6u6cL
Qwz30pgqWT8u1YjdtRTjdTP4LzWBUsaeOwol6bbgBGqp305mmYilYADMSFx94ogkRCLqWe2nRSyr
vXk28qWglTAtjUaNABfFnEGrcKhTNlRnvL4eRRkjoojFB64QNBh6QChZ9fGVG7NgSqBEhEN5SWmJ
UKzfJrdhCH8M0R2ZrGd+XbVjVdmkg9MNlffOii+Fr3fYURPsMx6ycFDXSkYWPjLzjYYDsi4MNjRA
rAklG7+NUMOhV9wAHCpBF2bqR9LYMCjhqkpNi/nOLwSPx31mDpL/1RSSt/dAyXfblmVnALe4l4eI
/me44d9id8kbI24ne2Iw7Uo2xwVIKIcgkw7wCg+Bk7V6gZAkiQk1T9wG3yVPngWth3UpSJYAHm3Z
BaMQ7A86Pj9dCXHYRAEir9DEmyJfMc4BbUfWM0j+AxfPvInkb1LXjpAcWTCvnSiHDnLYOEkCCvhz
I24f8womgJLeJs9kUvFut4wujYc+ps9381DlMuh1j/zjO3UkbUgAaZXbYpPDpfuS/p5qjL236v2n
mEHq3F0NSiO8P4vT6mEyOo3ub8J9zsM5fq6rVlhhuaHWYpzvn9OoQHr6yxikpXOhH+6Dk+FmdABj
tmHmpF+1Ib/HTa9OW+eaIxq4bUR4McSkXTbVN3iRvMOArM39FB5ZBlBfhWnb1nL8yeUxtiJArumS
wn6xA5Hk7ot22bvqzcLdcDAMAJI8ZsUpzRVSXCKK0Ea6tXBxa2/eWb+lKjxwnzkGxEBVMRDpBbIg
qY4AKhY2BiV9Uh0xKSzUpUqEEcq+LnX5YgsU/MQqv0kbQiWZpHIQf7tm6inUsAsbfxIdBjyTNh88
ue1bljLbsrg5r2n7Qvs1NyzU6piyERzfibVA905eC9MfsIgqBfQIgW9IEaLEqBocEwgAMIi04g+a
sI1xTS45T5tDzUpgjS7XWyi7PayzzLJa5IBa157kEsNz8hMzx3j2dkEwYHS/583Fzh6n+HsJG/ib
fpgcLsny7gJdGm8r02Rdxd+o84haW+jY1tOnzNa2q3w6/LNIPKn0gtuWNhAWQU2/BTBCmWscUcdY
9GVmTIVSbOxN/8BKGve1BYoJa5BpUGgdGGpVE/InJ5SxJDNnspFhzU2c6bL/lId+pe9ybQXkDaGM
R9nXmrb/V/0nGCHd58BFowpnqn8OS8k9Oz7FsX3QpMUJ39A/CuTij8EXE1I1njHlX9KZP4npzh0a
fVEhq1qwrCSFZdL+4etewiHWRUl7if5FMNrJoRdmSvgqx1H+hn/x3b4U9cCH1+x5d/GB3xc9WXrw
wdLLeihGVy5GQ1o3ArlgBeFkH4nYn4x9lJRl1FXCwcDmXTjsdWUj4QY+UOTd0uJ6ZD/ZdT+CPH19
WkUVMcwEgYOcQ/eQorYOm5Ynua6cLBjqccNhh1LB18GreGRMBzeMrzPeW5XAvHC2Ytr3i6ALBonl
6Fcz+Au/THLNSEutgVNW+4fYGgcH/y7wQ6KJ21WvGCftv1dkttbZGGskLXDlns3V6jQhBDHTHe5q
VMFB7ad7OLy4rFmLgwVU4tvuFmHYIQ9fXEwaF229OHxsSCNCsj6nqa1RJTaJPXUAdEfDy/aaOiyl
i0DfqgTmJy7y67SwCOtrJ+7g19GQfnpHOEI+sW840+NW/egVs0LnlhH0UZ8dtwIpVPMi9qB5BR4e
PVoaw37jO+fgBZzU7s/RB7Fkx+hWVZ4EQxu7yoaxmhb8NRsuzvthf2c26D12iBNVlFR5PPYmVSWF
fiBBOtwtQwYjUotISvqLK2ZNDe6gBOqBI/LVJs4MvrmFxDGRLlexfvw96/P4MJ6PplKLH/ev0UDC
Z7BGBtRGQlb4vXBfzo7yUk6JR8OHLUD6ZGWOtGwns9wh+VLpNpTrH4i2O0fQX/p86OaInBuI6vV0
L+Lq4sh4/JBXIh1LvBzzHJNkO/eZVGjgqxa3gREhxckm5TK6W7XueEhVhs3PiiBPX21mZz+GV1qB
88c7OAgx3tt3HIbIw3UqjRMNgLRciqdRHCaAXbz8a+PAgjwqX+knEdis8kdPoJVXcYq6ztS84Bf0
rgK+2e+sseJaRjuaVVLCceB22rH1Gj4PtYAm32C04HKMGMUrIAWNsXbDfu3364Sp7FXE32Ep4IWH
nYYr5ur7ZQVtLCEQjwnuYHeJ3bFOzfmydFHtExQDZnJYBaXG914o4GS3ha/BYsAsKZmwXNUE6sIi
cmFC5vN7VRjqTMDTtEWzwwjYUZLaK0adwQcWR0FOI2c1t6aAs8AB1O7tJ2lZMnu2mYFroFfNYjEY
IWDONMEy+FQ/uuFJrtWdAwEEM3yY7NusaB3nsBAWDhC/MuY0eYQkRyFa3obcRxM8nRmu0c40tuYk
I83cEht7A8ti1a6tmRh/IwLbb1KF/+uqzjKTCoks/j4db0PDKYNxiED9L0dZlJ1jmOGNPVy2yf5G
SJZRLJ68l+ikx5acZo89kIkYDnwgRWo7wzccvZ8jWBsgCtdBG/iD51p1Tu5poThcLzv2vErrcM/f
8JUKZ4H4cTukiOu4YkqT/TMY1SGajFeVvqzwe7ROGjfm3RhKcnolq5PyCpOLoASu+MoqpH/rR9H2
chEzsxFc8uKmbjSWMOqW8GGw0n9qUj1ewzpO2s0l/t5J5DKHmqv2jBL+iqCrWX7RPFvQLa7cCjIs
YdMV0PT6LreSF++0ikDboIlihNebToC58e8SPO5U8JcueVIlj+e4wzpBrnjuwQmYU3UWNOGZgxRE
987+i5RPS0llLtVDLYUArFjGBjEXoPMmjEskSaGA0fihInl6MAaKS9/SA91uV0qYFqrF9tyW/xT/
Oki0hcU1gd2nZys/yjDpd6Tev4C3VEsUUSY4i33VSKjThl3H8eVxdfHvjZBUad38BKV98JcJmLtO
ZVlJVwEYLCS7BYYGe07dRSLhbdlXiQE88sjNOY8GzSXMs8YpX4cKnf465W1kWJdYIbiVtBa/rkHO
iaS3xYlrg4HJGKg1QFT0+VI0a11PC/GpAdzUCJ4M+6bDuP21OZisVGIGsQG5fccdaZW67Cys2HWZ
vdROGGYUo3/CsYkwA6MmQfJ8rPla1dHUHNk9WhFWSRW2nYp+DK3P6mKrCCj+qsBknzu1J7iq5yWP
RqgP065jANIv3r83DuHa9izNmBw9Itf+hw9DnusNiJzCn4e3mcu8YCgorQ6DtrD8LzZ4t+gQ2Q/N
ri6DRHRkKaqcvXie9URcKHHh0ZsLK2PKgb5Vq6RE2FoLsPYp9YFYnjzTFIhKZCP8Wu6489u9S1JH
20LfJySXf78X00qe8f5z+wdwqWRT6XDvoUksV8kkB2OuqliP8DQIq4bl+hCubxQKoANhTfo2lzu+
038JygofzEC49hQ2QL8eSTfKhlXFSp5NqLTmRCZ+LiHTGsndTjAO3D/voegc1Yq8njaGuIAYF/Md
wpv6H2vPnO6Amxxn2Zy1SDZeRa+UgLsvKLLm4759JKsshcO+j0MLzPscYTOX5+23DsqAVH5Xi8WE
R5JJTaKBZSmh3NX5scCNeXEDI4Nxz7AhwGlX6jH/4Skot4PeatC0zYp1du9r1nR9my3Af1smucn9
vFEWZyskwUItcP9QRIG8Zk4fB5cw4d8ybiUijA+9NIGzmhbSBlej/NDQL88ESJzfpyYD58/lAKuE
AIyTXHPGs5Ec/1bEZkZU7DO7GVQa8dQ5Rta2I3ymG+VtaUmMQ0/dnyLkQ8o0zc9c1Jnhl8gyEhji
67sq+MGRe4wISGL/tNI/AXLrpn0rz3TGXpZUIlVfUq5Yf6rnIkVWs0seD+jDaV8iFCYkntFBNjbC
YLSsMxjRdDra/ZitmbaUM2A+jIA+xQh+5NUO35IzdhvvdOC9fzFvOLrOpCyfHEXrbPTMmG6ht/J5
GR+SrytVr+RJQpqw0NKfPxmocd/SgjZvBsQrae9vqM3wbdridviprTeF2JxuYQF/RI5AyUjIV4lY
gmGzogQv5Czm1SsVcooC/rSN/S3lG90TGJlkEQtoGitKqZFZ6+fGQRZ53+EXndnBqHKSHZY4muJM
TlssNypggtMOXJ/t9HSFDOMRjnHJ+642/kedwMT3SO3rTSDU++87Jgb+X67d4ozYv71SWjIi6fgv
c6aZNaxKMzYSy0gdywkRZBLX7hftKv6hEsG1XiL/OqNxj1tqt78eBzVR+rt61O2HHAz3qyKbAzUI
bY3LFBAsDRL3yWNVr4j1aYn/nRb0lfQAKI/NHPEMMJa6L8ERbXNdTpeSDCvCb85o83xBEBoMU+t+
5ovwvdi5/DgKBeg0KtCqvgwSC3aUD6MdxE/crsIEZnGBZG00iz9ZgSrogGx6Ij4nb2AMEpHJHOM/
2Sr3S5VUmutgJ6xYjuWAyOQUaowXKp5+pg0hZxFwfRhjeip9jXRmrhX1qbsQ5oiQecDnjEwszp9V
Y5uposyDrZUoYKQbwCQZ0Gf4P7yzcIt7JtsxOLNWPmF9eRXiKxnTX4jrIRB0732ZNK/ti9XCLWSD
fGNRYRvSG/TToPBOm+hL5xQe0MbBcx/vKsrNwOOOuWlJK/DLgaj+cHrAR+Zvc8cxJBAgTG5Yqkgv
1o4yh6nu2i3OHWa5ID3vIX/IjFZszE3TlGLa2M++qBJcT8+DRaTBHk4feOEZxS4hNyeZUfIr4cY9
5BbZyaVSW8J4cd/bLPRu+/Jq+CzwOJ40kid0Yesdz//aenIjNrQty1yIkieOM4ueki+WfTDdW6gm
rNYcJ6B+uv4tSwmP4aE3PGmcFh76XKT3FF+BTVZ44sllbvQUDiluVKYF8r4ln7y8EO0iMN1B358L
/OY0xFAk4VQN1obL0bSSjtqjhVlGQ5Hk/fhX6MZfLcSSqF7GiW4DuuElyNLKuEmPoYvP3Yn4L7x3
ppATWn4AFELibi88eqdlsgOpW3u2Z2PVO+qoC9LMTwB1UI7o+znzfAk+LK24zYrTB1j2OPdWBuvW
JIzriZ3PAwVZPf8jyfcq8SWXFKgJRm1FCzu3cSpJrwnwTh+4Noimewcs6aE0JUC6nNgUApRFXXMw
R6yRaUiUT3tK6Bi0TGskD5BrhsGzmsHkSjaqoI11Uw0zGMnc6hCv62JEUKHraml9s9WjVX45xYK/
UJm4Rbwl/QomqdTp/bHz+Z3u75BFjeoCs30mQpbEq25Temdp0cuEz9oPuuLE5omRUjbh2oiSHWqP
ZI2ELleYfpk8ewNFvMwh03wugor6UHjy+yRMzPfKQJ3HOqypgC/Cu+CzAIBEjEMESQKXKj4JOSoq
9u/o/bRu28NdpotAKROiiN2wE24oTDfkdWh8cctHelQ5QQ7nFAPhTBmSOqIb1pE+L+9mpciHaZUT
Bjt+3v4TJOgaWcsA6kx5VlXiIjO9LaNEAfTLeaVJuZEavlyLRqZirpeLnsYq6hNGyCtkJEaMmQAE
8RYm3v5yaMg7T93xT2ulwte3N4tcA/UdQzd3clujbtAVk66evum5NI4dcUzqIFzdKtNqVSNxaE0d
k3Ma8NKQIbhcPPUDjxBGKNwnHusBAqnk+Oht0Fbxl8e9LJVgkVDkZUBkH0A8EfYwuVIGHZsTpp41
fz/JMU1XWcf/VyddE6a+8pcazfOxbyoCU7BEHdvdLz8pYYf99X3jaV372g2l1Dc790tECd+rxozJ
z9alN3BOBxZ6ITk1lA5a/gTcqM34mp0Fi+my1in9PlUO/k7VHjEUbKSLGcw1KitJzOAcB8t9POjC
R+8arTKf96DiF2kWVJX2t2kp+BHwhp5MyTT8GIO+ETzzHnUqvyfJfUvZrJtAmRqjypqqS1E6KEjr
WotHyrqX/0O9W/B2ZkK3uPVVJBGlyLn+bEHbupTiHhgRaxs9sXxpoff9edbZbFowy3/pDD7xMdcK
9ysdM1tA3jqh2L+BBWrqCKfCXfhhoLa9LVtr1KZQKu0ycmMOaMQfly+dmkivG7Pxl1FXguR2wJML
Isc2LJUYAa03HIf+ITtsGYtjDAdbAP/KIy7Z6NihaTiMr0CkZOcVH9wkstC43Kv3LNkv1kD68LK7
6ieBgtfOPQcJBX+vZoGi5koRtcPu+mB1Wr0bkDSTOj25I3eRpX79QgrlrXKGuuPqP8nB9MF4So2B
xisfrrsIwNqD4da0KKg2PT3VR4ibApubaB0OQ8VGF7kuFHQAQun2Y4GcBE8E9tertPPmgCMab8PS
+cfA5CguV+42va9FR23iRBTSVB+ZQ0Dk6sUvcRl7mri6fdB+quCRp8iAhjpXXi0CsBZ0ewdYH7MF
LOYKQYTJbNv1mFqKMA04ELoqOL/W6rSpRjXm2DugdGjNsnPVynFB0Z4k8rGoojDV1JvACkm2x4Yh
ZMZQ4nxPNG5pquNMYyTunO143GLGzelWtb3CeL/GRjyMH+xP5VDCsVvjzg2ciHWNRJPoT69duGr/
ZuODSlSRY97MGB02INAdGf12Qjf+FSOI0XhhrMGGkBa0lDML8RNdoh8xT81hsf78fMffbI0Sdq2e
8YUCVj1zFNP8HWsEcwqSOYMUuWCxL+TO5gAoiGIUYZdB/o5rYgpi5tgBg/En0EKxGdI4RwlwFaPd
w4eCcN+fDiVBbQEzHlfhG69LRa8HaPvsUAg/WfWfef3EZ5ix7XIw6MYLsZI+K+b7qVkI96T10aHa
YEU/iDkvcPwX52wx1LxA3M+2O1Bw+4FIhppQ/X/sAAUHIDm8SCrnoo9k1lHFM+kZWowfHjUp5j7O
uFpeOpLgod3sc2UHoks9QBvRCFl2vGTSU7Gj5/upW483I4pQYC5yRVNOCKkeIdAU25mHwqvg3OHT
2gRsdkaGjeKIO3Cc4rM25cZvjR6364MfOcLCp6qg16QCptmzr42Dmt4lsbEWljEfhJFVV5kzP538
V8KUNYcmEgOkZ1GlsT2uYZoOl4wtsTeb2+51AuiS0PAEliavAU7HJeNOmDDWGYAa4VO/6pyeLQnM
RyP54ojd+LXyt030qhoKp4g8zwplrvz4OFWq5M7/xuf3EByGoTEWJ/Ep/sExe6ZqOYFDcQ/7uCMv
/FDWDlBuqdNMPfo5NxpA2ZiuQT+OJojtTnLc6MOe8Ql4aWOAub2u8gAADmPKSho1zB0rR67L0Q4z
OFHCYh/QfXx8ZDfaaG7lLcmHxGN5QVGVIhsmb/0bQFFtoSZtlV2n1bbhi1jpisipZ+ZBvpuzq0Ds
FQnYqm9Og6mTrDSU0PxJa1qv6UyJ5BQNESzsDbJzDvlDDUxQHkdO3zHgQexGLUJuKjkXziaOA1Za
Q913J970EjGsxEmWNSROWRWm1acEjhuA7//o6ubfFliHRyH+YfggFL4Tt0jmSLduXra6mHcJSZ6R
sa6H30CtroVN6RnYCzJu4caHuS+knY+ATQnJPXZUwBmmzDKrI8N1C+AuG9H9onoKDQ2QpvTSvaFJ
UNm1gvOjYtDrJ97gRbJEhP0/yt2jiPRqxF5ZttkQCDcqqmTlq/7GzP35eRMRJJAJenVvGO2HfPF+
w+6m/16uDXkHHS7NaxJYh1bS76sV6X1UxzQYCvxo4SZweBh/uS+WwpCwSBc340OnkcwQnKPBR0xp
C/sX1LVi/7JJlTRzfFPd1sQgGEQfOh+laC3U/iyRYHgKT/HZhoh7BWCJ8lzr6dDV1k152UzSXKIr
tOoE4jxy6imMNvsHx8r848twDERcXc8pUHNzni1djTbsN2mTLMw4c4t8FlBo7VSSgqg5zzj9arv6
VeWpdRuOagflP9JDJqRVZPBB9vvCIrpA12hY9D7h5GpT+f1Alb2eEatGoRN05cTpDqg2cZDXpnVP
bYAqQr7WmBVI1LE0UQOID0tFnjvBDdGRQcEvqZyPig9nZ8/SPQnj/jgJCZ6aLCzOSBagpV3CewMM
DmzTHhtZGshFpI3vUYCXhcZGmY2pdnKyoCaJkKkvcIHNYKxh/5bRW6hPa2xldMthJIGD2HQBBltz
amWDQ9f5bYouPvMM4vc0KGargDPuawwJ2uUp57UyF1JEExNIqHkFwS1Nul7HWNtTwKaWReanMK0z
3cXqz9/R7EonPmpYGkyANoTbEtm396a9QlW/KKcwp63e0Heth7/SNh5H42EycZAZ7X4JGDJR6COk
pIlYKmycVhaWP2QZouhGl1RJZBPZ8YZYsGZ5o76VqCaGVdc/Ka1m2OihB1o72bixRKvwCJ2OFInd
FKBJNs+UhzAu+sCwl6Ww7GMyjTZhkljnWcda9e4wFdFQP8J/v5lPcdRmkXssBCvblvdBjPcyVYs6
ijFDbx4ogJDPj83TwQxw7fQy7RYuu4Vm9OR9vEZlNCOmPspyMgHseobMIY6y0+anwQ8IJjUdSAUx
v7Dzpqg13Yqpla3u/+Prf5qHsVQvae2iMbO+R5OVO+M4MDHNCiDO8joE/8Ke0g1wI6Sgn6akxZVq
5v7TzPnhK0wKIEUckC0f1fR4iGESegnZr67lOSlN4MnupqMJa1etzfxz/Wc/YcHaBnbbt9qxXlC2
htYnJKGjsUWqMdCTCbJKLqvG17RGlcCZZ+Jf01I35k+EvQp3P6BRNLcBy/69MbKhTO6ABV3Ptq/3
VhwDenMDuwjhcm7uHUcneF6Fu24e+vkR81uzh21LNkgQ5sQsrK5V8bhkWNaqGnJTgn1rl9xabxCZ
m/xGX8VeRXNKFKJvFvrpWv8KwBmgBdHiNxKs6vLrOk2QsmII4T9wgo/RRucf8xg3V2wtLNnCBUZx
YSR9tCAj8hLELQG3KBNp66bAo3FA89l94fpNlRRGDU0CirF1sGUyOk95eNKhE/7Vw+M1VOrBFay0
3qoLcaHRq9vLq2sn9kdaRblLR7zavNhzUYaCh1dBc+RU/Uwto3l0K/e2tW7ylkvr81kJ+KxEK2uR
KAIKDWWHtG6/WlyXXwgK1CzfTJzC7UAZYbwc8g1kpqT6Eigvxk95uBzUYg/SG7m2qtDbBH1fEI3a
O6AL6UJlZ+XVlG4LM9crMNM/V7wV3iYSWonKFS1/SN9c9VaoVaiUvu5n/s9gwYFtqntBvONdZzM3
WFeVrRPrGKq2XKsDBu3rXQgF0Ca+Hui0nbn+caAaE4zucxWA9GTbH47EEz93nSntKsULpsAhylvZ
UE6zdMerZiTAB+GUJ6KW6Kq1E2fkhzrbI96r9gWwTHzOwBv2nM1BhBZn3jr+eU6JuEj25Sy/sZI5
NIEDkuEJpNsp5E8PmhQ0jQEnTqmOWdxv7S8By4OSmPPzftWo5kqvJjPngFoWcRxA/ai7fjeS6d2b
HgkwN7tCfjwW/cxWX9EvdK4xCPSkXT3fruPZhE/KBkTfOyOeomnJ2NAiXor9s7SSUJIk3OfO3kWO
EJ+1j3u+IGRAw8X10KZb8N6j05050xdAUhOh2/KKtGx2KnhiQOxYsuvJhExPH5Yaf9bsv135vxqj
OcJhD/pNO0pcPOlw6bqEkwq7PRxezgz+k11d6ILojImUhqxtyPxW8WdVHinxUVAopTXcriJncI9n
+7+ojcTMbBaM/bRIDU5r0+HsDOVf8rm8b1ZZP7jMvE1sWLletAfpDnvB/kiI2+/SnMaz7kQQgHjr
b2yD6k7ijSduQIsYWDLVgWimslxwho67e6PaGcPiTrzQDGHshdtvTQVtwEAa2WzqJs+cBatxeZcA
mqP5Ic2slYGC5Y0K2re6ty514knltJ0KXvH8OskogGIYFSfUvR7x5ame/kCWihc4cUaAfGeoA3FW
H7Q10+Qpk1nDPMHN3zXZ9Yw2yPAzrVS0Qv6Fgsto8cZuqBEw3gjLJVx81zQa+vHVvcAm0K5WZ0c3
gH50AeWRb1n/BKuBSbfccwOF+PLRVPLwNO6xVE6FKq5qgkNAe+n2vO4uTGpqCihWzvI3FPtcYjly
XqngL74KDRIE6nmqiO2rSMjJm060fsfZ0fH1voNe3q2yYWTJQtemFpVx3bsO2ohlWmaxD6FR8g0D
czNngVNSwCeaf6Wdvn39Ip3qXPrG/lcPMhmfAz5NEttHz2/8TGZQ696mZtN3lGZ9mIhWqrDm2BjQ
LPUsRlVc8F/ywa0CfKy4P4MWVCdgp1X6gHkZEfguqmHYcdxLYqW+Aq0Y6kxSpAhX/LI2YBeZ+C13
TFJ6SCiG0AFMHmu3HmbusxHFnp2rWBDN/Da/tSdtwVAAlRRtg42/iFCM5q9xeWLVKvzpyDySPOcE
mdnloDeYYaMeh5fDlwyZa6o/YbN2O9KI/FFdsTa0NieQrL+zL+hYNWO/6aEs1Xd/AlVFShPSNiiO
98kvfJofZIq+Vu4C2YnVodGKZALfIzdTKUWsBuu+aKe4d9DvsndSlurpRnMl0wcrBq0rcHPEU5cY
6PQ1juEswVYpobVMsC5c2sP8w+Ds+++ezWQUAQ6q6CV/4lJDMN+Iv6zG/S8DNjKnXqaRoZI9z40v
PhqTbMcZ1la2F3yIMuB+ZdlEBypzHm7X2H31kvb2PHQ8PXUIHqeY2+6+Es1hDJkrWZ5L69CSkauj
2kT8gdCaGqGt03cHezr46RoB4qjuziXBP6zi+2mGtReQWnxC0kc0EpJ5E+Kedwelm4Ia2ZOwoliK
VB1T4hUyWcdX7p5uPCYa/3HXUPam4zQvoMFVPAni0ZfpNteBMvnGE/CmcnXkALW8Aw/Uhn/5q4CR
IHTXPamgS+Dh8CQBkdOZCZVu6o+CIxCWDNmdgFhiQHLB//6PtJcrKMBCrn6Pn56eYrarqgXcwBRJ
ueYeXIyVpw5J26cZzpb8eiubbF5eoYkedGeWZ/8+44G3XOldB3Uk2tW9RHRxhXUo1FBLolIxH83i
2eZtrAbrAf7npKHaWduDpKGW3I7cU6J2Dp4K5DkSAKpmSXh9fMuH9B9Keile7KPgAH/iTXH2937B
FNnoACTeC3ZeP3/jxqMVhZNtsLKFmHl2Pz+JGcCtuP9dQFxviac9SkOAFdgHsr0m9+Kt7oKHeCx6
aE7Lo4p/5DyYson1PZA3X7+0LimwL/Tex6Yad9p38GFs7+cfmYmm1761A9VPyvBWu0/dLLreT30r
UlWIRfB+fYopLvvn2rXPVd7fnp7b4xtBG4Zb8shOaDrEcis07hcj9s0ZDGKxx3P/PpDonBVvj1WC
0+QN8FBLzO6YTpQwXpT64QDsaJy4D0wsvmgxngepbUHpLc60NZou1OJRnfThsUgtZtxiK2kXpPil
3v5xbF4YwoG/5k04B74zVt11O31/eM00iBWeou5AJ+vsMBb63SFV7f4YU15W0o+K3ijBCpFQBCJj
Nn16wEIjAiIkolUpAqlcOQew4dYoiu/K9U6iRxxmzMIBfz4Q3HUWE2I7Pe8xlhXmbE6qsJMTTvDG
dwD2CpG4anK/Z3InkyAPyZh5vqBQpd8cZxsNZASu5F3i/N0BZ+8P82H/8Yv86EH5+ZAMFlF0b1lV
GsAztRRKHUDN6UjszAtEVsPJYdFwX+1ifqv2mVz4+9YZXniTQpEqf7okCI/6OkI7NTepE8bvhLmC
iSaYeyWts5+gcm2Xzp8sT7wrXDqB86PmkzUeTnqQRvMjoJ8/epWrfsZdNNtrun0W2RMCN8d9TvB/
7YBvWK5ed+rLG3t18TFLgcg8r49hNKZhiFTh6RnKyF0Sx59jg5t7D9je/KbZyiF9vt5CqU0cAPtP
Sd0izfJfoO00QppvNiC3wG2k12TB2lv405q5nf5xCi3vWcH4f40MQE3/8vGUamvvmfhX530SZnnR
4ZUyyl3YXM+COKpyf0c/CHD7Hu7gI6PSxSZ6CWppH20LX2undNd8Q8qDxp4rK0IDPFd13iw0zCld
ogG2uwLvY3V8xrqCAIMYo6fUh+jbHF0Y/y+L9Yxolk/zpstFk4FxqjtgpnuOYnp0nU8mjoO1iKJi
AQfcv8bz9dl7kMpiPJnroS4FOYKZypx2XpGd4/JfKQvcH/TfS9zNoVv/c+1CMNpk82l4bO0y9wPo
iA5QPH2Gz6Qunn6FLEZAsBYAfYUyUAEpfPrdMnVZx6U2OzvSxGiC4OBt0vDQg0QBMUSJ7rDn1yd4
VG+42iArIkRhZZX+qLA+yVUZkTl+zitdEeFC/7Gq8f9KQGifMn+F4F5mG0xMnG5SbJhAc1ZLa7Fi
+oZ3Tg5L4hvuWabG/kPFSHFP3/voK1jx9quNpn/uKYFPu4HIv8WOzE1hn4ABk3qzJbw3K4dkkFSz
jRdY9IhJDppCYKfog5BQyj+B4C/pua8lcHQX9bwB1ExkHkRnUGkdMUGvdqeMPzrEV/+rm+lFOqOa
DcbGnt55KaQ7kzQEsVTZZ25idAhkkmWssRDyjrCBx2SzpmzLcJrm3EtGSZf137HMRwJDGdphQpt0
p2nebxp0cvDvOQtP/RndxKAzlCLsymAfYaNfcEkZbtS41CQSH0d+r2gD/LPWaLmObZgy00wWadOM
Av5QQE+k8xfq8Z5mG3yc3Bc7Cf6+kb3BjaM+Zf5EJBAcYqWYouFG29S6wwQ0RW9FOxPoD2f+BXOz
Ac+fDtRvDHegIiV0fM2Nw2bAg2WDeSVykb3u96AD63eT1CfXum04r70WiGXrHZzAa1b/vGPlqOyV
ehLqmvuXiy957Wn/bqc36MRy6V5LEw19d9RpN/uWNT7qVnDBsu2y389ZYX8xa41GHH/iAC2X4sVA
x45T5wTjWdzdfopjcuW0f3NynH+8eK1G4OetfSNq1OTsjfKgTG1uY5VfbMm1epabOfSjFMk+VjbR
1ll3QJkSdI51jfixp3f6w0Di+t3CMb5lpxx458DBu8pdkU66yojjL0BFZCvgzZqYC2Wt8cUxw5nw
zE6Sq/l6BuzBElDoYIxkYA9MabDuv6sYovJxL67hZCX6pty8eREEx+r7mjLEbui6GqyCY29Qcj9F
b33U1t4HgUOdhBvMGqYNwPhZIB2zijmfyWo5VBhzoRk5CU39/VEkDUE0zmU2qldI5qBZAqouYZfE
WvSIDLnQ1bkbBNxJCcGIZdGbTjhNkjfVP/8pr5ajmhMiGJONGRG0CZNr8KdqP9ksdLSmfHclQUS+
xmIjDjK15KHvS41gVANUWSTxXBaW83xZAdCA74XAPsHOaC/FXso15JkCnSxhrk9cAvBU9AMA2Kp+
v1Iq3Qb0cq2JnE5m0uFWRYW8qilI1Fx186NClJK7dR3G/8NX27OFikvGDL4Q4QZGAAhRSC+G8fax
Faq6TPDtqYVXFuToy+yRGdGb45Izqp4+7nhLBeyqK13xw6AoM8r3TUaHm9yAQ1QOW4Wcka5kDvlw
51EW6iearoVIeBIU3upXBJcVBVlUcU0yQOesQPNKl8i+t4KlFYWQuPPxbC2X+toPOlvIuOyAZlDh
V3iUik2UXY/WZI8/6MwoFbwBpOKmpowUl8W5BtWzvpx2EAgzsawW7sfdxJNSWlklmXe3w5W2PHsr
xH+qIwqLMwtG3U6gN1IqsFqggkqUj+spcM0PEdMeTOsqyCTN+J6GxvBSgoyaLVmhg3sN1o7Z4LfY
jKH/5l4y+D3Qvn/oUECQyhJ/Tejjf65zoRWkyFA1+cPTmQULMENo9M3JDgf9oLoOtsTzbyqC403m
VIEVpYTwDPHfV8YzKRvMfnbSA/HtWauwQoPV2+tKpNhnJ9G41tNfUm0qmvDTOrzHWddOt8qkoAkH
lpMGMNFjNP62z3lfpjHdY/PjxR8U1PG2DT897X+or8GoR7nThy8dPMwUgQId5xM8ew7R3qmbiQEK
TEtqbWxnjN9qP1z2IFGusYY7XKx6Je4yjFACCVlxDsj2Ts9viLLJDufkLlMI8nO8sNhzOez9pdiF
Hu9sd8M62+ZZ4pfPzoZhTLZURK64T9Qn5bucSWloxu8hEnqmISOQZTKssj1Cr1Z0NnhD/d9FTHJF
G2nj5alejjJ6rALXVpMCnbRprVs6Mm+Nz5cB04XsZJIsgeV+OFwH/Y+FzLoVVRUi3HljPH6XO4KD
2Mj5LV20AAMt+3oZwOizwvbo3b3fZupX4ngMdQdkVN6Usomxd2uS6apgJ6e92rvYDaEEndvNtr5n
Mv9awSwBPbAKZ3+/XKN/jfmBRH1RmBbXJ6dHsF1+aZ6SI/bEfbwgfjz99zcTSoEFVz0Ffn8pLRh1
rhtvWLPYcmrRKWg5R8UQu+dvuZUFACuh5QMRrA40/eJWvf+lOsbLbPxbqZwKLV4gK8+lS55ezHBx
ib3k+lUvENcUQo9wlOVXpNJNp5Bw0VxSTv59cea/fEGszgSCH+q4/gk+JHVZLW2E7ZpR0NPMZQD3
TKlDNkQWZ4q1jy7SIYVXKA+Eftk73zvzhwVtozLz8TCkuElBmW4mvz0ANq3zBwFuTmbOExWWJPbn
F3HZA/RLZ/4mAOHLLfd8IGkeJJbsj9AVLPpYyCcRDl2GauA6QCUMpnuUP00r5dvk4Oyf6YsoMga9
CqTK+YhUc4Nj2DPvggx45/tkTuSLUlqC7S03ENGtYaWD49QqTejA27AvR1Qlic7IN8T6QXyH/p+M
9zrD5rcStJJ53Y8znP5mEVIw+kSOtMhHChHF7RDbZinwyf1382N6xof08Ih4CjLdwJi8PE/eKqll
xdpLxxUGWEtfc653f3bDVes1IJ1F3mmLdNWVqySBItoKWcvhI6a1Pa9ksqh0kr6zsEYR8NaHHcKK
ejUchyfClBbAu4EhDf+B9UexOVUZVp9NufdAD176VQgu3adY3C/0PyYs1A3WMCc5v3Uo5lBB8J47
iwE2jrPcT2ySV2BvsfiRRoadET1NLlgBIS6eg55dg9omeHXLkQvdO1QRyKBwUjHVo78U72UJj91o
u2FFZW/blOpe8LEhVkTRMdEJCn3cpH8FoIQC4vW2dY3a2klScqXHe6HiUxQ9ScHFsUMC/KVsr0vX
QGM0kRUS250o183J2C39dw7F6T1G3/B5yXM889qfBrwNb/Wr04v4LzGezDkl8+9XZVzXHVbHhDE4
IyKp0MXlyxLrV/1lmfwLkqBj2aYU/0JKkAYu5uHoiYT0i//3TMZXKwaZR0R/29H8rXUL9dnq3kHU
VeY9Oen2rF65QBRsmv+Dm0PSNuT5s8dffcNX83DEJC55ed/wjqeg8yRHKm4TXYvzb8U9r7TelOpg
UOAWMXyHAsIZ7ZsroiIk2NQlQJfmzavtgXtpit8Uazi5CuY+9qnJ7jntN/LdHOwN26O1YMlnNzBq
xp7MdTJR/I8igaw7UaZRqN/+ngVMKcq6U71mNu8vKpEtldEV8xopSQkvkp0MSec8ueADzW7rrc86
nF/j/fei5GkqPGRrKmySnVGqW6eYD5xS4yAjU8aStnnH5ibkDswqA4wNoifEXNFf8U3c93MM4z4E
jn7N5wJbsN0ofkO6iTbeuhMvzwNKa7B+rmft1GGuofksamUM9eNs6uKTEOHUc6ri14tjKl2IYGnj
M0dV6gSpbA1peK2L0vx5HdrCtnFAx+T4aTMKHaYoOehWNJgQwcmIbq/aowYG1gZHvsbh1dHlpag/
tPT5rYt4KGP1Mfse1uNdz6YqKXNUxVjkK/+p8skrZH1qDRKaTBfdU6Eo3Uz6Bz/9fnlnmnniLeU5
QGK57mNO63J8hAYZy8J4QhRPTwJsJdl9ppDF8DrzH2lo1nlCDsBMppY+yQ7xhWSsFxEBVfTJMrXb
tQ/3UyOftQAw/s2GJBvQvQ7aTgOlbasAz7jXhtbt1L5GRg5EvGUwgqAWJiX3FfToEFQKJHMXTfkX
SNdfrs2V6UcOV6wSxR11T1hsgnEJpeHWn11p0fohtHK00IYVhF5I54sRK7HLlTUfLjtBDbbmCxxK
klTdKKCIaX24JjraQkW2zvOAIIbQaBMA3hbuUYZNXjFO8Smp5DSqedFK6nsqeuJrJhn+iKjeqCbY
wzZHRxAhFX8FB0KroS/hJuqnoAblxM9vLogEFmvSGK9onpNGq9e56H0C0cn1kFzlFYF5me9NCQ/O
0h/We/8IFtVxjB2xQ7gWaRwAgLhaXdy+LmjoASueoUwVwxBenfKDu6ld/5PnvOlYaHBhHMNl8gqq
nCEivh+/BWWZXVHfqBuB8qUhZ5jFBvdiAPjiLzu8xtRRHc6FmZBmLn2F9lQNc7ybslhr7Bq1z/kq
M5tRIeKU8w5D+UtdR7Vj1HakJyK0FZHV8h3ZPbh81wQtsgkk8N+t+6SiTvjmAM9nCjP8cyl/bXYe
hsvlzSVWM6Z4NGdqldqUMKvMovlTdolTwbLg4U42qY85cyKmoQCHNRtWndbTg4jePr1L7Kf5QfH/
g7KfdE9Po2GtMuDuCystsG0lWVb7vZngvgBPMMRmfisDq7uS0pgjVLPJqsYZAX1wMkJvRIM5jtA0
5ACBw4Z4OAe4abVf7z8nEe/7fb5i6oTIDCWLySTEZj8S7EaIjXAuS3CHhtyNTCKZqX9CCo6WUi0U
7oG/OibqKpevlH1nquzGxcVl6d57uupIrnTYZvkVjwszf8FwBZib54uqIga35FXHjrUw2j0zCb8l
wLEQr9XWEhurbkcNxsD3ee4R1JFF7m2gusNJIl+JatjCITN8qrLVO2MHRLMcq+GkolkYfgmyAJlQ
t59VS7/kSm+ImMe7l7dtBQXLDOoaVh6SHEWoAO4xX2FExbFM/FFkpDmpsA+tp02tV2Uc8Sg6JGqH
MlwCxjnTkpQY+L3LFDxin0IjVqJhzYAFfcQOPFNZFsuWfRNFM7ShfrA3MXIovyRPtZttyo5aicH7
Ufs20mZVWi4NyFU05306jYKSJKd/DG0unnOuVVem66jBkp4KUxCft6W+UanapD0+oAoY+Iy81UDK
FouAk3BWVjucV7VWifWLPjwQ6a5q1qpiJGkddu2JYEeMnhRUjBgM6mi9WK22WlovJyNtxpHJQjsX
rqedHFdKCY5J2TwxHJEq/717QFp92DzHjfMTvGeHC53Ohp1xb9MiVmo70xgYHHEKYesGUxsFLmYa
7EzjYtYkriqp0fPssf6VZkQspzhy5bxWI50u1Er5hhkCuzlHcKvm9Fa6trl8MBPmV+yRsJr2+Bk8
PxT+zzZ7jKeqViVe4XX3G9RQO1dvFNIyWZDPeWMtriBKlYcYK2aSNXcZFsgWdlpO8FDh/0vxM9OJ
buC9mV6QswFgetESrmlyoJ6hq+jWAS/f4YiUB04nSK9iKF9vtMNkhHR3d3jwWc9g9WAG4/UZI59C
7fIj6L3aCNXrD2ILPUz1Z7jKGQylN2KBjDa2AGPvz+kPDUr1UmLwPPNG8pSuPly0LvTMUuNRWv3H
sIZVNlblHd348rhI938lju7y9tAYQew/pInKamM2wRx0fpMIq9mAc3hO2SLMYynC+TnIyaTpVCj0
9Fb72BWqmnIhWzIQDpJfJcu79xbLVeHgpQn1mtfUmoHvwKxcqzOx+TJ9bfEa69rbBWktJ6krPa91
0lvSVL8WCht4ruQVh9UipMxYf4hfof2qKccj3AzSBZ2lyteqWb/c9QM/zDWQCxHoNY61GjC2IFbP
PET1/js3pMZzZNG12Vki4971DxenKzmSyFaR3oGlG1IxMkvaJCmZDUpSAzdQOa3s+HTeN2VnMbdm
uIX8uPUOA6x9q4UJ9rgLl7/QSPYlAerfhLz7L/LQpua1liBUYfOsrYtKDwH+e/ikdQABbiwNq4cL
keE4L6sN3hxZbEIKRic8KJgotyD4Gy0FDCMg1rZUWNXs5aGkJsx4iJMecHLPUkqeYunOEKng0Okj
QJ2qVJ//EHb0/DG46hWuRCVG+3tVBpvCiT1ac8snzPtk/tEcnFScWYnQplZpAWNRiIyAeZ6Kvzkm
zLtCmfcXcbLzRw/uDqZ4/UUmhEIBd66K//0Ggf97xT1qS+q7dm2VSC9QL7LTPqAig9h2gP3sbLna
yY1EPHUeG1p+BOYHHGTqtGqei9aUJWgxMZQGRSTJTmxqfpQo0KCowYBgQ88UTvAJlAAh49AZWBm+
ZE4kjXaFdxGMecnONGnyaUdz7IpwZ/oGNQz0OTna/05wy+zrLsTMddV01EPxMCBBBMYy3AbtRxYa
guvWWqRH+wK2MLHg0bmWIeEe1HA7ConIWPh5kElfXBwOC3SZ2iSmjwZGsaici3dkGOQPuabO7Y24
Wodyy5+4dI7gUmfxfMMQoqsovM72J9YJf9Fyt19b2Rat/f3ZFwpaUtk+f1dRP9ZVZ/0ziWu1ASug
CQBFPIJHmR98bq4knRfzq/hdQ2oywD9h1aCoskoniUC913fKIPkdFZakLrSbmCbelP6gi++qbawx
CH8S1ZxMqLAIBXQavJkrDkRw+qOxkPUTrGeBgrCUH/BEM8paHe1KD9zrQlQs5Tclk7etb7F/9Hkj
Iiv8etjMAR2yBaD+vxTDWe1H6u/2gywGBXVc41ODHByy5wFE9MbutO9Nuz1dwwbdZTRpvAIkdMFG
K9knhb2D5p6M24PfrIbpqaFG/nfQlQ7TmQYex4oQIPLZpj8fripNy06e1RiW41ET2IiFfIF9jkn9
ng1zsZereVNNt+OiL4jNvmQmGV3ajWZ8j64JjSktyy53Gk4e72JLUJzu82TJs8wA1wtdZVMIPHX9
igjggxmndzJ6QEliovKurEWFhDWIJP0PWLLO5jUHYrarLq9bBb4JVzijk1wqGeipme6vyEaaTPB8
kagZzwBkQh0eZxN8VndvhMRjuznXm9IWihpI8u81QRlxVbyPT6warZWZDI5xtp6pDnyqsHAEKeod
cL1jVi24uFYvZtfY6v9U1mO26MXL29jJxAQredbE/dc+855Fk0+4fiZYBcOfGfR5Hb5LWrzWS/GZ
G5akDbc9lJgfRfJAYd5kmL4/MIN0yb3V7frB3xW3+mJKbea1BsLqf76o3VvgvuZ5cvPyUJdPEH4w
vcjbY7iTlZbFWu5/otLXFUxeQofiLzfleotTaxN9gewI9/ih+rRNjhc94SfQmwuZ9XTPDwCKNRYg
/otHaeRroaxhdgu53IYBq16VKXXNlLNJD0M0oADwq1YEqOLYGdZU44XX3QILTohtbr+tuJwGw8zL
Fljk+Db/qdPx7X31bxBR7JAS79Z+5dxegOoaOOKuyOC6UeIAoQEl8I+3ZulPwxcFL+VPSKL5b7lz
131pAHnyzNxkOyVu0hMIgsPKqmIXClgFbhIc2nMOz4j1NsuFuMkcjACLsedWFU3V663FT9n0Khot
oOmdusOGlfiCSt1hXlZ0iigyaIWmb21ozB0Ap4G0hIur9pVGTRf7D7hSD9nEYAMQIOwrhmeuGtXP
G9eLgr2WXwHH40vOBBu1JRc4f+HjNefN84SKmxKnQ7QiBerj0MLk6FwvZIbjSsdwPW/jw8DdtX3d
t5Ukk+oAciumm+a0bAWbEEcBgYWabR8tkHJzn0JwAL/waxt2S5/DIcGA/Wtg0Q/5cRT+fiS94F7I
br5pWAD+YrTK94VUqgLzJ0YecVnF9vJSok+6WyP5IACQADxMet1+MIPDZ9wjhCC34Q3kmw+ILCMN
y0/awYgV6P7H4WWQgrk1Fh2DsCh5xcoLjwrETKVl+T43Q6USVu4nS4MtEOf4HslYoxyBsNA1eJ9d
Hvrtk3VcSc/nHZjXJ5oD84p6GpV8ByqU7t5SNUinSB8D1fU0DIiwaLeXRlMKIgwskQi9Sddldrn8
Sp81hcXVF3Nlh5DWAhXM38968Tkobs0KnPKHa+bQpyY47zl7c/Oqc2whiid3fM6fQgzqDb69l58u
NQfyQleNZqi1nWSYN+fyGhak2w3LhIhOQGhstKHsdsA/X6FCvBO6zFURydTf2M8TI7Nhv4DiqT6Y
4VaA6rkQfKz80Ngm0/R4JYXyBpcc1SYLkETcG9S+WbTeqJyOQawWiF7rYtafsphUoRxIcMECFEQX
x+Mg4DtNHK75LhOMuRTU0OBQLRr7g71nizLTMhmLZFv+M2edWpJwS0YnQhhhHsOgSGLz+ggLs7wW
CZzaSnjjeY7qm1rG8LQxxOd4XZAver4cLokFb9t43XbSNSeht3T4zZajW+itaTUQY3HZOFo07nM7
hl710HGwdlQF4iZsYOhDCxRfvG12eZPNfbg4AVqDhQl0TDSjIybPWGFgXLSfmXuvWLii0xQKhrRe
oGhlfZW/r52WfGQ+mE97gNpQ7tp8aas/6BdI5BhRyhGWpsjFYJsUwaansRXWN7EGartIVatLdEl9
SjC4Wf8GwYCz7ACoOTD7nZDF57hrsHPLsT6z/1HuiPJfntjctLyUeyw4ld7hg6Ec4O0dCkEZUwZo
+hfscDUYNRrh2ioD4FzJ31cc5hKVDuWJuDVErwQr6af6iscDK9AQk4F9CbOhhWDd7d0WiJ6+J8wg
982rA0MyBLbrZy4DHZ9kxF046yWYYQRssJJNwAGnffUgFNqXyQ1U3QgePXbiVuytQIq0vLx+fAxG
5zacwK1gIXbaRdpVwhmOhWe8quPjdXoMVbiEWrklaOdxHAVUxPQmTF8bHJfodsS7DZa58MGZaUxn
rEAcEWJK5nfpmgQZyFd52OtBfe0C0JJmonrGk7bl69fSMT9ZiZa5sdSEljTt6rF2xXB0qgGZUaBS
xHuzdyGIsX9+RAqCBLAz8tb1UrJsg+S0puLvJwRx3ybQV8w6CT4x7MuZaBg/SduV9Sa0rBGABDds
15/Blenx0RMQ6LZ7IgkiXqwiPYo5biqw/Oa3CgpGizrP0Nopis9vzaSHEqckswvaRtW9bxKicGX5
W/Yq/R8hp7DyZiBmpQwuyh4/0ETIuqMRkE9yrT4W+QBXP/BxXsfrKCjNB369eh24f4q4k4WVMi9J
7ZHM6ikcg4GnFax6GYhz2GWihIKA25N1E6u0xrGBKCX0qfvGdJv2dKa88A8X3+sdUj56fLIKXO0c
SNWfTaJDx1zFMakSp+LZb8KjY74sd2ebmnHQPHo0hi8lMl9uqaRx//xgUNj3jVXply7YwFJ1iyEO
6nK4x4hOxGIXMGtDrbxCFU5Kf+Sh1FK9V0Y5Na4gE2ttB4KwrEBFmmEkpP1bPGTA9U3m6VUkoZ6/
MhFUvw4bODFkxP6KIupNFZxpCga2E/EmibiGgpcmZgYgiC4rkZteylLGvaiKMhDxWfvxrX3CNgTM
LplHDSvJwzmiffCoRWXg04JXc4FXYZufYM5Sd0u3m4y7sLi8a2H4Fy6+btSW6N4Yn11jCPH87m6b
6hWddgS1rou/b8CdkhUPR1hYEUMCqCryZPgg2/ByJIbZrw3kvgwNJ2WXcrwo96nYQ21Dl4H0YfBS
BQyLkfyLZlbFWbDLgzlajaccgyWC0I2WDJkNDUKGNk5fhPYQlDwWWTHfGLs1rzPvD4D1kMWsw9mZ
p1rN5iSwRtZj4/yx0tBPVJJl4j+Z+/awKPfKtbcu/rF/Ms8RkqGTZ22whGeO0XkNX225ulxPhfd0
pssga5Uk3ActH4YaCyYVTpTgK842WBGLKFE3vZfEXGoQSOYR17Fgta3aYaRcPmm80K3FLhpfrMVb
duZWe65zRG8fycO/lUoXiNyeoPKU5DLs0WT1aUGJeVSMHmPfgEcqxR5riZJmwc++A3Z+k75bBrCy
m0Fit8DJrE536V1Ftp1AOVEnp1ks/L7OnTV8y+b7bGmBBXXK7UW+TvrF4AvNP6KKtFj7bVamKyge
zuJGsbbN445GwCxWoSLyTxu1EA1e0yatLzeevffc0gXmyQURelAxHaURIlHKY+vgtusqK6r1/noF
Y/qDgDXgiTX5hkNe8AQmm07+JnwfVoRkwJzTj2z0hqMqJ4ZQMiBWCPVRIQnoY9hE2WsBi+Ci3qQt
QbFRkerUg+imzuZk0ns0BFbibCbUJpkpZjZco1c7+3kvcHH6/xtKqxxIhj7K2eCsXocwII53i7aG
PJ/7y0rrPtWhmrk7v7sQq/L4GqhVz99hNI8YUxHYGAKnqHgUUpDKlY1KLrKIOvZ8fj0YtHxvSojC
c0mypp0Ykje/eU/zLH8osZp9gw+L1wRJf7P27H3dJckyZJYUtCf3zXhGa6OiG4JhG03QwIUZCAaA
GS+OcILuViLGhFLKMeYxuMe3663JqFzlPn5olvEi9EFY5xgMWcVejv7p9T97ulVQDXUhaFoQaG4l
mAq47sAq6fh+QbxJA6SEDaic8vbD5Z+NZo4Z2E4ry5FAtXMz5dGcvXsCsl8bWuEVdPrm/ODkqiT9
rKWXDrB1NXzDCVfA9bwtZ22cbHQCDLVdEYdJqGZG/ruFM+1WHZRN6ocSmJHeW8DEmQV49U0+HcgV
97dshzTGww6se8VLTikxWcmCu8D0qpYEk94kMP3eVZMc2Jwp0SHQZWxUWFUn3JT8Mwmcky7PGb2z
ZLGe6/r0cdeAy/rU8C1TUOHyP35Ev6phh2aTspNjUQvoKbX2hpioGO5hHB4kdeYZOUpFXPCaN2Zi
w9HR5MPY9V2JRgj/xOCGi6JEGnU9a2rmogebGMIRe1INv3YZ7CMX/yArFPQ2s9t3OgPghQnT7z0u
N81sitZFVC52D30Hf5IkaFZKoYvKctZhOXHV1HwoSlADqyhH4RCe66Bdykq5B93K9Hhv9Zw0ff3D
iGNXJOFNYH7vrgx+jSvEf7O3p55gTPwhtaitLIXYSF7NeQK5POYNyO4jlycCfhPLp5aFcmA9IVzO
sBBIUxmOATBE8961QEp+PQXpvPQ1QgLslqq1N5b8U3OIC/srPVF/suUS07wCc9A3lkdOdqKH1ovr
04+ouN3k4w4njAiArdPvKWfO0AZLDdrTLqZlJFR2Q5dc52q3iq7tyMXnGyYpRnoxYMIBMDJCKgsS
mTmborZtsiuKSswZQntcFcDhn1EDOFQbHBQqokAw8EWkYUsVT+GPam8CfGTLb8BkwXUZe9qlmXAu
gmxvVQhWx3WdKpnKiM3gY4Aa6g+sNhU7w+/gl+iBuGVC0VPsp6+90erBNBJcSjnlbXHY8DVQtRRC
HALxEFQfFja4PZ30MygV6D4tYdDymz7/05k8kpihD7G0gHiP/dAKVWs96/ERLAL/VFNwaiZ0XEbR
4nvmukhj2JPkm7qVC78i+oc/DXj6Bb0SwJrV+pG13QQS3wW/FwNkgtPcO8sAh2xujBO8AOUM2DVY
OpXfLPbK/srafB/y/JVfZHhLlg3e3XNZIwJM59Q+qfnSMSYk0N3IDhfz18b276AymKOq7ocUIZc7
/S2Oe/r4WEyJ8ZVlEGnzELhFjikEWG7GYLj1quT+KKPA1kvGFdYbRKELkLU9XeNgt5u2ZOAKjzcq
JGXQZCiBNOL4Q7ctLmwWhK17spz+WXLN7To/t4GSVRZ1N3JfBA2JmADO7z5HQfF3IEYDhQp0ajVb
QmTqeXTE2s1ZIgkEr1bTjZ5QzUgmuu0d/XeOBRH8NiIY+D2fLWC1n7oh56JE//sCTQwatV/rO/Y8
Ntr9azxJYXFrFg5yQHzHUKEPkkdz6g/ceGHGfKBqpCaVbXRes4pJOFpx2/oSl7hfXAEYzCoPQWaW
HwzIbk6OOIc1Jv+IWTlkNz61MyLlfhlkoRaua6NpDd0nZ15I2xoxqxBEKwycQ2D5wf+esp3Ul8mk
2Ywz5Il+c68cf4pTmZa1Af+/xg1QKJiw3wMAFT4JzriUkmHAQ5uThy+Fvwfwb+IfnhdlKmJkdgC0
QK6/O9+YJ07u5g2shyu1mdDpaYJkz7ytJIlsP/e73Do+5goRwrkkF9CxPb9MDqxuFqbqFGe/UXDU
rS3QZ3TiFeGL7dab0npGII4tC5lQfD9sa4wFLWz0GCsp0skeDJxanYwl9tucLg5tIhFcbaRC3Dwl
prefpelqDP9xULDQbEgolB2uvxA3kURnXNdmfSZox1PUwxPA0zd4TW5fjyaj/yVixm8lF95bjWqN
479343lPZzar0pIOW5i9809egxLK8YO1xH8PpUnG1YYDrdW+9a5et6fxvVLkAVT0rj2NepW5B7G7
0EOe1oLdnQBBP+Ml//4vYxSfl/V8w6fYTvd8CoU14bfoajz28ab5CB4EGzPB4RMo8gQFNbHF8OHW
rsDKn+S+/L2Vyx1LlF8LQvFM1kyAMTcOuyoKADxDGMcYshqu53b+7GOU0n9fPgI3nJPlO6D2tLJG
iLwF8yExopL1TPmDYrG/eluoRBEit9DC6zFSUFrshVFblGp6XYnn6b+h6IUdvPax/qhATk2tNzDo
5zkfs7jFjps1E7xPAdQoas1hww+hQUE6BLrVTrxs5e9cfbF8vnelEgn8OWUSIf9mUnjpSy8a7j97
Lqz57M+WfYDKbaFrYk9msUIcQFPaoZgHf7KSbWI04QMih9QGnEwY8UrOp6G/u+S2TL7G2W7w7W00
KK1SFmoNNbU9rTs5xsmTk9km8yGajlCwle5RXNHQLSla63c+dnihDwscXDlrSypBRhrnbAxw1vro
OJOKN7/xpm90LIkud9Qo4D5Wv6gVzRplQ2tsnSFAlA/dHUIU82H492Udj2NJ2aW/7X4CuIkS1B5/
CjyxnqTU18LHVqvJcKnLyT59YEnJKSbgH0tyNB7RF7IItwNouM33JeQB8nS8t1aH3buDpWLRUqpg
49TSMRzNnHNVfjlD84S3ZY70iLTszeHgzoNRbws5WDFbEW2QcyOU0kzyUGDd8QYtmUeb4jUqDv+p
tmNThjYxxrC7xRrQOO5zh+qD4sZM5Yik/vFI1YcRjbHPbAXD3k372c2OYppKEXNAtTtuO4li1sIH
0ayPkpgpEstXq/C6twVondWa401Yvt51uDlYsYXVXT3BwqLrNBA4aQj/cELWMn6YwFlAj8yqQeU7
rsThFWtjurNWStAJk+waJ7NWVtsgyjHInjuJLxDGMyesj6EDRpSD4mLAwZnkHsOiIHd+pbyjlmfa
qSyP1FMydbK02Rh5ZhXX6fbBhxGQGNsTGFkQHnh8Lza2yyGD18V1mGIRATB2ktVfOMokxA39lk1E
/9D5N22qWJMjulwcLHtXjbkr+pnn36J3IyWkqlvJldAYJuWIr0cl4WvAdzdH1JcLt7YneQUzw3wl
opfY9E3V5uvI1KE/aJtud/RJntcQ0b//VnzS6HWI8bEQiTBfNu0nnZUsARDre3V8+WuuALfhtY9m
7/syDk4ppGCS73PgzT4NVfvogL2gUowP3B2jhhZEzxPDAc8WmU5OyDWy9UPX/8VvOl0R5/Nf0NtY
ysL+FdVglE01AA1UTUc4pdLOjsrkxwaS/55eVioEAW00FZ5JA1cv9NghcuGwZRsb/Nl0NDR1aspy
Oj5Y3ia0GDmM3GLrSF3A/uv9z1LWvSuwxZwBsqRiLiiOK5kq2fmMHY9fAoi5YSnyNkK06D2UFgIP
dlvfJViWXKxqNNFsnFWYYi7xN4TWSl0LRphkKNi88vGF7v43lJSoKhSYEkQSPrSKWQ/uactHbPLj
qMtVqtKAsj9hrccBJCEbV7Re82KSAbFSTmieZqfpr4LzRFPw7dcyP+Md44zYP3A4O18HK5H++MYJ
W24Et8WaEYYnHlwwPM7wsrC3/3tA9AhdaCds1zMjGxqfCN9V0qvQipN5zXe6Le/TM6ldHF6bM41R
3Ns2482WIqchIr+rM1WC6rLo/gEJwhWBQ2ApOuXECsb2w2FJA5TBEPN4DQXQ4IYDO+3NJhDJdAp0
m8S1m0n9h0j6gv7+prfoHx0n2jtO8ybqVqyN6T8ncIkMmkQnuESNyHUyrTOPhsTyXXtEz5adKmDM
NWth5JqH1bfYFOa9nRZ/NSn4XBzEg2TLmR4Y4ITS13l5YGXxv15YejXZOI74rY9dopTxOeiNu1oj
jwhQoPlewfKQRRH+jdwxOS8U0Sx1Plg3aRKhuoQShIAqTDeYggreM9+t7Jf7PSGSrltdovy8SRor
gX6eDaAXT8vfu4mUUbeVQJPqr/lWaUQBHqp9NzAVsAQGPQ+Is0FSe5KYOuW+L4ZC9VFPsFWqPIk9
u6y6a14B0mFbmAnqgCFse+TQatMfV6t3Sv/95nVXeRK87A/aQ0sZMiBUO+BzNopbFIpZN2zBQa6e
5dRhGLu915MgrJSp1K3Q7cyug/C9ISvSVQDBvw5Hq8alXmZhbN1b93uNvGx2NN9stWtHO5nsgCw0
9LgQbhTuiFv2iaJhUkcaEbpXATBIOXBjjEPQ+5F+0tGjZ659Amrj0fB9sIJJwkhtKAAVLFAOOzS3
Sq0yXM0lDb0Ny7xkFR7oXfZRqwAEBZy0FH1djS484tUTmw4vS9HrcKq/TLyzLTzcgGKCMvjYKBNF
xPpfRA7V9mTNDvhDhNbm6gOyrfZomR8xzOmBtpIBWODeN5XNfGC3IWx1pudVvUbzYuSwGV8dyLhC
JX3Hl5aabv/l8fekCczds4JpfjpAWxzf1T+R/P1hDl0p6yYgH78IK3GDF3lyWEc/5KXbY/Dg10Ph
fG71NNc2ilkYnf+jcsb3ojRYZ4T3cOCYg6o1XYvaCWNL+KySA/5Os2CufXQJj3lmJBE/4WF435FP
N7TW2W3DbZ9E+sa8GR8FjHyH6dYjfSAZEjNmoT5yG4442ROY/bQZtk6fHIhGN2E5KvQrVJEjMSah
2mqykUh7hYBFdnCp5S5PYF9ngHuZ+xPtaFvvyQh2dj2V+CWo9Dca663dFbtKSvoiKz1wcAARxhEj
Ta5dJ2a6XYsNejZbqR3Vo4vyTtTV2DyhvBDvXomWI/Kr1x/kfPH0+FP2EpVjDR8m/XTYIFfNNzzZ
4NQ9qIPVNur7yyYPmk0OuTDz2m+971UdyLepL9gZJTDOYPotA1kCOXqH2rWRljW2BWtjO2+Xd6Cy
cs7oxAzisX1t/bEAdLOwvbIRaGPEYTLWJu6H/mJLlJL5/NUjhG5OehpVFq67F25Am12Fw2IM85KA
DgY8NA8X1vs3/wddvrdKKvn40gPHhxx+vyZP2m7FV153oKVlwyUeGYSxsze2Bo9/t9kU20MlXqyQ
pF6+b8C6ed72Rru/B57eDOCyA5rAgpVqCj0KSdiQaYh5IDaSuBNdY2SFLfs7QgwIVHK3qIzhzpGY
SajIl7K7D48olvwCa4sYtTSC4uggMb0YeyEshAi3f4C1573CK6uMTQPLzJWjp21efkV7s8MVXhv4
nD1mEFYfC8PfTptpUcbaOQzUV5Ghb4v4gWz2iAkjiMjCU4g9T/Pg7upE/9ZH8IR0DoLMSyQveWKY
Q24uU0M1wRzde3wjLncWD0vCchQRkEnobDZSFSCjsxEMZQeDSBuMY/xiZW+MhwDIrhIQpn19/bjy
z1wQr39cxWpbEzDEGOXbibnpLAQnFIgMP58NNht3Wb1P9mgrkI8drcdziAVuzkTdvYJ3+4w/MQT0
/4VogRaTugulKxgq/eWNuYoWzm8RDv6EdU/kKWrar/0F37PCY9vNioi0HJ1weaDx0c3GqyZU173T
BveE5SlmBoGD/3Tqj1k+2gpY6U1Sm7+ZgjD3VKMyUS2IT6ergbnWtsO9wXfGd1V+YOWedRhhOb7Q
xZtlLUzJzzyWpHrZV1U7yt/1+hnxO3XNeiSOMftl0V4dgzXVIyeraLoDafXx8+YngYyBMTPrBrnP
N1+Z28ZikKM2LdELoJpXaYYC8e1kn8v2HebzJEoCQIAZMBFx1sUYr/p9FOwPdb6fK6dobeoe/mYG
eIhWf3LX9nQRDussxDehdY4tNBtBwwh3vTbUqE4aYR2Dcy3pWBrrf/M0lZR7ZxVrnqsDJKyNGL9K
YWMo2IW/GHqrAZt0KX0Pi5nX0+BOQBiUeqCOG7D+IOYAnnb6bfwHDuh7Q7c09P5KKYuqBr5g7/jU
d9ahguvdUPCvRMZULc/zgNIKIylr75/Rms+bvuzl2k7U6/HSJoTd8ja/e4YFvPvY6yiNIS4IGzUv
n3Erl6w6kqZ2IJTBTQSOQe79iIIxww2vrahyrT8BRLtRvK6NLeTq7FIN85KMv3l+STavYLpZ+y81
HB7VN+J913qAwEG8C/rOwaLA1a6h0z0Q93HFH0PNBfFChC2wimutoMXVh5zQseYzPd/3gUpyxEnN
Jr8Y4eqMQlnR7jXuDAycadH+EcZPgzzd9IUCO88TwQuWWce8VOm2iu2YStW6jEGsxmFBjKi10ID7
WqgY0epygjpsresZQuwmNgLCud8cnCTCmhbja+Xq798Jl3km4N1FlGF2S7aCCKybEvuJYJnGilXo
fEUjW9E0R3Q4wk6Xn5K0h+COURxJiX9Ts+YAvJ8qxgZ/HtAdJTDDk+cl9Bs8CIc4P8hO93Jn/Koo
eXTFN+y/xg6MWD0DdksG6BC6qqFt5KmPbkF2wzbr7qG+Jj6dxFCmgTcd8j1hOp2iAtsvuMRfCQ+8
y+POwaQCqDPccGXrzpYLwptci4fCBNySPIZqEmr2qjozsVCyPWsa3qRagFjz+VgXMkxqUlzFdSzd
OsPFHdfcdSvSsXI8wC6bes2EyuF8eotacRibVDDaCNn7yKqcS+vvEz5X/AWgcZyvPmhvLGZ5bjwR
n8ZMPIktRZfSZfWQDofGPb0+NDab4PdmIxD7C5tb/DkKRCKmaTxUsy4xfMTLMAGeUzk5hTD1tNOh
T40Vo0eyC982HrbAhx6UiyX/w7Ry9lUljQt9bYrBkaLmOlvB+tzj4eD1JtAaSlBtJvXpYKlzttgg
nBjLXExSDEp9xZ8SyoHcUnH7pxCgZvDVXHQooO0sfcBx/fp7tr2JophRZwLWm88XxTLJ25oVaOOx
RqyxilcN4YHEVMyfCi4xDmvGmNFM+vCrkAHmtj7hEJyrON826xgbrouSO3yfbTtswpgP32Jj8bmY
RiwkWNhvtxBO1EK/advxsTRGyaYRYVp3oT7qOI8tOpe8F8D2UUxj0F1NPz9WF0mpMb4GURs81vLV
k67MoF+ovNTJuMyEZ3LWkOiAkVz3GeVMSyzXvJ624fOLAMCyBCZ0jmkCYlyxzWeWTH5ytcShKlVh
ImdzooWvo53hwpEfCMsUfVisXgSFMXEqsBpE2X62Ast1dEbLdbuEZI+DSeQPJ/qQBNTWYARcKuuF
+wblr/4pFB83jPMbLActNXOFVqUXWFDxDexqVynxaJvD5M45wEoCROKZgd+BYE2Y8KpuVo+hDxyG
lQTnMWGctM/9jRYNCKryZJPyPaD1J8pmmrvaaDF6w7UwWPQKY8FMXo0Zw1+chM86K0dDOkcpPK4U
2r4BaiBAuyxYDMKS/+uf/qv0Musf978CBJPR7LKd89h0o4omNLURy07dC8IcYpLe5+mSjZ6+dtuM
n+Gl2PjugrYriZYHkK7CEj6t6xPkM3llGO4MiV/2l+PhLNscaafYmSlp6/L/iGq2uUk3at3Ipp0V
N1/IHoGPZ1jYHvsCIzi0x2ZJLfXNoTQxS2RbKWw3OgF/yez6U/LeMCPMSE1D22/tQ+3WGtG0lgO2
IaTLDt6I2ioGr4OlCzLMCqIR7mCnvdlt9jYfHO6oFgQMlG/mnYFHs6qNs3bMmDmyefYeuwtRBaeV
+9oJ1X4vDbxCIM0SzCEkzwMZ2OxYST6Ga+xt8PFY3PFPfVcgmWlzuCrFgkXX82oskRysCI2o5xgq
0jr+6O1m5RGonObGtnwWFYxb10VcHgFng7oqI/Vg/r6oKBjQgd28IgmjwiFKethpzy6sVQPtU5gC
zoVmTMjWkSCcPSFhs5s0A5E4lWlxtGTFayEDVN2opidO/uCazZLlHi6ZlNkEiod7p9EzEXO14rM2
iU8q4xg/EOqVwuhTiX/5cfFmo+ps7iDQU0lZexK/buRE08YGeYXcC3OWH9nqYUn5xlt/bjbMAU0x
CCTXWEvPEfxmhXXV39V8leEi4wBMxjOiog/yjFQwJmi+OMl9ay1uNEYp25x0myyaPPPkFCfgf8vP
baXucnpXi5JeIRalmyau/McmqY37+fp8GCLuP2hPWyUN/g3meGW8MBSAbUS57qYuuRZXwAihwrYM
5OoY/BG7AOCsd3P+jxJNcneWk/co8InkiidyLKUshv1oHwmvX5ZEEOaEdRnWOsu0GPsJ0T9fOVtV
zwlsGcdICujABMQqf6ztAQI8wbWOxzYn7fJ/NbFtJlQfv4nqqze9TzHIbRR8bqctgu1s6ypF8pkp
Cdu9HZcvP19xgWpdDEQHqGsnZhTVDhuLZFmy1IVcVICZmxeUknJg3Sb92HUY/Yr843jQdHtOcSbO
qk/bfwo8fs6GVE40ADFZDekRrTFCBlTkoyQ/u1/azVzrJB6g/t3owxw/ZOwFa2ErrCjMffas5OPL
jVZOEND0QstpMhpnh+VnjIl9LQjKzXl+/mvYLQyZlRrbolvfZ6D9ZU4zqIn7JYdRk7biqDlSUWB0
INQrdUubbOFvULCt4M6VFdE2e0twfmSmpBczrPwVaZP9NbpZYcP1rGHDIveX3bfBEjokPEa9mjQN
t5woU49oUTu/o8s19puuJjNAUWJcuBWTk5q8Eev4afUpO42SGpemKcoqeD8R1LAxWdrp/sq/W4XW
bozqNZNUkogL2iDPKe+fG3asl6TKXIFazZ+uEO15mbBtAQ1nE/x8dmbN8GhnFkFLBSvIlN5Pvi+a
vNRWMaHSEQD3eQAr6KzlbJXhfHSdPMG6SbA2yGiPNK6yS+vYnTEtNzXDDMR4fmQWTqD5xRmcoefB
hEaTH+CtE4YFMWPgmRXSPJ2doSMI1xgI/8vT5i4jBZjRizgodzgFdxxckJDsdsMDpZ7IPMZDfrhl
hkb+qsovqVGBDGOGfLCOQbz3CQ6pVLQPf44FML5GbURVR6H7X30T6VqfsTuQC5S9sOG2ejrdFSF+
Mz7NFA7kfc1vIFOE39tm1geBPd0yp1ZZfKZPlkQ1b0btQ6G/Yi/N2BOXWdHPBJGrq8vzWxTwTswJ
LBY23jHF6WFGX3rgBbORgNBufQMVGJWm/cghcV9T68xWPvp24NmvYHoqZsrV7lU7EEjljDo3OkhM
IEwLjILqOu6540+8Bc3HH7gts3sHCxaaKoKzWtJaM9CB7BG9KzfTDRGjUL7ngOMZNV6ZsJR+5/C2
e7gxQUQyKDK9SRoGMkHBY8jW0WMpSmCWu7r1uzIj1jl5ZzIH4Wh0JsFybtHyEK+dnMCEq4Sw5DBS
6YKeCa/5Cja0rpFKSDoYdWjmxhfmkLt8CgOv1jz0CgjUqDNeAvSmJ4G20/WNIcIVbCFkz2YPHPdM
3gZCYe1V9rL3n6a+4Mc3zcBGMbBz3au07aXD1GWXB7Zzd52W6LZylVv0LRdfXZEKdq4tsGPxBbTV
wTfjVZEqKn0+K+HP4u/TbL2Y2CssMSZ9wXh6m4okBMj2VPfTvbHoeU0Ilbd7mw4RqCT6p0zDbRIv
EZAzmjFLOOMk2cRU2/DO1A2a0o2QWA1JVJTJmUiOeKwlDAJBEmWx72ejexSBrkOk5pmjTkLa9T0N
pMB3pMXNyUCps+lUZn+YzAiOxHg63EuQxTJCTGaA2V0YYyHRaUUFuACkBVJzqK0gsv6/7hVrR4h2
pu+1odGJGehrXx1SxWkh7BHD4armYtoHtBAoMCJbFK1TB4/WBtKnLcvOoTojEEWBhmqFvXR9OmWa
47Tt4AkqHGsvgdBUdz7gQ2ux/jFbO8LJ+lM+mcTMoQoKcL3PcPg24X5DYQG+HpJl6lSaTNQcqyhL
gHL2t8JxNACMohq7UEKVXH+U8Tj/46dz8BaFCNLRULOITUPUFcX/jF8fKwyyCRAgjykaMTrcwoZZ
XJi8X8ZJu8ZGUVAMe3/ACpglS/Orj7mhMoVPf8nB8KP3vSrwIDBHpCLqVc9MoK4RVxGTh7OZSTPD
MiQGnvUsWRIEg7+T8aNgPbOuD28/MU1Mikh+ugeUMReTuTnV73WsuqO7KjuytDhoUEPetBeg2VAR
Vo/TpIBMimqTDq9qcSHmXROc0eDgnDsDKfHBESJucd0SKhtpCnMyfCvE3i02lR0IUcj6dQBzivZ/
Acg5O0dVeFdHzRZKV0H4AKVyDsskTXhz+/9g6jEH1Px+hxny6vKUBNK4VYSwOzbyoaIlfcsrlc+x
mXcPnL+S3287qAvEoYAzu7t29Ipltle+l7OcG8DRYw7FuUZsXuFz6B9ppWK6oMDOeV2QWoix/qau
dnGo/y1nLZsB5/TO/zyoYKujHKwAtYOUkaLs3vxyptBKK3E8n4aHOXwDxV0UbYuimKsxpdnRKcP4
lAOztT6qNlodcDvAE2j0fCwnLj4bRkq8AaOwNtWHtp7k6HgLbNa1oS+221RYGWbNMhrYWigYtKah
NcC2XxWUBVLP5LuKSdSJNlzI4NfFgBasCtZxxSLk1mZWg95UveJC4bY6xPyiSxERH4wyuMIhRAIQ
SybEztOiNocvGZk+2V+3W6FT38PI1v5In+HQA6K6kIhdygCVflqh3/2luO9MSxAHrdLJw2YyIE9j
qESeDo5RGLCJLad6uPrlDomHDs5sv28RTfUVV00BGzFIK3XfApHKkmzkgXbj1TY9ryJFmey7/s+9
+qSimkQTZZ6TTGIpjfa6j5ba1JPg4HqdLHd348wKylHLWdL62Q3SW+8FPhfVz3iF9A4O5CwZZkan
d3/t/tJCKE0YxekNtLbitrp65UYoUyOpvSawUmo52V2Z2QAbtLk4iitvTuhbqWlN0E9cHKFNmq66
IJZLdWc4u173zDPJlpJ5W7aYxnpGHDa0eg8QlhNgqhLI8ma/g/bBLl9y62gy6EgHA8aS/JLQBECY
jfyxHPUN6XNt7IMB/easwiVGTksDKyAc5xhajPoeVSgx+3iWDwd1aSJEY6covBBQYMxgZ9Edk1xQ
wYXoP34uwKYJXkgTS/TBLjNv/NGXhmFlI+1lwRLUQnBmVMkoNxuwzuuDtcSlFgnGZ5dTc7FTe0H9
fjGfoh1FpzHUdFHeoPWUWg71kCdTszecz6vz17Q8SbZyzBGp56vpO90pcsLoLzy8XnC84F9ul4nN
JpidhULHe0LjNgC5op4hiwMm6ZXqs27SgNq7pabNQJS7yZA8pBX/SeDhZZL9rwEQZ890w9D0pWMo
jZhttPL4zS1R8eLp9PxjSwr1YnAASUbeRsUxyjg+fu95Da7l2LdRwRXq8rwQA8bvYOvWi0gGajGB
qilQhmjpQfUPA9OlbeM5+XNI1Y/0/N4ibYBJ8+xdSYXPLeiQSIhgtTK4dUEJm4yRsh5wEwhjQRLi
m86aYOr5BwvCOhX+sL8P/BsnBOLx3VIYu/h0iJf3pxvDI7aEMYHJuVty5jJtEAp98IDxiCpfBIwQ
/31Z//6onxGbniwAlbiLmDMj7KA399P3wikw2GrYg8/MDV+vMy3lcrRPFA+6O8qRhzwXwuEwWYjB
BHRDdEKpKtvENeinpNdIJFjToOLwXiRaOakYFWM9wH4EshkRLKRE2jHiJYwuOGyfvWVaI7D2BtFN
1fBV1txY06ILSikXuK5fLHmByUt0yCmWHU2QAFwVss2copu8rZdKXdz/738SaqGN73ylv4JF/1/4
3pXbXuzzkpE061dH1CZLT02qbeYnN1Av/oTC0anGo6TWxMzzl+7fHI56rxL5exzz2l++MuJzNNne
3lXV5LJHfLrCAdvGj8/N+UFCJr7/mnEmdFo56kDgX6q5+HYAJKRdQa12/34a/TiGwgEgdUBeISsO
PVNZNPzC1/8JZWcB0FYqI3XDKRJ9dU8ldgQ3z8+e42CnPUY5yAtcCF1EsRigXAtdMHvg0jdT0NGw
xXDxWtji+PqTBLjkWMODiGBauAAfyjfAzhacGl8it2wDlBbMRduAg+22TZO4vdpTWM2PF5PDQX0T
gjydDd/r0SRKio1yS18y2GJRuUUN2NIVJ8jEVHVnKZ9AWZpex9VVRHcNy0xoLWtF/yXu7UN1SToA
ZgSTr/4EA+Oj4Qy3gHREySLP6UPaScOeogmx9RLveenFRMWhhuf7OtBZSXdRU7yRhgeRwPfhjmk/
1xFruxVETOlhh95AzqbrxO7dFHsy0Qyvk2YrXnyqVygXdRMDVFGnNlsev5OmdE7LKJ97tuAHip+4
7d7LW4rA/FQe9dcy3CvXVo4I/x7LDluIc5NC/xcKKf3+MVulItJgIKBYwksKexRL3xjzgYyLvX/K
A1ndQcDjJ1q6LnWHKayq1SCXkw0l6UBlYxdo4hsctuGpTQQyU9VZ5EaVCzDl9//6B4hzJj36DfW4
9y7x8k9QSztdGNzqgy0vzCECKQMq/uOChMSAhvbM+WU4mqGeCN+6TYsJOSWjGeAQsyFKMS033OO8
mW7DLwa6uKHrcwnpbfj+WJixaxYsjzj/T1nbOGDkl+yIZ8M3mkDsRzcazDGJZrJx67XINCnIsMLS
cyLOw280DhZeRncddzset3MCNvwDzyxhD10g/TLSdFViFQxole2Kq/5f0wHRL9kuZBUAEmgerO08
ALmfHd8UE2Y6vfT4kKOW49N/p41+bGMafgbUPHqTvHFGtSYRaVC84I1lPGSaz9FlA+6wjIHeuRgK
AJ1YTHWMsupBSRHPqDiBVOCjt9oDIyCN0YwCO8l5dkmHb3wBr88yBSApDzBbN0Vea8cBGjD+Ruzp
m9uZ59v/bDgLpOHcUxDgXVQdlow/evPUKSfd4aw4XFji0CXzZZ5rj4yTr4h4sCTxCi3lChbYDSJJ
HBudK1R4AjR4CpxvziuFzp/hpY6lBSLDYeMjcd9Ns3zpQgJJL7uWDP6VQ3C+0iV580Kjpg9SBbEd
aayl1u6nFCLUwhayXoW03L7vhQAqyTjFB/rnvR71c1dzh0eamyZzet960kPVXTwXt7jS2FoYIkfm
4ddOFgWM04C2m2ovIes6qZX0VduweN/w010yNwF9zPrtSbtNsEqSFF+Pum1goXVQ1mejYvlmN839
E6fy0n/j1sL/o+wqW5drdGDV6Y3zW1XO9Etc/9ZN1ZqyuFjqhDzX8kx8gm9aPBMNQtcedg8Xy9m4
qlMcT/zdGUbFEUC1lNycPjwZj4tfVDTm1PY5bFg1Q2LIjESosfSuyrswRfJ5LDjzPCZS5IjQI4up
X0YkZ+dsQarl3HwqtnClr7jJmeZc76xZNGhXbv1PeO/YbLxyDlPR//QXEMPXkto4wausPW2y7bWf
C9Gjfl4LqE1NJIr+dwEojrCIWklJYePq35UJl0JgbOX9+fm6I/WivzfqcCqiaHGcASTnXlQ+5SJB
Ch7xAGNEnS17CqeqDVo2kBBbmChq9O7nJ8fk4aV/mLCTWmorwNg0ayjQbwHjqTmakcpIeorBP/g1
KnctZ5hKXmioIFDXzuneT9JEYUf53WJAMJzkQRJk2amb2gQDiG6Cr57QjBU6xGSxxc4ugYswIyCb
lbEzQEG1jUN72vIvSh54jg0CZ/PRcgaaNa9iC0qw4x4MdeCkUDB8jcKUcc3622BfHAHjDFz+D3sI
e9XPPd23579nL3GBi2eMH5pQS0xOmjzyNcoYU4QJ7VZ1OHiSL87xAuzQic/k9A7i4vWk3pt5erzr
i3yTInhRgD1DfgDEXA70mL58VpdYOdWWQ5Tr6mw5mXwv9kQMboqQoH/xmvpwL6AHKTiF8au7bTAx
tguCvEo7ejzZdGaMvHXUbiFHj3YWWl6ymMBaX7myKjIYeIxipi0qui5/eXu3p7uO3Ri8/YcYYlJW
0Pq8Awp50pVNmz5KOpOQBW+v3jtquf+Sh32uP9MKR9MwauTNGgio1v+6u3et/H29ZvSJaBJm0AzB
FsjXVZ0jEM7ANQqXvwOTmLgWZVSPVGkyZYL5fOWT5lnI74m0pJR09f5Lu48N6r/n01VVrtZUnkwF
LK6a89LwZv/9yoEAj7rK150/T3etDzC9ZuLGXEBUCh9lfDGRzNAP9ApCXrrRUo7mg50liiCIhcuI
nFfQ6MukYxRKYzH8zaPKLkL+P7PuMBfcrFrQE0mB8045xpDQbXmvS6LXyJRuaL9/7bK99UN34udz
caVColDU58Yr5kEFbIJ8XDccva1WcXupNBRHvCMinF4ujYsWIGNyOmR8sruJDRajYtkQojEoyLYe
iT0Gf/lv0GAXr4XO53dSUa+sm7WnrCSpKkq77dZgA/3fH8BHFTPHyaCRG1WfVGHjy56CUGd75I9H
eui7Z4sLzQs9qHn58dZmj71hHmYSdP/BN0VzG6zQW0ZjBMT64zCsj1YbWawT5NRRZsUSjGy6V01t
svJ7OoPmWgT1S5IouKXKNRWsnW8UJiZAqKO3ngSg5wXr+ci9AZGohYGfjokipjKx6GzGACtvKMjx
oZYHO5dN1ojVlsIJpWD+2KJhBRuWrf1hS4TpxIVNvy4kJnPnbTfaVvjG18NriLHtpzW8Y6A/MPRv
tOc37yapx0tIbegWExxODIE9uTfQPQa3Htb7c6AJAPzhfC3ytCPaisbFbF1xd+RhwSVpFVqmdLca
aPHoZfU+3eW4tYvODDdFiX779OLVkNpdTWlE8aVULofPAtCf9/CXt72TL4RAMCpCEU/dHBB64+rv
d2AkE+Zi8mCnTdbZ5iwI+wDj7ttEd3P5rU7hB/gHqHS8BjPcVmvMawUwUXD463RcL4mF4ar7CE+X
eU6QHejnPSaEL7Ndw2WaTXN/l/XtOViPKqD65/zMD4dHxrYeGHhxY6TZFGg+3miTQgO6pfccfpr2
ZEpt3eUap4XtPGOTLO7QPF92EQj3XAhSfddXJsco5tSnhmGcS2X3YnpJ0Kktp3fH//M9kvMTfLrf
H3TDxrWNnQMXHXlDed6bEYmOYgMJFnvTNRCqE1pYfvVuBUqG9TW/SYM/B0SfIm5wb7Q8bWglCJS/
BWNLQoOIEt94kXWNzvMbG+q3Lqn9LICc/9o2f5FZ2IG5Ow0NICOoLQlM5koAFjnhv18UoeOhq8rs
lLJ2+6EhE7vAenv2/5PSPPLxXULvRNnRpwU/8gFMJZqNJNRbVA3CnmE/AJrm4fbHOfW9ooGt6D/x
7JbI6gxyjocIAkmJf/aOX/05MiMfHAhDA0iGo1KNbmpAZL+qjd88KpGDyYbxswruMotRzjLDVJTb
eQkZn1oTMcLKL5PPxRZcSLnDhqwN+kpegR4AQdpi+BLCBh6B946KMFzPS5qHS0X7tV1w9YeRUj0b
JzrEsa2fwtMLIr50Uh4jghENnl0Mpeme2uWryWB1r8RPd9hWAToZ91UMFNBpUN+MLMKbKJ2fXkOe
hvzlKeHEEF8pPhWSF6Kc25PeZ0Cwd9UFS+hV2Vhi7ouLYC8EH31X7gItONukkuU3eB2nZr9zNlT7
mKBrezeLTWI/e3XhBA/wkLb5cTs7rAG8IWk8L+xBVM5memi0fBSagpOoMYNs+Y7euXlHe8UrgJ49
eJwgdMwES3CbkrnbbN7L/+HkVzNFdEGUJ9AnDEb2SpsTirngMSeXm71qtCiK2AbFamm9S0wDftuy
JQJhIhfsyHHZcg9/BeMSJLjW3+RM2uXR0DRHPvNLNLqQauNlc9NDaglpLqNzypNpME55suk0XYkh
YiSieisqSii4tezrAnw4ba9qqi/Kq3QBDqGXS6t6e0ARaAOUvwz4+eyHfVlr+dSZgHuF9KEek+ZU
nqNc6JDLlwbt1Aby4CNkoDhK891CIVsbegB1syAFmTY3UCdF0q3faJo7UHjbjuMW81Q2cVz+l37+
BVKAr0imiV8r4YuylYK1fkmbS17SsO5h/h3yK6WhyAHCDd/RbA4oyh2eWxGwy5m4vX+MF353IxVo
bfwiXM5p5IqhJZB9YtwUh0xSdyErruJmCUk2ljRtl4zoExP7TYa0z/suMOXD7Yr2pu3ZVHoOMZkf
RRS65R+9++k1bkWNwbPxKV6CWFIfZHNKLlKIAt7QWIyRg7Y62wHloh5+qeqgv0i8CEdSvPc5AXFr
YbS/H8xKwDIelT+x3Lz9EAEuw4v/MkrSk23zDSlprBwAHl8mE7+okZPx1zeqTMy2RT//8PjmC+bv
hEmJHp7Ay2jmUrCiXB7UuUZhVzXuPeIXPLMcBLCQB8CCIKAOPPdtku1q6ber74jyoYrXoMIgvf0A
nsUJPHqbSPDFog23DBBPQK7V5Q0cI5h2WosGo8aIkT2ek+/nM6ysFKRIA1M+uvEt7F7ZtN2uoxgk
mTFNfWApJ1OF8yAhy8h0HzfioGz7bNwBSZGJoYv7++0O6g0aWM30RDQI09NLiKgsUe1njjpAtFK5
PTvAHRWOonFdJNc/2rUfXsJxkTnQbzSa+8v0s9k2/YttAL+ar+217yADiyorEXVeJMRn7ZgHLOOi
x2C569FEz54T9W0HsYqx1XjHeDfYPwgJtubD2LWmWBXKsdcT5HKABAJo/PHDBisToIZDcMYB2SG/
FoOA9Xk7koXtDdcro0WyGH6z5KHseCRFHcBdkoIp1jXdMTmUme4KHTs06JgDGYCnFXhev0DeLq3N
qwSlpjfR0XCHYhNP+WhN3HV2KQAA5SjU942rlDxy5DRb724yrLcQqXWUN33aUnjwpSCPmHI5hVat
8EJ0E6rx7KYRVXdZuBEBzP+t23lTq73w2qLDdBZRmGYo/E8q3RM1TbzzeAycUGwT8IZEKeICyAjn
RBWoxKRh08EsQ4Mdfxa3tXTaZ2uXbN1wdWTqXoAnmhaRQeuu5P2U/L3z7AruNOKIS7XdkZe9V6IZ
WNvSE+0zEde4Fo4+p0vI9+4Mp5YOEcWXggY+hznPjvxmHE0rW0N+2BVXoXercRDnSzbVNOMdpAYM
P6TDC4/QNf7DoHerbgotsfrYzt9FjHJ/ILBx60plY1iDdjBazunIHP4EbgCWwJhDC2I1g02tIySU
FlcEdo5eT2TggSek8tSbCfc2rPmgle4i6A0sqCWSW2mAG44+FTXl7vJlWtA8gZXUYj/wSTysEn9d
/A7KuoxbMIJ3zDlOX0D6RJM1iq+tdbX9Z3ciqOr7vtS4oEsX1/yoGYTey4Lp/Dj6S8vUQ6dlmWj6
p5OI5DR+D4n3ucTN9kqLg8hmVOTo1egapjBpDC0mCPxBq/+8pziO2zSHnoM2N1+nH6GLSkjdr/Nt
ofAEG7VUuAtmCa6cbFw/aqbibDMNCZNmuTabaNwdGApIkdat4ZnVLmouFtd/rZkCKF+GHETeF1Ol
MuG/P5mOFPQ/wfGp8cg1zi/yX+DxNefwe4l7WwS2OAIkOm4bwFJyf0vRpcld9fkhClwXTXYrAcaQ
aZglpwocrznI/7di3Frp421PRYvAnc97J9nVBOhiLbVjEE8vQ+nsEqdUUs0/AVb5Ay5cMRERc5+n
GkbZxVeYtuZw0fkRZawI85mIPegFEsY7uqi/WR6PHmAVDfu/ZacRoX/k6Ci/eUUH3oL2aeMBam86
gexiCIFtHS5TzhO/7LD6FikhPgfqpgAmg/VhHtJpXlluEFXoEnZYKhZmebVu04e8HwAZo7lLWEXo
CsaULx4gLf4QaUiSQraRqkZc2fVrPMLd+1CMAMHMomWmsU9BjcIf1aal2+cq/KFs4GRDl5KJRBOq
HnZIEtTAD01Maz0U4TIKh+lpZtmH4YSV3p3rJs0GBrImEaUdiBzC+eOPJpD1VqAl0QoE57wk3byw
XOqwuaiC1PWp3xxr+om2jw3eJTDB8jpXLq12/FPIi5lUjMnolOPcwLNwg2l10n3PfQJFNnfQOwE8
Qs1RV/EUowzbLGfDnzNpjclOjfvM1KQYxuztPnoGTS3/DV9G+SdbHYHPdDhNYWj+S59i45CRPtCB
KvgKAhwZQ/TIwqwB3yLyQ1RdjWPr/uD6xSebMPPstTDreatr9u8V+hLMUULJfuhybaTClo67QUsB
RR+WnfvdZolJzh3fUxEtuCtvIwOiaVA6qZ6/CMViWvh5U1BlhwQqgfLS/ETddRP41rEZBLPZOR7r
2J2B5xVDLThc09H+OhGrHH7WF4wCu7r0+DdOyCzRFLLYU7PJVDOGOt21Mxetkee7fDa1KsmRKkYI
gqL7WWQW6G5deBE+hTdy660Xt4xwjcDu7z8BB/Ue+G83pjGkpEuW/FDB69fNKLQdeZYcBGZUSS/J
tUKonTfPRx0vX1syK2jfRX+biEKG9kPJzcUSE+XsDvWhnmXW+VYq9dB2X4fWiAswjMvgW5NCQaPi
M7f0FI3I1f+l16oJD+VCjMPIvsw8HPy4LW/+w5hW1I9GfKS+TMTqJPvnww5Uz9YRgeX4Q6/JiFuo
lVWuIKE9x8F1Uqj6JRccG1SwjDO6/xrCt2TLmlTzrgg4zrx5rSVnZGpgVwQMW1vWcnhvmZguVH1o
dM1qiTF4K9S9X5DZrwb9Tv+fzSQ9MXl0vbaeZmNl9ioDLHFiraP8pEWcWZq2Kw/FDdrGkXsjpiaY
CFhs6GBC2iSFnjdzXgGBaXzhwKutxnzdQwHRz1sgf9XvNbcigGEodte/IzOBmfq0xUHKt5dCtZ/x
tQKf/VddwM6ZQbDtc4yQn2oyrxWP5+OVfa7aFnCKvQp0pYBfR0ZKVr47sw/X0Q6famLgsRVC2Gcd
lLYVWRBjLiB9vYbPWfrNTNBjR1Lc4BE/IIIYeSHFVY92yggpeI75aXYxGH5C6KxEQMhWl5ri++pQ
ZLcyzWKu3VAnDEVz92kyToYDNtODN/TW6w2Cc+SZ9/C1xY77V3F/8zTSlo6YAqlAyEmbW+rb3rdD
WbYeJlhCb1oTN9vB+zprawR4ekgwsA9ldtfg9bk3KJusV9diJGgCfDV+qMigFplQrjOG60xkgm7i
Th3jyHaLL1wcjCQF/aORAtXv8MYTd+d1TFkyh4CdgIjAKgCLQsH+2+PqSSuBJDzkwQWG7brpJYRZ
T00jbHYYazETWQ2L+9sDA9GcxweOgSupFLPEoY3G9UXktc5IWbVsxL+2NpiCREFY0XS6nLrBlA2s
4NAUYo4kLjlOY4/yohsDNpZqaqEbqJPfrAG8oK7KnfmVuI7kVKJQmD85HmsvLbI1pxl0DseZ+qbx
6m2KHuvPuTstOaXP0FxpkmuMKJtkSVK8OqIVj9Wscb8rwBARP1swVBeOYulglCjgkc/goed5tzI6
yJKw2ewsxgicwsC5UR7TIkY8TnPna+VMqkJOpwpAUF0SaZZsfDP8TjPrRD3WxHQZ7eu5yaJlA4bu
hulMyIeAsdcP9Tq3OXEIZkgZyvIkPsmfJkKXp08d2RFiSBXFzULPouc0EZd9mEEdp8ChgEnxOD81
Atc5hXBctbiKh6XuRn/8SF+3ccT0hjrXFHZ7ZO8KPtLbI1DrmXU2ijUNcdfbndE9fGkhdUTvECQW
Mq5/j476yhrvMIVVgmSX4KNMMF3imyXZgmEK/ySGDcmw3t8DFtqmVUDZb77Ds0ZG3RcjBpf3BqBh
iVoQ6wmI6MqzMnEi3ezKnlm+Cw3RMzDOkUB6mkalRa8v6v2e54333GUgX4qks7WILYwcV8r3ZM8i
/tvYN4j9PsbjNke0gVv+yEpOuR4s447Z4YyWiYZc4hqt3/tCy3A1hRW1YQhU6G7XCjsNiI4rwr8E
7BuvZuXxYBV/sP1buWe3BoreCmRCVR+GZMAwvNiXgU00qYv5bNcVJ3irXCp8KMvRrLWjf6KJGRyT
yJUkEGtqq7FhKFXCWuCmhAYNly0GDDussqbDEPb2xo7kWZAnPrciyIi5bZjBAcUN4lmrNHxikc7v
762/LY0O+kgKnOFAtZB6jWBnSFlvhdLnGpQkiOkDOrQ3Grx0L6jh5TNv2aiW5SLOo0oiSibdIpUF
JqgDYsaH7/0kPsE1JZ8dCouhyPPp+b4YFKm0ySjrPPop8DPvrADpLeLtQHp6u4jlnoJPStX2yYfa
0mTqjf0iuM0osubV5/xjSvtBZJn2C+8nTR953GWA09wqg83BqigpP4OgagF4eNrqDS4k5AgAPxlz
e1to1git0sLqpxqos0FDdXMKpU/kW1PP8rJvCPlHyDM3/FMInbKpLHew/1XL1Q8gq+WKZEHhPktu
4ddhcxLzA4fuDMKYvAfrtyb2sLD0m0kbVBqfIxO9RuWxLbRRuwdW6NRArIFXtaTBJpozBSuOZLgK
fJwAIJ0cPT4EW15KRWQD3iRO88DHGRh/iQM4hhk6XOqgB59HjSK6HgwA0NWUu47wtGY1/0j6MtLx
qxhmfTMX5hfHZejsD+3swW609y60mQfI4Mfk1IHmR9UQmKuufEhVm8tVu3U3i85GMPQjCvMkszBQ
068zovOTrgTdnODinstjG/qzw2BETyMaQDkZ4smnPQ5oOnVTJggrfcF0t82gJuempuVG9UkCJXdY
yt01f1wLJwC3wK5Mc4+hWmu7a2LSVP1Ga0nyvNg9PiePEYqCT90THiWvBl5Rze6ZH8l40BMAF3T6
JNg4090AgBQWAgL6qoGzaMZDcOSFgc5WAxXMPTB5D/514b7c+/7oKN6GOWgkOd7VND7uyGkPlT60
3ypLMfyfosGEwoFrYPdrjVSbk6jQ+2UsQwLsvOoEF1KE6FhbR5M0wlNITy/p/rHS7lLDr8+LtUrk
tJmWIORnteOErZ5WD2ULuLsBZx+vlSxcOdBiEmLt98oSyb1rrlEFr0osQBZ3/lurakP2+4Kbnit+
KP90KUweEGCG6+8Gx5FBKyWJuh000cVuIubunwgu768eW9DE3IY7JwTApdaXSsDg2rioAPT9cZVr
u5KzxrTXQopP16uxIeM1GgTGPM12Q+0jgT1DMwKYWE+gclD4XGks7fAFmH6H7lowK8znpCfZR7LI
FkvBvjFXzRaZE/4OH9iRYmGOYc+CtFS8rFgukJZjd9xvPGwMxKMJJf0k/chFIwyJpRHWT8EWuB+1
igokeKVnB3SbbvVFqHCryFRJFpOg2eCpzidhdaDYROTioeFS0FoNptdOzMtcU4wcmacGTi9F5ulm
+dwGEGOXXttFXZeRbDBd46jpeoITykZkHhy3wCD7ewcWYGT31MbsbGgpK+1IzC6Lz/AYYysSCuY+
xSo8kjQeFDCqGpOHxDVSC3rZpFs3KXygq8ivNj8JzPV9fogHIPrQXvccZw4Z/BS5HjNY7d943IfB
HCLZtucjDoQ9oNYCjtRFcz+XJ7h1kxmUlW1ftpWdfpkrJag9ldE9v4P4Um1df1tGeCg3p7rOxglx
Bu7rMiKwfYC1DOG6753BU3STQNCRPpuzkCPOUdgy+mQT2/e23DfALORs1icbTSj/4eMV0aFyGkQY
QMZS09eYD4jCrMdoMjBFUy4yOLwUyO+HJCyyOGRxPMPoeuCaXszGc0l0mGZI1u3/kqCCs4QmPgG9
WxRHRX2tkuNRSDcnRoV8FbU5+YArFWriAXgWUX0/o3Wl5KulNbMVzm/k7+LzsOSdaOfCXOVL3tHD
JJOCXUATj2hRTSpAMyPhegE+O7l8ZITU1DRfelrIo08eQTqcKStSdTtFCmCeGuLFjskv+YEHWbtW
0PKYHPvcYmqILteuLDUJ0d576Hsfk+CrHiJg3JMU93A8bLodSv57o1RW3Mg+X/0sWJRQKb15DnMU
+ai2xMGtxbk8nWQl03MCCitnNJjF3xdyHD338nt0KPMhhFqdWabjS2diBMzsUQfjeoQctE++SAaG
K98FF1LWJPT1HXwDjhIK1F22DRffX02CM+Z//zapPVqBpxIOa6tNEGZ+e1A2CpYbD2jsgFDBlNj9
hPrpVHZ+d1YbPMbvBhI+VCK10HoKpP0NoXXf0353Nj7UEToL8974MrVJX0TR0iisEEnXt8vTR21x
0Zr6YleSPpzBALVauS2K4Wdoot5rJNbhOScQUV3OS7B+j6QmdfpQARC8pgKHPy6QrnTnPL6kvdlI
hxXizZKvYU/uFn0stT6HmV7oIlTno+sWnXj046z3LdEABhjQ9nNM+Uud6Cqwe0KMHlFqrdxUoXHV
94lzrTzqr/9D2Xq9eBtCe0C1aFbStK38VmA7VTSCzrJkECKuO+E0P9jtMf3fV0gsmXOeU9qvO2no
ADWexPXSoJ5b6tgqYkWnn6VU0llHw2cUeg1oPepHt45cBSxLikyRZORLCao7CLPcPqKSL47boLNA
+WIPB/+f1Hw0Gpn96XbUvO77H35kRXrqlCMrrUIZQtJ7x68GljgEVR3WaNNAT4J9vHixgJRuGdi8
jbVMSJL8PuzdohDX5N/FzQE7kCI2StpjzPjBfRgp9Fk581XSiRgNJ7LSaxmqFnjmjGA28kgOVnky
th3VaP0UVNCn+3LK0SB/V5IlKY7snO/OexwUYcfF32nji9PHeP8QR4mtegvZciyLA3p1/BWJLHlE
ZLoBrEmovU6GpbQ3GTEBaRxC0DiSDSRrXtYOpMv6a1g4UejeyX2+9q4fNqgC8MZ4TYu+xA9nNXgr
/5zErU9Bvj2CjU7lkXfZ8DQsOZXO/TU6fKK4c1BCV96l3S1LI6IS1STFFRlfSjADxqj6Ar/DYIzU
hRhmF7t/bwYcuOIZUkbmXCiFqNheqHBGP2hmFYk3zNHrI3b6rp/Xjgs3p7PhVRTYd5Rtmel9KDK4
QTB1GKW6GtJePStqT5nuYzyX4i8BQEAHB0nZgAN/OX0oI0SN+amsAlf7Odo364B1L3UgAF90KTh/
XW7ybXruVWxW73CMHgC+rNf5pdk+/b36p80RHlrtFR+2rEJVabhkOboARMUIbimuJ9vxLkiNqc5g
XhbXAioM6G1jfFUoU7AKPqOksM/DLypPvQWQ+D5N5m+ML1JP0bUpEA1gZPBVnT64MEqDDM1BIPRV
y1fvs8CdtrRvQUi5RF9r6LV1PcYcIaWG0eAJPpeYRdVsG+ygcFv4LXhCYZIlV6MQtzwsYcWH5C+c
PtgdTSQuJxVLQG+OtUTKB7Jqm4ANBTHdFdpnuAW1RBjriE9HwK+qwjxS5Xkvn5gjS3iafaY+8zhJ
FFXHGZ4qydZNGM4++sKY4Cy60mKNaDLabNQ9dup331hBTQ9U08m3spj1AI8A2C3bO47vC3hWeEH8
CXxLDCxRp9LNcF53rgfdSSRnlGPxyDYg4CXBqv/7a0ABzEbzEEV6uV+5yY4Uqff3v+UUWzsjdh+H
uZQGEUCaLf7SnvxI2HPRmZekBfUZ1e/rqts/DgVeh05Rc6xc1MwSVcDra3gqHkb1EFKJvryKOVcA
OLvjy7Dgln6Wem9xZfjLeE1wl543TOZZ4xbjet7yEpba2W4BJySRyL5wQMAn8cNxLKfFe2wPudjL
jyIbnHqH13VOiJI+oiyE86AAaT3cV0LqVLaCJm67KOVH7qQ4oiZnEF6tb5lReICbjiXLLY/R2asw
XVZadYQ197S9PnAYiduVsS8MadfoX2fDMOtKlfM7thAu65ROcG2v3hDlrW84jpcNjnzTEzeemPqV
ARyvXKx1jOulQulSz14VzW02WXvH7GIhoHD+KwlldwXT6kRX0mnOvxoKRY9dBLIMx6c3AKZ3ZbX0
BP67VxCSVnVJw0uRoDsEDpF30SkHUssLQp+y51kIGcwmPQO6VzlttMX4XOdPgug3vQ5j3b4cjZ9n
zB+PlUm5csQ5frypcJkPdUI+HOJPg+vwxdNbTbO/x2ZAKDh8ViNm+ON6bgUNxuDL5CjSUYPLFAwz
cFlc8OtntPthMCWUWYLEph37f3ThvJQsS1afwSdNdi2KYTM37gKpxrWs3WUi0L6hwwAcvNqRjaVS
7atYkgaWV/Orz576cdEhGuTfAsDLq8eX2gorMaZQgRNO3jTuV9/80gYSV0ZTbhWqQkHtl4GM4Fme
Jjes1aj3+rXBAi8yz7sYMQV98xAmWfAxtFn2Tsw6YH3DmbVhLKNE4g90hkAQcd4EFrlrzjyRd7fI
PNfg8O8VZMnDRQb7leuF/+9GZqmsfCoAUNFqauBOYSQY6uCWBhZHRL5lKxt0S9KV0JN5AykpTOwU
SrdgRixgn3qa4ZLkHuXYdbhFAuX7hWMmceguNM3hyaCW513dTBpg9BgsXOpyXK+VwdnI6DGSVRSX
Sdc0vkSUEUnH28Gxg1Tk5FFhTiDbZsv0IJBs92JkpOlf1NgIBck8+VJQgb1AR8KiWLzQ8c2K7UuE
VmSkBPtlGgGhM9/le4Nl2oaX3rwy0Sg6BPt0SNuquwH2MKtxKhR1nb9PKQD8PZmfylA/g/m+DZX9
Fjeol0D+8lV6ZHCZ9tWzhjFwBXsgaJhAqO5Xqwd6PAel0sBkiT6Q19MYCMQOP98s6eY3RD06tjXd
bGLHqXcNafF9ZGXLwnQEwt0tfrbSmNHpEkyhdMvGOcK1sqmpJnoP+RtNx11JCtDzxM2OFbUOSA6U
R7fqKqFuuAdGNIKdyX+kHnmG8+ZBw1Va/D/Ji9hREr3S/Gs7ZM0h9V95SN7KFR/z42PrmKyWNjKg
WEdifB+BNYK5dliFa+gklPy/ZrT6AUrltQku6iwVXaBnr720if7GGPZAPMv8OALWPzXfgKb0IaOn
unCqbje9zYSNIMznxJdsOaVo8Ipdez/j5KU+pp0jvBhMFNxdQ99cqvDu7J0KeE4AmZLVWCshDXvX
gvgEdZsK1P3kXaQKeGpdRNPhmdGrjvzTET9ekIvnIaAE9uu1eLLNnPssO3X+7S0dqHMEhShwVHd4
gDyysUK+ZMWH4zHyRaFeoqX/pAFe/keOCkVbVAMOWs6+Tptw6qor8ZoGmc5VL6j+kRvPrJQEgYVb
DUYM1sNKUini5Guq58U8M/HZsZvlfcrzf9yUebrCItFexgtkbpitvuOvaAQfAKDExqZEozMLQS+u
vjAlAGEfwM7y86Ab3yQOzPtXiaqiP/vv9zgEQwKA9pToaX+TiKZzkGklw5Ws4OpSXaDWQuOms8jN
b9v9Xc6aopkdpDMNE8oEbqsgEJB1VTuAXz4cqEvmBVYsMYJ33Pt4Yvtx9wvbaxiQvGlXfji6Hao6
/biTbL4iATrQqePAlR5Q+ajtW58xIccAHinRjGxrOPtJCWa6KQQAx9J1C9zUjVUu7WxiXmdHE15T
CBJZugUup4n6Cfn5NzuJKh4MajqOY7LPOAtncmCJs3o/ebfxe08fCs/GZx9565Qx7Yf0Yw2HJ6Ht
Q1IyhzLbD0i2I1/4Md9gB6EI8LloDIIPzOa1kS4B9AZpdGeC4gIEmqSCxZkZxhnrmGza/JksbyC8
ORPpKK3Y7sIVOQMxrEq3kQVUZz9uCtKjaS70xh983KkrhzTIkR8huTeJgMGS6/TcPrQTX1EbMjFj
Fa4q//C7NayLaTAb/Nx1n/zRGQexUpQ+8PDIpItBA2Lklk96mkN4o1bbsTI/SyFkMNf/prYDoKVe
tQlSnF4FjfGo0jeqG6fg5zdD7slALjNCYXxA6OU/IIoRs3XnssuJ26pIb372sqREorT7U7wID1v+
PsRE9l+8Sz+CNmyUxHbIErYUcB83DDVY+mD6ull9uOrkojYh4s9H3YAPEEz1ZjswWeZQyzZK18Oq
Y4VqXQtPTVkbfIiI4ewP6g6Ger/jiipezxCxR2EL2pqzsNQTq/rvGUtUQcT6DZMMggQbaHe9exEh
YqSjEYIli5zY0S7adbN/gr131/Nqg2IZLdk+Ii+NJd0bWdfMLmPUADVZmeNY0xQuecLkcwdMC3nu
7OiVbOeRKSqPx9Hf4ztx3SCvjH/h3bJzw/LODaXcKVQdYzfGYxOxkuifgFmN1JkcHobDIiSxwTNc
udZl2uDSfZEtwY7Yoj9MMWDFvytR28+U1f3JHjjFNS1DWmRrP5Alr3okjSHnB23KSRh+phO0XCl3
e1gE/MHR9GunbTfP/E1G6WiI68waJNGC2aUW3O1YORg7RSKmewW42diyobO7zro5cIfUB9GWo6o8
C0mY6Dm2YPyhGt27Ddt8B5m3DXdKQ0d7YyOCqyAsFcLieIiAn/f2s6fq8tgveUh4xvDgxUV2N1wZ
kRq777uKzbdNTEviT/9rqFoXdH81xlEt3CbC9SD8hdyZ6sOdKESn3h6KYVqzLpVu4KN/V/Ku93qC
kmD3s+SujQag/7TSw7hDdpgEBW3wlvdxSlyBlkyoU2H5LpnQLeBjQlYrlq4NURDibEnyh4c84Hcu
pxnPbN5tJqCPFMVWD/qN21U/uuwuoXN4GXXkAuJrcduUjMZameYH0YepkTz7a4cb5o3WLptJBW33
V/HRMVIswP4KyMrf7H1wlsnpHjqWl2FeeJngIA6jzbJc/DCtNkM3No1TtUBeJprLkWng6uHbRxGf
bbl/djueg7xAPaRO2srLtDbHOa8hxT+WrfBREmLmo3SvWpNK7mEoEDbUXLZBnQHJHAMpnZ+WAbnK
4HbTFIXLeJNq3RN5p7QTJ+BrLmSk6UyEb1L/Rmy87jJorhwU4jydS74XYnRB3l7Kf9cM1Yw/N/IZ
AD/8g3j68OmE5b9sfXXYorg5DM3myW0YVL63UQShbClpaQqjIXcnEnj07QzA5Ndq3siwbcXd7FaM
s9cCoYxJY5RMIFxosL5NUntSnCwQooqMun22s7ASrk5OPZSxNaADVlzqNOHMV4DCZ9HgQfVFNvqw
DATBomJGwBq8jmXumsvUIIH5dC+Ku5zpiifKNbUflM0QffeLpLXjBfyGDURlBNHKDxUn4epM6So0
JXwPJ7ZWCrOj7HECwupRS56puAY2g3aV/VsVORd0Wt5Q3ZJMY0qTQdvcP87lprphPTBfQ+EdxpkI
dGAeRn1eexjrs+2R+zCd9P+C+I5/sCUiSQlMOVjd9vOZGJ4JuyV3S41TOfr1pYlvPp1x6wxUopVU
pNyMZ0VG8KxNkr6a6BF+g4QldTL3nQf4UjSpAYgYidq8sMq85rEMEPSjwRCcisna7FEwHG2yL8K8
606uf1MU2vpEnrSfBSuXmhsJ8fGphfDekRL/UceDoAZqbxrcjyhQ/H1XqaapVLtomuAAUIkPe+83
kBQuX/RqzhTzzzGwkM8ZLjcKQZooCbgV54SqJRCJErH/umWA30MIEbc2rZCh3w9+Yql9A2IgX0c8
b+l+cIpny/lbntgNuhCA1u8wlUNNxtlwtJSlIHaiIhvvtlIPOheuzFKWmQSKraQjfNeaJ4DESOuq
B7SWQba/jrF39Dp+E/CpRGdQc7ylFTZdwR2PEEWL5FiD6hQdd5jOKThUIvfLIiLZKXFYHOuMMXa8
uDrkscQZ+MEg+c6nJQpiD2NOYhMJo0WKVkpLSvsGzr1agHYy+I1u9ajm1UMh17JFZ8w4GhFE+hyd
p4O1CPQ1U8wu1aLMWIjcLvBBiBdRdVnRraw5Kxdust42HQqTryrV6swwxCbQs4EUiSxA14hK7W+u
+SVfZCmL8cr0Rbg4qdste+umhRKU35XxrTLKK+tSgFovbuWqfuumS1oMZVG2df7A1Cxg5QgpMKsa
4QYB+2/wCAxOtjvAJCca82WOPMeome6lZaEw0oTqBYvmNiUYXK/rP2wxTPP1IVjN490MnoZaYUY4
pKsGKA8NWqLAacyc+YSfQpG4okT57cwr3iAraa0+bDSzCVxiBpkFuI56cXa9tspGv3gKT5lgpERu
lGOLhv2iKn460Pgwd6gkkLMp0+ZUX7B/fyj7b0RpAsJ0Mf8NRy+sCVDtAB5lPkPAd9k3QYDWrxhi
/AzF6YFn+RzOb0giNZFQJuS6cN+hZmXJXXb2t5r/r/axCLjgRtHLWB0JbL0ysztyE4vXZqFkkyf0
UfhkHgH+ZMOrWpilXj4rpRYBFMuu8k0lnmzOjvnrFhUSllM+cLj6Yu8/0vpiu4zXSz54YRBtJbJA
CPuuWFLsUCjjL7PZuB/9OexMSib0Z9W9qM2JRHzqhFVhEeW8vxwr6Ffn+mpGjViP2z65yLmfa8V8
fVGu0lcz7fC6EBEWhl9geY2axdiuXz6Qzh46Vwa/n9a8MWVJhuo8I081JSwLe7HLILgPW9XE39nG
qXy+6b8vIgf4ahGpXdAMZafSYfsDcZ6PHIkIO8lrA+xL7iEiTWqOwiA/SKWEuTGVf/CKZC/abybc
0mvoWgLGeqsNiXmYuTA1N7cQzQVtHjToVgMeIadRUdykWCY29i2019HXdTfRUAzzY6qjYqmslUpK
z3TzEPsfseVjiI4/b1Db0LutPYok7j0cMerVb+Yf+z9bAnwQwDs2A0mbO3LFDgHB5Z6RnSuzTzXG
JqV+qe4vvq8JpEYG9AnxU7m7lihkFZ7EM/MBnT9fY1F42WhXh4tQ03L4ZdNXer5r3ANClQ6qjZvK
I7/sOEliyFj7LXbg8Mb15v/3Za/Re1+KdRiYeb66myC0Xbicl6MuInfW518w6hwPIBXZ7zrCwRHt
ht5wVTI4WpH9Z9OqItgsPwWP7M/msVfbi15bhGed3kMglpGfNBczGOSKzhOjOH67OKGM0T6/nEZ3
MijDsUqOe5I6PjJ973GXy+0nu0tihadVa8czB1ov1euwpw6+sdBEH87k8Yn8VHjhKi9omYphPGUV
dTgd+J6EYdQMHFl85Tp5h2QJEocoms4VViLHnYIrye3zU3XCTZ/TwBlqp2NeETr/Gq22Bv+hsC8U
XLVuC/cuBEvtiEUTCyLTqgsWw8tFZUAwDqUY4b+46j/05P/6XVD+yUrbbZ+KHycSvfrYdxenepnx
i5492bw3611TZxnnEGKZpWPmVagOT0Slti7GgiijDM60L40LH4LWEQCBOvZ3KwUlQ4dH9LHW0Evv
r7SLplon/ys1VlHkQp44hkA5wBobhdAvVc1uuBk49IGTTz/h9UqKJCi5NH9wIJQKHafnCWhZMhdU
tOZwPBl1UeLLSWoEaOCFY06bGc4gNU6rs78RZ64Op2KSX8Ac6tse+TzTdLrApma9DTbo26KHqmV6
+1pAK+7G9MvCZM+tCwRI+5YupdihBNl34sBac6KYvlO8DCeythsizW0Rv5Ipwx0/zM0EqJelIjby
sd7hzEdZmdEmAeWz7jv3fnPbf7Tt4/Li79poI01y0cIyWnYHgy1L0Em5Qe4V261UIw+8rv5IuNwG
7/viG5tCmzIZCSMkeMEiDPJvwdZ1MBStKhkDlIXL7dqZF5nxpRMGgSvTPk5sGaG/vrxbHkQJFkAl
nuRO+UlD0OurF5eZvXZ6gpKJ9V5rs3zYfpsA6SVGV2KeRn4OiMRRe1QE3n+HaNE/bb7DDVtNfQrA
1GYl1Cda7OelD+o7wSQK3CAwllf1KzW4VMx815dnrWWrFUQEWBbEVHXgi08opFhZjIWHuXSoMfWn
fsXVtFJgE9JeG2jgZWm75Yx6dNCYAp2k17t/q3GFRx3qsyBG3Z1KiorDCjQ7i3Vejb88ud2SRt4l
+Y5dtPHyIGujFHDoqcJK+YJIaHBIf2XbBQPSbzYe1t/kdY/bW7ne2N7YAqKyjjRNVk8KW3yS4OgB
qrnGJszrXBUGdPVFAmZBuIDpxu/Y8sKxSGPlvN9p9faZP2557swQVDsFbwuesdWVr1e6NghpWt+d
oNw8LtN2RC6HQgOg/xZCiOmCCCEJ6sU6riUeuidUVD4pnEAVXkKQhXqrD4WXE25ZKF/tyjE4lYOa
1hZOJQr2904++vDnx0kyeEXu6yRYueD+6LVoR1+2eT0B5OSsJzkMyicM1rs0gplqY/+haTStvlhE
poBhYg8s6GuS1COvgSHDtZ1Iu7+Qsh1ArGisTn5fVtp4nLw6eNCg1xkcdd27kI0B5N6wJ0hp25wq
FdFFaTQ6VyFRRe5/vqs+vyiZThteVmDKI3D5JZwlcaJHQwd/kb4NFdkm6yCZKwKaEn8PyKBR7b7n
Ra864MqpNRBq8p9sZVH6wb6W2IQdm3qmHcqRucxcTAez+RIIFU1uKPBrmxtqhb3eU2rehnaGukKs
vOD4XtPWxCSrXoLUmkKnqdwpL0reox2eXLxMp/RPA4fEwq7EkXGDeSwNZjnQUOp0Rq0qrarDXSwx
g/YThopa7WdSXm4mazQUPdOHLsbR5QozGbWVmjgcZoi8fthbZ/qzz9ycGp3n5ac0PE/4mlA0Cn2d
EKN+Tyrq7ifgfKuCHJkK+dIo5BDmt3z3ViL/Jmcc/iB2MKmypzN+w8vPu7tazrz13ocRJ122LQ8P
u9C/61/61Ccumq3c1ZNtAzNEqk+uVmmnvJ8AVSmhzhJ9vnRGnszIKd0HAvH8BBG4Ma3mJ59XsNlz
XjfwGDgv5JBYaCHCIB4DNDnlIjucIKHoDLKI6MF5V4bj6bpwUXesH9jRMpIJ9sjWqlPJdtwHcXSl
MAkyCgflE6B86+j/gViajsWnYL86GYZgqJJ6anj+0tm62HjuMPTMmQ4UwZyj6BxyGywUE8nH+/Fc
BxXcxkTH/wuoi0wC2I9qDo0UStvPdxi6k2ohTKaU5NNh6v0PoDTAV0di12M3uEAtC+Z5xzRE1YvW
gRFEkWJmdFHQpwOIZ9bFmiKYReFDrHkGm1YgTJtmJ8hAE5ORTiRqMkWgJYygF2WF7EnHl1T6tdtE
d10lAq4Q0qtK99ZD+TglmRCnJsdF10s1KFEdtgh79f5zoyPkabVgnYGQCJh4Ab0rxYIvucwN4CA4
g2Ia9uOek/8Q3e6HerHe9oFc9RuBiMrAENVXjSRozprDtMmDcgJENHAi556eGJwh8wSI1/r2NCox
uaz25OFBJ/90vqfnC7YZv3kN3JLU3rtVAFAIWvi1W99GNYo/kfDCGlbGfirUhsPrvmgk5k5QyhN8
YcW4K3cwIyD+p9bdJh2P3QvDKYGAcHojHr5wMJfM8SxIQgI7WcrIb+vK1BoWBrbFJ82tJRACGkDc
53bKINwlIoJcrZPG07R/oX2egMi2jl1KEoo1SS/HaG/zibAE74YZEh/5mhHPq5Rf9P9jxLAACK1N
skSBFHd17aT8zKfKgIpzuGrI9xiQuJoVuuuGi6JQIhuBsSgilZc5mMeY+z9jfmcI0t7d6GRahx7y
i6nK3dxTkUpfTTrUysi2d3rcUSGZeJNnBU2xSLseK8MmBfdMlu1SyKmqX1JkyZKkdCbN68+xuGbT
17Vn+y9AAShfNgXKRTIUQZsAC/LeVL5MuEHNp0LhR1lM6nlUCu+muPTAGV94F1CGezoKCEOi1exl
dIK8zVlMPcjSCY3hjQvxnLlTujVvDTMA9Z3Kvt+S3aerRaoMpLmMDsSh8xUxT5pT7pKelTTe12U0
qNceD0UL2jQdt/IRbFFwp6DjTJ+czbfQrCWxAifYY5CyqkPsZA2NVc5Ovs1yljNnlC3VmFnsR0EC
iE/wds5iDcFjcW0dJ7X2kKWu/rB1ccvaRS9m6gs5vimI145gmPlM9kW9TQyTTPh+80/Sodqdixj4
Ce7S/XUZTcWzLaJkREmvAveuuxalE7Qoj6iauZwToN7km2GPl0n8jhpilIGdFlOXPVoSnvhQlEET
Vaws1ZcnZoeIlRA3s8ZTQnyP1HGRl31bpnMjZCuFBMeELmpsEc7U8RukK/0YYGcmEWmK+pHym0Jw
LF77HwbMpz+t1zS3RYsKjgFXZ/dogx/44MN27EHmahfTIjt5nVUivOIn7M0prtn+JeJZZp7DX/FA
ru8BflOwbDosyNZqTKXne38WipwpIETPqvzauU9hU+5YgfuEd4VwmkfFEgQFOBTrw0ZD6c8cOt6n
28cVJzHtsTG6wt0sXRv7Bq6zuKJ8CBTZEe94mLIl1nDsTaiGy/SDzrxs9a9TNkbBDT/dLw+z7LF6
FIhHtrokHoDoJbAlwifIF3ys/5S4TDf+oSRI9SGFfjZ26z90CCREUh+6jfCiCdvqj00qYN0oqkZb
gxRjtfm0/Yza537/1nzfbkcqgOvo5r5Zlk6/yeyNiKjTfFvXmcmJExgph8g9qTXBeHWtB6Z1UetV
hUSx07KvxDQ0a6sB0/dLCSStuvmmWZhNEinu2WrTOnVmsR7JZRq6UdAjREQOf9G476sCl0OxZeyv
TMvHGnYsMJt/Q4cvlw1zUc8YMCKKc6AXy1hGKf+PjYJYGvQNgNuUHTI7zSpb4QokXODQXYAkEKsW
pGWNxQPr6aBeU16bdWH6bxgwQkCntVHZZZ4SWxtgxFKnXD9lzj6o0mOeydTMziSTDSjiM+8d0nR0
g0RPFIuD+jXJYDTaaB4NSBZzyVJMDs7JPhAwX9eim0IIAdpAoMFEjUG6+GKaitbsjkfzfNKMNwno
iR0Mt24u7PP+lkk3AG0LbrNaRT855V4TOz04JgdHciDO2iWo7i1qxkhH3kiQ4Ls3cnd6NQRj1VVD
iWkcvtJ6tEt0zU7pT9qiRhed5UFKcFHb739GjHOKtd02dBkjkvuuAMFxv1JUWEmNq2meva9znRly
UcZO1pKUXSjmxuxbukvwnOz4nW1ZM1ZYBcfI5jJwfVD/7E/xfC22UnRzAZADImiNQh7Kx8cIi0LY
5KRmLLpxuMWD2tO9v4nz8xyddtE9DTlEOim7JNZE2bZFARPT3e2heptlCLiy+BcgYDdO3tbtEtgg
3TSys4cl4bdV60eaL0SR0ajQ98X1lcCrFSAA9/keaP9GNeFGOO8QDYT+iB/8gvqg74zLx/KcayaS
LlKmfk3YNKdsGodm73977kib3OINhznQz6gBZhn2Edy/7KrjUYibnYp93a/bKhtnttbuPPhGllM7
NRgJT/Bg2nqy0WvYJezujm0TQZ6fDDHYAraL7VmpsYWVyz9s3RgrmX0A8INWzmYUPTefbjX6mJ+R
IjUh2Oe9CO1Ngj3jjSCS3mlAhfYa7rhcLmhZVssUY6bfzcQ84e1zZ6ajGT8GHENtNJEsNnQOIyIB
LVLWR+evdjC7VteBypZi4lkTN0pDYIukJ6yy4aQe5OXHzIo8jcPWjh3ziGDFuFl04RCtfbNzgvZA
vR+GmLTZU1QhQc/d8qBPW+kY72TenujxXJnLoaE/dfF2UFq9wd0tozynyjcoyJpnO0qxdzpHbRpA
LPGTdSh8YezAztpq/fNf3LX1D61vLYLgXSaWWor8SYmJ+37Pm+pHIt5T5/PbzdSbytlziaufx9HG
Dm6KbfNFNJU9M2FsIXxU4ZZ67OjWZLopzux/AMO0zkNofO3Aa3TPnWmS4XWqneuXw8n6H9wNOPR2
h1Q9rqrEOQVvqY63m3rqm9+iwrP3Xq5bN+I8kTgq82G/lgLKubU2TWuNHZDvjf4+ouzbp/VUEeBw
RaJMWgQf+mXAF4/3lpnEdlT/D9ouAmM1+szgHEr+OiL9rnOLKZOb8YtJzaxECRI+/d5b3QVMqe0h
pzKMquC04PMGzWOsRu+xNqbw2skbe+LFAWiKpcqmn5N3PSJKdyksntnB4ubmLpL1Ku7kPrIAwXtd
ZoccSJuSb/WCItIDUwnSSOjwCphw+eWg2ki6oa4/fJ7PVPxY0hacr5Vj+3S2cC3U1UBqgxqvIr42
masMwrknFB/PSUUTz8128zn59DGDwLjwgsdRvduK+hjkcG2q9loO/8stSfx5NBGJre+8CrY9NcbT
roaflfqo/VROzzNSnzwgyAgI+6gN3pUyuOuIb0HyTOefCNc6Bc36dxivVQz1iM+kTRqq8iEDcS8e
t8nHbSlfzp69bwU3G+q2LCLS9wbCRF2MH//d2Eswyi6nfC7W+FcUWvy25C4q7T/ql936YVlkQVNA
S3wsfT0U0gCEoXYUA1mOjC/FrVyXN1GxfvFBLf1nipeT1MTsUYFUO6XpWh6tXefYIJsIOPKX1ypb
5QkEgdYLcVzKz2k5WNpDY8pvacSCdTUVR9YVHiFMdJDMFQZcWVm0EOKYYwH+ebSvUkjjHLS4sG0y
GKM0mZvgjQWRYA/V/hXVIKxumI8XOAitZRslk+DJpJPwwG6qQlmvMm2LoE2a+TICM0/BMbtiU18d
B1mpWzTP31Lcj/r0iNYbtQ/LaCKQkZFOS0ryMqJNuKi/DzCMXm/EGEG2xpEoh3sSE1SJNF7vcXDQ
XR6/0aIzJs/rdVc5Gth0mfOfmdm35z07y2+KLToSKy6uhNgzDLJcL9FMDRYZFJWubqCTG5RmcpU1
mDyl+enslhmbEfRODvNnusWrE1UOcnGXQuAb/YHAlWGxWAbTUxNUCJbnXZXfJD/n7ZREMPZHeP7P
OVWMF9WsSuM+JFfmL85zUn75XBPmbvjEeVKPcbRqITqzpsptyxzbCd9McPYTjD9g4VzoX9dtyXuL
fHCTTZfOWT3Fbud4buZ//yeuu+67+pSLP03hPKmjODKPOJSxoYyQHSG3X/LmHMhfSz6S8KXmFlRP
xH0jiCwOQCyrS3EZbPlzxhOh7yYAGa8/D7JYfdKvfB8f/UQqTuoFKNqFxMZbXuOqoWFF6S1U8Ab3
BMznlFwdS7xEdWZ5hOFULEwtzwuoJ+uV1n0xfRb62DQlOXVne6h/5w+zlmava2Yl7+7hS3Jkf7Op
PzoFdXA2Ngryqi+YljDGHcgfck3r61EsgIXh1gbfP7ODy/KVpTu7aM0R3kDAaXSJMn0Kv92P5AvJ
Y/kXyh41s/UqzNpvzCA6YqoL7ukzuaAdwgELrFMTtoOSRZLUvMpshypkHLEqn9OphC0qD3rbtfMC
m1RnrKg2OrzNzVqsxa2Ndx+Uc2E5JnsKr1oPIFmW6v7lhKggRryuloEqJoMHTSNnkc8Kap7dAtFp
KEMmtseF2fw5x945AIl1s17CuCVJ9oB2z1NRmyihbM+NP0JjO9CzXiUiR1zl8/HTN0gMMeSFa3wY
wYfwlIWylySAj2gtBoIK+vJXmIVRunFLfecKdHHb/CohL1ZxcSwwt/1S/QSz5FhUzxm+M/BOQgCc
/Dn6foccgU/ZApZP4mVejaLVbWkJATpRKtLfmmf+jnUmvso5IM2FR58t/206HbqCKdlP8zefiYiE
BJ9VBCPQXc2K+VM1LrtebZ6BWb40D4qJARkMz0VmdUjcK0ZLCE3A+HcaAOi+O12U2azDTQ1wazzP
gkLrfT+n/z2mC5hVGPVhp0obxCylY7d8VCbKozB+eVBJWGIalNPkWAuOTZ69yJsE3qe7NsLecL98
xmIgLm6wzTK6S0KLK/GD4hIQQ2HjxwKzMaFUl1g0dgRmrKmgkGPBd2sg+CRFFqeJT8EHieLtJg14
UXP7y3xwr7WuOWJ5123pnQetRNRbUr+wyIlnNDtigCr9Z1gzSSoE7F/5Em16eenlJUwc6QdEPrNb
oh9pRRdJ3j8B4xtTiOBHbk75AAOs4/Rtii8LfhhJjBkaWXn6zDXDHGu0Jnzb8NHKHmj2p4ZQzBYt
8qUHfgrH6a13fLNuFujNGf6pcHmINe9Ogww7kDZ5GeJfYE9QIeraBBhXCsDAY0kJabN2BByuUYSl
Kq4ttogmibYUkgXxar5xgNE2ZLIgbUUMPmSz7Zi88sgD6Yl+cx8H3oXz5ka2PFPFazzBphS644ph
FYpkM2lNOtkIRpjOVytNHTQfeCLU+v7Blm1PJrxiRzM5QG+2kXKaKYLlNyxfwVDY/h/DLVP4wswO
OQN6MsiJcBgxDST8KvHuI3u/W1zP70ST6CBCVUDh7yESplENYVgEM6wgZxeAyqC4kxo6krKjJhBi
77CC+3jLgIlN0mFZm/7A4vRQ8DLIQFhsQw7A4Ug1g+WKaKkvTk2jgNvKncvLgjbT2yuv7sZqSrrL
izRapjCD9VHYo5Wk4VaVI2BhXlSYpAUZrzW5khvYAxSd+gvW7SFF2A9Fli5DNn1QL2YEm/2NOQ1a
5I6+gYKupDn8+fDiMO5ooT+WAt3rAU4PhzPP9Oqn4+OIba9/ES4KVeD67KETbD3NzQnsBanlXPQF
J6DS2oJtAz+vJgsVzrj5USyVis4aBeNUKwOm7jG1HBDmTpacccp06CoMbKiF5DB7byL4XtldDfnl
M66DwbAJP76eqghsIYvPn/ryTX25j+kAg+RDno2aRpV45DRNw2TL4hRF9rrWtEktLGTlY6LaGRoT
m37JiepowHB0NmzMJiLnlpVYyGihMSESrOVvnPGQG0mNS2gQQhhKh0ZSayY67TvLwr0ZZUUWRdAT
13blkEvV+HxzvsFHJBMmxmBSFnDZCQwqQPUswL91VWr/a0n5kbP3qQNwGptovvlOCMOYQTWOc7KD
twd+H1ApkSeaN/xXzhp9+hChyfouX/L3NaoECSHP6bMSQ+pz9qSEClm8qOQ9k1TMaBTAf0nFbrqg
BfdMM9YEY0hC2GLbWwk9/TpAxwbe2d022gXpCuoSnyH+9NS3KQwK19rG9z1qy31bwIPIP0bPA6m6
P4kFfXIXR+PoFNwXbTC+zvmZnZ4y3jn98IbLWReJUUHVgBTc/ysX2R8209KQB3neuoJbGF9S/iuX
ai/20pNnt8+QUFL8+kwOhHgR36yBTHLthqZgmEvIZeMGpQIWW2qh8IAjfeGKwgIQ2mnAU7xtjjnB
8hZfnJ1AR8SlDpne582rLqjJGp3MUtlyTJsvBCmX3DBtPqF8+Pmw8im+09HZydvwbZ9pXHCXhnCd
VMSKCZ/XL50cfYa4rZ7x5azgEeN1uqcxfE65pbh0MRx2wRHNVEuzpmkaQjUTXyNMP65ATzS4IIxU
UKS0jv+ujbCcJEf1VQ1CDRkkghDfg0HB42M69fxi3/Qtu5N6gFNNlXWKWO36ZVWeiv9/W3ZX+Q84
3s96o8l+KJu8vWh8qdhMHadurE+3zmocXVJYkLDtLOvXtBjCAgSPti7u/DA9ezgZD8cLFiCM/6t8
tTHwkYqoKf0O2wnWA5Bh4odOFRoNdaLtIdTK/MaMvKHBbDRtnahWOwwOVa+lWwDmJt+QcD5n68UP
Yep+BgWqpErSxilbviqhvqG+kHhVc8ihoO7kxa9hDjKI7UN5M/MZuYL8YHuuAUfA8fZF1YndUV2E
/iU1YOmB4Hvv25dq9BDe9JB54IATPWKBVDMZXRJ7FQgVS4sAxw99fX0R2MZQbPzjya+oyMc2OGsc
blq4JrWEOdQEjajkheDE2Nvxphvh99cjDdc1rAIIzj0s9jLKXKwUJtjpTq+qr3RdazxnsuFJ80+8
OyIlfC/dq6EOvwiBPerXDHqEphjkfGNjxgJo/EHscAUULQi1luZlYrftzsUfTSDevObYoOnC33WN
Hz1u7I4qWAvoioP+ibC/1YannyHWCW9/1kwTXW3XSWuTYkQqi/yWQgxTzL01szR57R384QDZ2io3
IAAdNTZAtzKBu9HORGQSvuxJvSfqRdyRzRX7oODOyhnCufN4q+f+cCZ/Du+egZbW/nh+fjU/w/H4
SL90oZtdO/queJpkq4SG+VJbny5UuyNj5FiCMCIJWyTK4BxUF7RGUfV/ftaxwe3x9UDBK9zXmbYx
+kbUS02KUosSy7yfdF+NfAg5oV1EYmSH2o0Y/C2tR+35206FAYwFAwKpgyZz3kDfTGpUELFaI9rZ
EcQriKW+focPegBasKbSPlbqAPqLyZbwgYz+v5yDdGdpNIWH1gr5ps+i8cfVsFHw9J7R/UNe78o4
O+yzRcKSbSL0yzY2kaIHhBBtZTo5sEIg+bkFxArNg9bRfhPOaBFL2IM5AiT6bX3sq78Ioin/dPFG
CAhdvNrqRqlzQEbmk4pFGT2neeYcUrCZhCdyq6BFW7GBXIBvBnMvQGCM7bEBv07/OODIdRO2yKMO
98Z0DG18G1Vn0CkWnLnNMTbYyerS1yn+xhLQ6yN+kcCw/s2DJINww87LxAF4LPWRNfGyZBrD+6rq
/6JCHugDN18VezkdtgvP+MwAaQAmq5B36j4R7EulWf9CZf8oWfYsw24MtzuCe1yywVJEE6zKKFeI
0sipQ0nlqB/k4iIKuebOVzVUL3s50FCINxTo1jef+gWZHq05ftt4g1H8fltkJgTYTn9itF5CQeZq
Mvr+WhqrqM7NVo9rgR2bJmQm3mC+YlSeyNKzlkKGXQOf3yY1tJ0hNwQ58T2REtnK8Fb33Df1Sm/p
WfRicXsIMD1rkoCUqLFNu2b60d1WAp4O2RGTg42v4fG4jEpLouxGlWcKh4527QYmOB3AzBN2DN4s
QvzF19u6gbFWSB2uC64b2C0lXFjaja01FBSEL14m3u65/1c+oX+ELQ2TDTy7wvhjt6/G31ebDodd
KSV6w+tTop4QGmDt+PbJCdMFGHUrLyGHHCVkqM+vuEIMYqMPR4wbaVhFvzskRkaGc3ypE/lJitdn
muqdHCXzA9zkMS1i3Pr/6r3L7kPYmBvXSlYyn6LRB3WL9ZDfHozK87V/RrTA5AZHMgZ/E00e34mp
njiDjNFn963ZJvM3Rf/VqjunQ2sx1UFCFA5/5m6N2mYYfTe3sDep1IfZ+Vu3zkm5iwGwCZgcwGxt
rI8VHbRCAZymaI1oUp4W7yFFvcsTiDd5Q7iDHY2j8Z4Y60g6eOePBq0B2nlyQiQdzORSWwTOm+jP
DqXOpMqTG+UZOt2wytLqTvGCKrFZ4lGjpiYGmH4NuJ9fczu8wYiJqhDgfIjQUeCUF0wYetT2oRtX
YaIUpnt0O5MBBXDoK6eSAxhYboUe1OanAD+br/WY4OZm1Wh/E1Hqw4FfW9G4WrTnN1JPKrzPIDF/
a7weAicYg50KlL9fLIqSnbnJ+AcUfdQvO5fBXMsHk86gh+RijcQLgkCdxhmuerbZuxaN27bnxryU
uzoqJvjOokvnu4EwusOHVw4aEpCJ9jgeLj/Ttjh4kyJz1dWYXp/lM/+DLwVl5tLJ1dFN3drqQTIb
IpzLq7N/KTWLO5QUWZTnI8U43+/PpBoYGbSgTXHaaLmzyla61oSw9QVfBI7B6negxtDFHQ7caj68
QFoI5LlBsvXalrWwZ7InQmJ9x1NIdYI9PZJffhx54X4b9TXr51zIu/eWw7RAw6gb6tSa36Zv3ofs
4UX9jb5KSHmiqN5pfgnaCJVoZFCVObs+pitPZl1+q5G1VoiBDb7Po5c7zzTIvvx8S9CVRgO/Flya
oNklR15qboSVa8k3R4zhiKZ9mg9GBy5nFd2vV5aVGQnXLswQM8kbaYiMLSzwva8slcpJJ04iLn9x
Cp94Ee5UIrY41hkV0f4jyoB+hdy4E9SL22zmzM7E3sQoWhIFUZahaLnoioriLygHEUAJyTAPAHFe
6fvTt/etOcAfpLw2+b/XwFdobiyEs7WLcUQV98KAX0P24jNWwzNyMjpgBNcMiFH8STBi05FdghXZ
EOmbxXO+cQQC8+Wtfy8o0J3ElNp8O5inbeLxlnylcckRuMRHihsmpLqg2jY80Z/S2eGi/HPN/OSY
FAw8rpY22OKMo7RWw1p6KVQTSdEgo3ueMFL/12KgWSSP6xn69QDupg1oHzpAKl2Zc6MpbEhHRoYn
9U1goenmM9X4fhVF5a2oTepT3LrkU9/jsHJunnpAKDJOL4rQOT18+cGayvDIMi3n8iksKndKOGtO
9ecAJ4h3kykX7P7e7vk+kXv2a4bJNK7rtBmaB+vZQI4o1wl7k2I0o+ythiwJ1BBdCCtFZsWuq8xP
ZQAgGQ4fFiVa/m7kaWm9tFdV7muScOugFKJ8uMxDwPOWEY/OydAspdwZnIvXp9cICHRmKMJi2H12
4iI4VyyqVoTn+fiqF8LRvhb9E+gkvnHUJjPt0hqPQGlyH3TbiCC8frFuKcKU7EGtgJ2qhntB3jyC
nWn3KUZaaKehFG5LKm6eEfkdPxm3yXDuyOv+gGSCIIghTNV8QTZNW1v0JKNWNQGPJjyLV9gfk12c
es2ojgG6mrMJxkKhY/vHhArzb5A1GOGwjLFsCBOh/t4uXhoG9/RJBpupgbqEHJy4gUhP/7Om9aPD
iTLz1z236mLae9dYNn+ivOYLAoL2rrtwjNOpc/ypjdF+6We4VM+13E2qAYvl+Lqt1io2/fBKXcEM
5HiIHZZweG0JFCG0XrpwgaC22ryAap/r0NJyT89G2bcVrfjUCOcvYsShYtk1lrXlt9xorzKEF99Y
ohMXLA9Rtt45QCGvuSfhfPTf2duOHKooFPBcyp50WN4OAmQu8od5QnNXiTKojqRF57RjSB/2s+DY
j0v/v61XNLhOesDklOAsdaX3jzUyvjEP4fZYe9gGKMHR+aCcI71Z3+5R/8j70GXlskYMsZWIXKvs
6eHk5zr2XGg2QTGbPFimthwsQ54UNI/VAXa2iiu2dVdvD1EbJlA85hXUvWWQeQdXRYwYGLzq7Puz
Fwy3tHQ7UfwcGkDtGHsTwmzq5wD0Au+GZKv7BlcbvhAGvj36o3MgERJ9iJSiPAiiePzMqIpL4SgE
4JxZ8TWvjpFkcEkslyxNeDel9t18bBxFLTN9JaYSwBQCjKcXuc90dHxxFF6wnFEtItqOZZVrUGww
JtQ9ixLQmVMIh8lCpMBzkQRO/AaVFmK2QgtEA0zxNabN9EJUnttS28N+t60CBT/nQHYE0B6FduqX
IcE5fLPcqmxXEJsJjFK2p5zuQ16Gl/FZJQeORqNq1jUWM5obCKAK4o+5hb2epgqx/pSfARPc4Zn/
cyWrgvK2UqFhG6aSTQqyoGEQxCydiDFBCm01dQJ0PJj1DDe1lgVU2y5a5g/J/SA1B+DVstxZzQ8n
4VsfAr2YqXpsZCewVGbGHgzzHf+Nfs+ODpKeR2sdCEvMTfxjVqjuFehLKa0R0Kz24qPW+P5Mg9ND
X4T0eMeFQN1cZzCU3mUHJvKswg+qiFEleK14aVaaLAZRFdNpeWeCBGLgq7jYLx/FyupmaHzNkiT4
rnz6V4qkVeOb3g0KeuhMmsLx+CSPBIOCAWphgV4Roy3EULhQzFU6FBhh9TYyQj8LO6JIwYkKPvQk
7Od/eZmELBVeBzOS4DEF/Y5ztwKIQxCKrjEylG96HiZeGspNTpuLZ5w9+3IJK2tJE+kg38Robes7
wU+h2nzHXJkCSWo7IMDWtDnhRfdnds1R6G/ASeO6rxi/qCkRcFtu4eGTKMlHy1VCyU+aaHLOHNdF
5uACa/yMXSB2ME+sNtSyblY7TUaR78tIXGBbjZY7FtX0x2abzDK2Cbg855sAJ24cSzICLUd7q5VO
1mmuh5KcBkdxuHf1iP2DNIM2FWIVEBb35jnbCr202Nw7JHcgwbgutNXP6g8QgM63i4cBKDDPgZCw
7INEjVPAdbVa5vk+1GeP795N7N6HYlYDvkctSiEyvOOFBnZLkuoqZIQpb5Z1/i5o5koiWm2UoIc7
Cq108sf9Nv2dO8Y9kVgw8QRDNMD+0MiHzxDD0djfzWDNQrQTeq6IiyNooN+GfnDfSXBE0VxfCHWZ
KDFDdJHk4L7LYsX/2NAN6Fim0gtBbtBttQyCZ2S0MYh+idhmai0azITZFAbWgt12AjQAfsZkBfOT
jZUKANMF6hJhB/ongd/yFWRaGbbBmTLrhE4p3h5Cdef6EqtQx4vaDJnf6GZUyzp8Q80a6eOrd6a5
lMcR6eKCoXF6SHquJy8ULBaJfCX5ZNFQmOpPHrA7tmIw5EnGIORGdO2j6xbcZlHVvSry3bbg8ffH
bmOqvx/dM8zYfegnt/6ffZ0VgWtsQsUMYoCZfCTavednBuop8SmGV6X+WU275O63ZWLqPfi4C3nP
rUmX7OabTHfGKOQ5PcjEORKvZsq3eGAt/3COy82AfUI9p3lJXoJOJWk32FJQnPucmGNIv9XFmgn/
D0KL2E9K7Xr5LCbAFs6sCntE/h/5eCD9HrfVrsAkHr6hzahP5EWUnEQ5cF4QnAkNkl4XmVieKrrM
0MXfScNDWRaTF/XebwhFVSOUODz/jiIK+hV5ChR0BZiWekP1bSqDTqqfZPI8WOGfdKiSi5wM7FBN
0B8wq6arGYYWC01+qWR8xJSChVZrqO0JHnTTXXt7jCQguHnZKCzRVnBavpg4UhCk3PMa8kWutpJz
Ya56uEN3OUcdfL3ZUe6sj7V7GwWPU4YWCyV//SUujf41GrNkztqCsQb4FsPT10/5AgRKhXb6pk0r
D+Btu5lxjBjLsmfO/vUKrG/A9IQ4dYBqMgYKakbwMV0Q5t6CVL/g3fTQTVKyol834z9SNWgDvHaf
GbVVNsi9M8HIySz6cYk4JKNSmDI6oid2moLx7jclvC8w1hN8Ssjb3prcgymjE1wKzmPHuO2FiqnY
qaOVHHHV6+phEpUYkwMGJplux6+BviYxRsBjycQ59eetAw4R5rpVbd2EaTy56uYswHnw+6KeDP8+
mdVeMth0WlQ+aEI9zIn8k5G4sX3X/wWYN+K8muUhYNioMia/k8bWv/AjYR1qQ+Wxx5ee41ZWbi3V
8dNzxxpjMn9gXXf6cwkGC8ynlTrHacxLNf0SWzwWUokCZikJv6/J/GVHJmOJHbAUo5Pex2TQ/edd
gLtfXY8iWj9usXFn/tq52NXjF7PvuBDpQ9zmWITSKdSZLAjiiZVhK/lMSWErCnb3j2Jkf7GlrRns
umqRcCU2JsxIJUd/iMABNC7wtcyPMI/VOLpL5dqhYBzlavbnpDWflOD16aQvQq9W5NGSAJWb4ypJ
9YVi9MLPO72GdE+iVd6ftAtwaadMfooY21xiSeWN5IN6U+uBMLAfdDxIkb4klSymlf/EjDglmzCf
dTpJy3tRURvCIPpPY35LWmvc//dryGoyei0NPGCTRgjsV+FlzScDY64ePnFI3N8wohYH3EIwTs/n
7oM1ksN79XY4Uav0i7cv9HwKIXu44ywM3mmvavO3yQ3+mi5e28YjF0BYBGl6DymrdBBUbvAadq2x
JFRPEFjCXmuafRjhcHE8IGxfJSB8HecDWbwwdcjs/2Rvlj6tiYx/s/Z2BYqHlw2WEk5B66NeU5Ue
2vEmDqOUdfxkqSarS7XXIiyzrs52+wcK2RDmmYsfc1SOJUsw9QqwwKzhC8y3aJs4vJn3nvWpzSMN
tZfXTzgjZAM5XgxRia55MzmkZ1co34TUBMhTT36DcXvanYXcu4ZkBguFJ9gXnvlDs93sCQ0QVBp9
FfmhyjkAV+gmfrdGstRJ+hJ9IyE3jZAltn9Kfr/kEX21wkQZArmk8wUfcua/NUlbNys9BZ+oMig+
F0B1nKRtbnYEOON6LHvACPqKdnfwTNN0qh/iFJQuf29OQKCsC0fVNC0Jzb6EyIgMSCAsUBH+ulo4
AxtPA6yOiqG/XeA2WBH+wedHT37bQ4e0Y84s1QQRSo5cIdPd5Pdo1oKkkn1e160TNvze6AGjGeDq
v4HLvFROR0Hf3BhmT4Qvwa+WJ0AtP8cIDEmQvaPtWzVUng1caoYEiOH2IcJsA7uS473JlSibWlVX
M8Hvh6mV1nFnGdrCY3SuswOR91jtmEDLgmydQir7KRA3uDiHps6gH1yOXeHok4dlMROaBfU3ZflY
xvndA/UU8c2A5hdCEYtZnTZBOQ2qqhNuVh3bfCNNvk7mTWJXnSfauNjQ/UwYyx4HiT6lFQjXwd3y
KL6Y7nqCDjYeehTnk9sPMRHFJfTR0TFqh7dkHB12PuXHwvntSa9kpMpCHvLSgAlF+XOXzzg16Uaf
2WzqO1REj7MoFmKevkR3hd9Z+YzJMah3Z+6LNTYiSAAzYopGTEytpdQkiyTKATdyb8OU/XqGZXXV
9LxQX4OhUuQ0ArJ5fSiGgeYTgF0JAdzuSGD8qyu8b6Dla6X6FIiN2ciDE7+oeEQXU8Son0HrEgvx
oceRUoAMcP69+BqBo0LADr3CJd1AqQLAug+fCTkuNu0B9iAaMhWVTGUQGddMQM7Sv6WaXNcnWekx
ySco1t85dBX/2CwaNNosGdV9EX7FL1aAyAHBQDiGuE691Jj3QE6bbcmT1PffGMduKnrsiK+wdST1
sZ+j8vHa5sTpS6B59JyR3kZfLi+sWOzSruPwIjQNWjF44WMWD+Tx2PTXCGqg9gS/3G46sS0sfaRe
wC4CH1E/tMG33EVnKEOM5DMpiK+KVSP9bMem0lLC5AzhGOjuHVwijCNIYHR2T2us16R+0tTOQvTo
yu3BANTBqr2QdW/c9kb7pXexHzBZeVz6pYMp6n6RYsA098tqf37V/DdZgapO5kBAOs4RLkV5h2Yk
q7HPqPVvNwY8oHVnPY8ALnEAi1+kt7q/DhRcNArr0f6C7CR+isOVAiGiIY1sQVxovElVJviYrvSG
SJB6kkMjwq2sPgslYlM/r8BkHbh1x6uzGbi5jd1RPdMIdTT21kJN8ANZiRhGYpyiUc/nY3UsAcat
4OUghA6zCkzAqynxzdXSDY3UB6avW7lhZsTtw3Yd+oupQbQ8jbLykDB+Op1Hg5deKuFu03qADvKt
n5RhKqPI3HSBqyzQsLbFmg/Bicj8mdn9QD7NcLAk2vFFKScArbQVvRU4Z0tJlig6LsBSoUKQ0g9v
UvDg3CC2bJhwVZ8cxND0q7JBsGbGvXiFpxUtMZaCzE1PNAFotX67uSLXdAp0UKOGS6upL+tLHhEE
9XtNo3/XvRTsEnits37laszdyNlWTRKzEOjMSF3Qu3inQnhODDyIq2Of2RI0899MRjvuW+FB25lY
sofzTj4CEmeHhF/j4AA9jD8aDxxE5Jc3pI5ClPVgQdmTT8ysB3ToxCIzUL+xjdzqCvJjNMBdRlLk
c7vkfdiDxdcMeSal8Wq+PGlVr4lLGkKqVueUt43MSzi8VciIUXBZIPwHpzy4ct4V8LgQPEh/XsR7
OMk3HSpw+OmY4udglx5byd1QpLqhc2NBvsdHpdbn4ZjXU553aW2kZz+qISq+JxJECuGMf0ahkOLM
xxdpJGBuF8KzU0ce9oompNubcMXRTqZ6faKcSEOz6cFCkxiCfTVFFj1kalVKbozrXGgT5Ttp9Enc
lwL4PscJG5WbwoOEROr+404trSivTocLkw/jDFfhEmTiyc+l467s9GuLpZiOAFJyvtmcli1p1TS7
T3yFOAblL5fUP39T5rjgDiM6bB90lIVXpmgTXyBqfKE+VerLk+RtxarWIZx4YZXT5HeNwEx3KgeG
hojZIRB3jnTXNiyC7BHofJ1B134dPh10rdUlAQrmVHrzdlteqk4TWcIxNxyOYwdfEirx9qVYpyGW
ByW2mSYlug+Ae9A9eFetiqy0SqhrjCr0LIqQv3gG/fuUDLQK0gPcyF/t8TIFtGyVOirdZp1cZa8J
+KkLDBDQEp03JCHRBoW/LSULHybczLbQrzgFNbv8nA0RIX7cSr1041jcv4XPrR29Nykj2a/QuERH
sVid4iSoh7GkvujM5B6hogTfkaaE1EPPTgzIyvHvNznZuF66nQXdjRQsDt22rpIhA/SZt+nZvY6f
hIqlKvDi4mpfC1ONnxdyqIOhV+P/qlClyfc+i+JuWTNX0H6aUmXJS4bISBHyV/IBVudst8xeTSOR
XDDKu0L7p/VBeYHVtNR3FetTw9csd8v2sUyf+b59Qs7ykLt6oH1VVbD5PvN4N7zyDzR3ZFsYe3j8
7xaXIK+agsi79/Gg4UP3/OYcJ8qboNlY7UJWGaTWo2Od6NEH/Nlk6dB7+qbC2IRo7bn/XviL5KBs
kPukZcQcF6SWW7uaA/JzP/pI2pKENWerU1JwiDS4hmf7SqfBZL+4lVOqmHcrwMTGbPEL4yQ/t+q9
d5xLASjH3q/VTYpaI4BUHELiLoWoYgfBBkxx9DNQJiLp5ETPraxEqtgdLTfbVh5WFDVEVe93LXZI
3ztVfSn4jvkcKIPxrdfkX+oDhUWAhbsLgbNkAONUypafhsa8K9JibqlkFo0+7QtYeSBmeHm9Q5UU
swu5KBApRVY5lo1BXiYcbj3GZJnAQkZ84ZbMV5g2QLIcQTI9eUoSH7vrcGYTD+grvgsJ1QVGLYkq
GkqXvfYCusmeSbLb3SPjYMJ6f9VRmO8i5a0sP/MC1MeVG02CV6GdwZ2zqflXOrYNFTE/Gbn76NDh
30QimHw7cu4U36kDZUHjlANN9ynU1UmxywNwhf/ecAD4C0BKWP5ibFnRMkW20ruHpjzE6puhQyj9
kCjT4rcETuLZO1nCsqLBYeYn0ZkTXxKYHJixfSeFDPYCCtth4SUFR38VOjYw63gm2QUItczQValM
aXQr9Ah7JpbrlT5pnosM5epiVqrQbrBcnKAZBwiYp5BQ0jjVzQagjgQ8c09o33S1MJ2QvjtOtBol
hFCE7Dw7Qly5sbTEh1gCwxcE2OgUsdh8RXm2OnW0DtMG6KNQs5w6bRbWUo9goZz+Xv+gWugNsIRQ
6dq1IISGCz9sHJnvHpZmneqgUS2sNJqTTOBr7H0Y4cJDrZEqYgAftn2XDpqXuj1Jy0PJquTmZva5
QxQ33dRObAEFrfiwIiVDfiRFKBUC29lxAweoYzJHKba0vimKVhIqqRRvoiVjoKy+1zESwccbB8Nf
IYJMhoO2qNmjuhkCgdqhZEEAHJxytUbzSJyBjn6H0PCSodid+zSeMec0SE9tN6WFdGUjbKGXAsBa
ZMMJ1jbrPQcI4DO9NBchxQBqKVCv2Dt7tAmkXqmMVafpTbYDemGelQM4xs7xO8Cn1bSbqw7/fNq7
EnMM92NiBDupPhzBnxwLd/Ml6u7Tn3n+KcQ+0G9Q7tmeznUvgmN1ULos21FJkTaqh0ZmJsgorSZk
elRL1UNG8hh6o7UNEAMtfaTDhyLdtoPXQ2LIcediDiNmjPRxYO7Ms1NutQzdRIt72P4oRowdOV1N
G+C3brdKAT4Ff9EIfXjyOko5xweoEZUCP37yCW0itk31fmTSHnSF9PAZ3nzEFjJgdus0y4Ec3+Wc
pj6xhT7FTL8Bre8suT+9THWO2KaoBRBAshunKzSYgowAc42kh4/C4/mMq0zoYj9R92EZszWJEaU+
McdKYh+9AnyjDm8rDPSMseed6PXTp+fdNTpFzYpySqMvPyomKOVLYyd1OcPNljeV83LyBnwp1oTI
1x06S43SzwSr2R9PbYMgTcrhUdmhGifhOrxt+CerTg0VoGyoSliMnqjhxhKcGtt4JF7QcLGp1oaE
yYl75Aeejford+kCaY4f08yFDeiKZJofemOFuhRJXtMNVKuJZGqTkM88JdCO6aQ9q2fYTcviIl0X
SKK8Od6icCV0KsM9pitYgYaRyj0Z3xKZ57fl3XbSr0hc7JOOj0Kt/8gOwgGIbgAQGTDN8uMwqzoC
VV0nCC9R6GeQ7MJPRnJWEOBHDruyITrwYOVLLzn8Cpz141r//YuH2VWL0WTEwPzyXT0AKb7mtjtN
YdkGxyGqZqxWK5dnROMLGwI0noH/00x9oXqNcLbmlRmEyLVAFTgbKuNeohtM+hr5EwEgbK1ntsM2
pu3mrei1yX56waDCZg+xds5Z48yPnNByzS9CHy9bcSd2fYotmjuUkIwzmJXCfY3w2enfr0IpWta7
fj+Nees5/H5v6RqtPmL/cNsOjN4xTgFvQ9wxBfIRNALqgHw/oKrOn04qimYNxlx9sZZhOulrYqlK
PgBh2UGW6QQhUd5D3+ARopA2/qY5JZm7tXosv+rnGaY2S5NnILfCwo8Xnrd475Xr+vu/ohXvYqRP
q5uNczj9ao/Rk54Mq15XRhXch2BK+zWD90eeggPrZBn4NKX73uo/hc5nZafiCuzd861/FKnROQEc
wzB+elOhy45KIRGobSb5I4c2j7IkP7+MqdVetsLHQIKHfkV/eFU3WLuYnQEMKQrVY4ZCflgQmPLV
su+4/ztmQCGFLojWzLDXq2H/QG8saBYIxykigztnn7gM/1QpTCNr4F9Aa4GCKNVkXVhWRP0JHdRg
d2wVN2yC7I4xjNUqgRskuoNvFumjeXMCKWOsvPae+obrJYKhkRuWnWw+FToU0DNosJuYfKpthzvB
U4+o2VbQgyWFE9D9rxDEODpbd0vqTVgyEgNjG/mAr3h83oA8NB3oedu5niy8WpNTIgQE3YRhwoA+
h40e7q8qCKdQqhZr/BCvJ70aFZv1VLAvnxaxj0a1pNhL9qT90SCAVcZ9yLC804jSvfve9PXah2Ms
5dhMpGIK54/mdmfgPOKH/XtcNO258rM1RwjK7+WTLSx3eA34UU71ltSSN40a5/9h4T2fEG/dPEQB
eFqfe6AXNhb1lI25wgy6iv1Sv6I83K2VXh191RmLlbX9Z/ScOFHNhwfxvhQr1T7aOOVkspqwp96i
+3p+sKoSDYJ1XL448fnlJkSOjUz28UsR6hRLg2ObluBUIdpGwz1iIcxrbrHu4lH4LvZjeOKaNOQy
BYE2roc8El8xMK+XO4YP8qCOiy+yeCOnGje8Wt70Xoi8KJJhvrgwtfgGRxxmxwXRU0lDAiesBaP/
qThIcdV8J+GC44dEBTqSY8A2ikQl1XisKCaTgsf9BAkunLNtTCxEF8Aml998mX/5KXMlXoc848wH
+SexDTQDVJL4X9PVss/wqXebwSxiinkZW0FDXUol0b7caPGWAuYyfTZv6bpFPoVJxVHL5Qnp2lhU
6rjUlKObF5g5ptJfrxcglzA23RzxiZsr2jvxKFqgUZdz+SxFgISRBtYWl95sjMld16ooxeDRUK1u
VerUin6nvJfCsu9b0nlgnrbzrbEr3iAS7aqkI1h7/Om2+AlHrKkx5t/eFe6fJdO+FamYFyOb1wk+
o14WOSome/ruxaeP3OpbNEXaJ0DXGKh8JBkD/aDuanzbVV+3+0YSPkX6vLzu6DMbHrgrpUXtPJ7g
YkX8gkEeN0qTnejgNNJpSykhht2K8xZAYVjuho0RWk/1ISlM0byeyGyZ8Yjc4ul7/80tiiLROhmD
mY2SGnhd3lqK42Npvlx/fQ4+nwFM+IKaONhiZisH5n4qJQUajEwOsthhEzhSooLYpdu4reTY2Ozi
0yqHk4UocHv1XTR1psfip4B6aqjEPmlYVCgDt3wAMn+W99gw4ra8UtCpYINKQWGs/55ChPAN/5ob
iKC6JhzgvtqsR0C/gLckdZs+1l09jjYGGoOkQY/CmlgoElIFBLWvaC7DNlC7Xoa1Kuam/j52TcFS
O5YxwVstdAvZGuwSDemQJPkwQcefXhcMssmHT2LcNn17AcOSMznBli/tUN1Q8EQtC6vViJG2y0x/
0JgRUN2FT4liv70uCtr4kEnq9O9/KXtyjahcf/jlV/agoSah5SBsQ20Ex8Wu8WithjMGMy+waHND
SZE2xI/j2z2uUgRXl3+mlnX8L5TlC1PKjooXO7Dn0n7cCkrltw718uiRDmIkrpm4jcZAg2y0wENx
fzOfuaAKnSolUP3bx7e7qTrv+m6Le/4qUi3oTXF8DZUvPfQQBQtRE1CHaio46ylJ9kWMo6mlV5HN
YOdfxyPgrosOdS9LXlf1mMxHK5qqSJIowru6TisrUeArcDKuhOowoGe7t+BGiIBixsHnVKiCD4zO
sZgJ5RKE2Lmw0NRZUQF/3F5Bpt2QKePgBosRc2JlpigY3ee+nBUgLgW4lV4mnO03y20tRHffT3fD
YVOhrO3yDCr+YW0nRREjfHFoxwf5GUIhN4riKGna5PFBr6BmAJKuVA74LzpbWPWEKbdHzfHn31WL
m9bFCz852JPnH2k1sBAfPPNPvOYxeun8FpoB59o70iUZ5kc+pYw/h+htweN/Hz8f6lFeVpCrMyvY
mG8TlhD43THQ/hMtBw3Nm1CtsnlPMAl/wUlzPVkb7DyEDchzTjWExzccCgI7UDC55VduIuaBncAQ
laISjHWk3fup6d+93NYctQuL8IOfL5XrEI7Uu9cB+dZ8ZavRAZEQBsHXnM26P0CQQeG1bmWHlD7/
/BvQiSwfauVfTqdH+dOgV4xFRag25ia83VXlsBmDv4kj0ORAnVBtkVK5/hSHYWQlAF2P+1ES8hFF
sszuhx+QZ3XnoPSlsvWR/ChHQlWUhBVb+zso/yAAcxfmcaef2a2hB6j6UN7ONj0SuEkmq9MfZ7YT
JmU0BTgda0VBInW/RZfmIZY/AoRR/GdAmIN4vHVDTovpusPPXfJqa+qnMu9IO4mbuIIYLckI8Y3+
F6SV2E43NUJ4Nl3D5gZDA8+PvXQXdxI1oftAds5QrPK5f4JHXtui64KOnq8OPrYNVqB12ik8o5pL
S8DuM4sxHXyrSgDd2HkADmxcDoVYlZGGM0ErFZ0NlVR1dKFssSxttdlGmrf1G7NBLJHGloF/8Jvo
j5EZNB/FP2uXu9B/aV81a7RHqlrdwWN+MeHkrUa8gwINIGxep3tkN8cIZDFdgOXZS+kVs6tbJrdJ
/AItITfuxrP+TEtQCOqEE4uEeAnLP9aXcHuWihq3zCik55vk7c8vnB2oDv3CVALFRW5/9Ugxda5T
UrIYMUysroTMnlKpcsbDdS5ZQoYwYv+UlhNwuDhx5UrqeW4rNebNYzi8zXq368S3pw8IYVTl96vI
NeyR70xjWFVul1IKH3RdiEeirGMpV7JsKCw1NU3Yj13WlLJWOrwRTm6/7MAdDVhsZfMaLRreBO+n
W/gvLq7cHp2+71K2afNtiF0hpAldw4+Kzh09Wia4FUfg+7/xBZxyzPq2VeSSUNVfsFGyhSqEaPho
oSQ31bWI1zz055kvLXjgvE9nNEhgOilmmYexIFiLyrBzzBW6qeUpX4h0PYm+W8xOIPzscF1Chp0e
1fTIhdrNm3vvTmbIk06MO0tV/f8cMcm47nDSPZyiEwiNw+oz9AsPLJJ8sCXvxnPC9qOTZG3+Dmzo
8zOq3IvK46wK3jzueivdll5+qguMSSHZcbYf8+RMWy7mk7pzixPgc/XTvLQzqi4/FNn2ibvTwNqQ
R/g/WINdC7LLNIFQlkiYAKZ5uS62Yb7mcWDhkOaWsPcPXjSZZtmo60uVYmYqf3wtnArTEGkIUA5N
8VJTE58u9Ec1nS8vT6nbJX64SFGbH0gZ0WZSoAjA+CsrD/DgjUcxu1Xbr7boSYT078vAyf6bwOWu
mbBpW9v9dl4zJcOZvcRo9F/+0ZjdiOdkZZr+shMvLr9FO0P9Km9h/r8OEJ+wwiJUGcMrhOsku09d
nsZCEYSQt7c9uiUOn/Am883I5/uIg42w5vgcWHZFX/GpKKeycwXp5f1Hjq12g2itOCWpu9n1M9pi
cR/sTkgGABII0xUcwEa045O6UQmZ5HeHl8rG9i5u1cvpdNbIF9tDx7Nyzk5fUiQJSyZmBNAk1Jfo
wOzn35/8IQYDMimYCZIcTdNE834n7YU4YXEe7FtGO2GF9jWswEDEIF7kVIPgNrEOPtIaUZ6NXjkF
47TQhKxe/kZ67AVY3gtG2t/mKXJUaXMAp9KybVePeF15galpUeYzcouG1LPNvaC6dOdgrUytU9NQ
P4zsjgwr9EVYFg8p5I5z7GFGP+pYfe4v50ZGtnYa2+0+4ZQcRmuVruC7aWe40LqMcPfdCCp6LrvB
Rhh5x6lthF9sZvU/mH3LIegkDOk9uMd9ce9AwewWmZp5jS0aBB4pvczh/qnlDDr2m+v3Y0Kv+ZF0
HnFZOlx88duXyrcYTFczgfLWuL/xLUU8rl/baq+VJRIv67fqtyg9Ck9Wa+wAvK51zfk1xx5FFk7v
GytEIODIt94ZXXkmnM9Pp3NIqzLD4QW3wp9NjfIswZ4gr7iswo7R+9/Xuc1d2BZpYG8RcCkvSUfA
0pVBb0Vhf3ZbjTX4au73qS9SXfF/S231IYBAo4pbjCj00JOAOVS6q1I29BgcJodU7SVPxqm5Q+cx
+wX94RZ8OJzIsfomrUDDrs0wgVTp+9FXwpxEE8JBIIbbJEWA1/xquKmUPOhTD+dgk8KHBEnHszpA
W4GbVmpPLYOA9+fNeHbMUFPXY62XbH5FQGs4GN9JDjkcEqmnoMbLB8cp5SuasgbdzJvYE3bQDFUK
0hB2xNYFR+hcKcUJ19H0r4jjqcz5oD0HkH7Rj2LqafS110L0FeqCOnD6lcB7iU8nuGyDh4dFcLl1
UPG3jfpG5Fgm9B8hvd9/CNrAsJOEIijHxP39slV5XqSXIF8W7VI39Yyt1hdzyRWZxIWhJI7XE+XO
GGLaRKkHV9nMLCqn5QJgvfPZ28ccgUkNp/hkp6Vmt70YnTxOwBZ7XlxRyoIj6s2Pyhx5GvUgJRyQ
GpDPyR9+2/kbrGxBzhYUao6RHwGtDt4mzzopc77HJ9K37KLeZdgc9MQ49Pqh1r39CU9ui9607W/l
r+tJWJ6G8+xx+YB0sH2oTnBF+7skeoYA0qsh65eQw0UJsQdBEe+EZWdmY4+hL8EwRdPvaJcwWLiv
SmgqDhlejGyzQRDnnvn0jMMbUZBwX6AIrYHv/esWmdQR5ikzGVDANvwGLlbs8+rSJhjDVpxrTv9Z
eAOeIVuX0lKmqdbALUISsGTkz3chialYODnLKaHwLpG33BsDwjvCi8QRJRLajIqYOtl/zHRg1wBJ
pve0Je+NgFkaD5Qcyu6JQrf3Ax8so5xGWVtf19QujSW8+KaTHYkEk+Rjc9Li0Xl7KMU9xYKidbw3
RA1W6NVhbgit8wKYl1ERTyRdnm+4BdzbjHwuvP/yAaxZL0qkpoOskPeIDnlpEoH7scb3R0nL1ZyY
djObAYzQpx8AHgYiPlfElZv1WnVePoDxI4rUqMnbadM92K/UW/Jey7mxuTeMz+Tf9dcgWzfr7JWo
MiDBI/yjTxyIMziDCVjGX4yYGMIpNIRbLnswUjXJ9gRHGc5nakHYa2GIwUxZywo6/Ti5W/KW6m27
CVBmZcUjuGHz5y9GvOyUKfqiMwm1nGID+8Pn0G2ZOG2Kp/FjTMrtTSTQykwskr8FjSonF81clXZ6
R170k07xd9ru4yqtOFJI81nsb2DTPG3VkjBHyFfYTNV6D8Zq2xlkyqSCKifd7JpcVSJEPn/FJfYp
HIdqX6Jav3a4bXnISqxEZanXe0Gm2tNEga7IOcE/GAGJDkV+8oFkmX289KBQ6tUtW/kxoeKISYKv
Do/7WA1DCyA9vU7XiSn6YcdIUFVL/4MFmV7UjxIwp2pa42XYe0/EAEnX4mx5Sw4qn9J6zMZEIjUm
43cwX4/Dd5qsW6bBFXJg2OwklaiZUx1Za8wJ4h6iIKrWL7etyssJRzg2lWaKTVqqmaitE3DkcrR7
Tleu7/Wlf1HSWUSR1fqFq05IOfq4TdYqmYqo2X6ZoOdWFw//ovuVBN64zMdhIaPqUl6VcEVoBKVV
brSScF1sbVJzDUaAflfsHQPz562MBe0eldJLAndhIGZfCQd+nOg8Actec80BWN8zN5WB/aHkVSCs
a1SwKMGEQY7h/UW7Cgt3f2D/TAAehVSGtno2u584sXnS/Y9+7pk2MoBL0JCAuNlfPgZf92bSr9eO
3S1lGy7JIu1iGaackomBcLVcjFURY8vhSo1Qqsw6xxPvtMqMGexMkPfK5UE+G97D+zn+V5FCWMko
NpEHD2tmLKGUxTSd1TQ3zPyerax751U6PfQMLCgSU+AOUp7HwBUM/h5nOc09Fn+ZG1R4vNc0C0VY
2qFADoMQ3H3/rkQuZZwinwqbYwVlfH9bfrt60zB+zMbsBeEzU3qbGYe+1yspgktPtUz/YruLRrE7
2ME1wZfFJs1SyYyMW8O9bRkhedeedDf4HVX19k9hdVqONjey7zR71fE2Rfnq3w0Nhyi06UgOxCwC
sNAe6lesSSnpCCUjCCR4WqBP9NbTllNE29T0wTZ4XmYINPaD1PD8O1xsMUs3/EGFZiuyBzgCIFG2
KmWzgrIKr3NaAyzX9vDdYf3OMxXfQNWoJQj6GJ36jtZixLLrnagsK22k5F+zk3S0mc6TxJap9/KV
52PPj8tw23aEeODpdPToh+NTI0l5K0mvXRgRLlpFrUGdr4LifforBv0dwh10xqae+BHIjGTd+dNm
HMBJw6/IenrnBLsbjwqmEGMtbxZdC8kzrO8UoyXlpTlecmd1RhXlu2tnu+dQqb4kOUVp/Tffz6d+
tGgJzVr6LceE3YhU/XWDosSlIb+sbeeFez+MwyZqhfXnzC0YecvZ00bw69ZXLuxu1w9F1SEdofzM
QWgfSIQXaImq8rgLA1+6tzrHksdmZiAkXwwx9PkDs1IEhwFusAQrCh7zFdTFAB8XiyKVkykx61vH
gYhWllLqdkD3VR8IKQ09gFllmfXx4ntBi6KgHR9XglpYTMf4nOoC0xab9k7/VWj9g7Ji7LQxIksw
D9PqekP/nv5WCjRM2F7pONGaPIGAQJmP2hX/6y/iGf1XN40GBaVFVKjmO+TGJpu/axuGxfAdYAvj
hldxHaBe/+m19C6xSM0StqOfIJ0QE8Ya3x+KpyJzg2MERaRP3fBBgotdN4R+wjH5DtK7Y6cOwh5y
M1nkq8hewU2F8ui+Nng6F2Z1F/U+e5HD/nrRjmbylBgh+vq+2cPO6OotDyU13JbrVdhBAuqu88ms
iGJ6F7zH0dXyi5r5Z339dVf7AkYNroWn3RQUhe9XAkmSRp6ElOyypNe0hzyW8YdFl3zuUR8kSCpE
2kOzL9zw7KdsjCD4UutvnKgnC3e9p7bYteVUIC+L4yuvsaow1L2pVUYFxi2l3FfYC62BsrLqcFoq
DDMuXC8jozChBVqMD4YyyX2AgwM3OqsftsARkKnIbiaGv8sqt0FfTv3ufl3i9tRvHQL13LPRPle5
lWlVHt/gt0juQj2hPpX+r5gVh8ytVP32wni5o96k4zxy+NcICGg26TtrK+25naTn4XeWIOjyKEVS
06vBRb+gugOrA++xubmU2WbP5z9Pe6qWaEILl4wn3xqNBRtvW1i5+fyQJmIaZyKdu2zoxlabCImH
NIpmAbfFquwksevMIzLXtd4cEcw1EE+5/Q4Z/lGggcM+fYemRts9MX7L+Med5OdjVkzPC3sc2puy
BN2fb/rwl+rHelB3sPfgmj1XgkPpjwOjZ2BCc5ETaGZ3KOIBdOUIqdYpofbkTvk8DL8s0BCPoCEs
GacIeZTLzHe7KlW3PSShDpxtk+Ji8Dq2jvBJ9F69vh3SxyEO2PZGCGNPnDfUESnwWWToytBInuz9
woYncgYFegQdvtm3EzPiWsB+RWeEIiVarJTfPZ33pA1AQchxjQDVKmFMH5tT6S4WUbTeFazfpX7H
oGc+buZf58hOAcLwE3tGvg1YovPA5vZ63hOovCbQMkiEyK0wbkmq0zRZEvGZ6VDzWmwv5flKv2b4
u7ukVXZUW4sjDt3WRLapbDNmkkbi04I+FGGUNF4Ub6Jz8DsBSuBdzsrCwuGsfI3QlLmhfk6SRGMU
9nhWfB6LlAE+ePrgRQhfkqlP+3BDcCZj8uFgGWF70d0z88zkVt7vBovw8gyDAYEbyxGwSmBHlTzG
/TfAYljloGOqbTCPEVrtUHi35NdyGnkcpCDjK1eq9vHQnX87vaZGhJk2249pQ91pkel4t7ustonG
V4p9VTB4yV2gCOe59wf7uG9gNTqVsqMrsVPi/z7aa/iUmVT0Oo6xuDATbjC3cADHQYKt9NGlij8G
UjBL91MFrSdFz/sojfUuFOJNYf12d6QB27NtgqtsJU6nxE57tKw0VsHTTgLqzdkpxinNjQ7E4Vsz
rW1e0Sv7h0Vg8g2v4SNJefMAoqZS5A73xigZ2aRfVWQsvOKT13p40ozznCU7KkhlrPfEr25dZRGM
t0eFjkTvalxWCI2oPs6qgdtwTf/oZ8lyBQ8He8w2lqz6eEOkMK7fN9AcPzKfKL6Qx8Lf0RfJrXFd
fx18yk5mDuILyEx8ffrVwbFh+roOGHgBnDOw+mcJKtQWjYSM+/z2wakCKZFke9lHpmiHO73uTcPK
sOf62Av+o3n7mvtcRyt6NcezIr11Q2lAQd4CF53Pb9BaikFjP9iMZzoi3vNTETH1twrXFURETE/V
qQbBq4kKko8lXFZjoTirGLFssJEF4HjssSt+wQusOZWhWo8uql0K1ndN2aXV7cp2YkEeKf8KUk0h
xbTzxWdjgGCrlfpyhBJnsLWDn7X8xfPuODNEQlJDaGP3ueVY8c489UmRmVojDtyKyYwNi/5GtG+w
UrW8TnMvUaEHuyJaCssMJpzDY22+Gnp/6LMjT3sCWsSzPbj5KSuo9OCNvq3GXP/Iupjmy9VIi7ie
t2VW3J27db2Sioz0LbYkbwzW5By5NBJDuc+WnyQlbiW4D4BqCADg8W8XtoRaEVog15NVFlI0Uf1x
+u3xbQwiAUpMREJRoWaurTSGv2esqSYQMBkJR22eL/N1soHYeo+riE67VNUir8mYbYdDvmPkl/5c
hJnRQdtHlYZaG8m5WslDr/sJlpw2rnEWtG8vKAUiW352qtF90DKypOF+QVBHdgxFwhEj5VWgsEY8
UGkEayRqoXIBvTa2sGG+zJG5r0yH63Mga2FIMH20jvn2lwraMwbs3v9VS/KVU1R/GcoSMhtX26b9
R86T05uvuiOM5YPiGWA/NZNUnK1kvE7q4v474GndsOZNDbw0KOF7PsEBLOpqYicPUCDUdkUAvxLM
3ClcDqB78bv2N1oIKnQNdOZCfKT1eI7ZjH4C7EW8oUq0Ke38Qr/oUumv3JFU3/NQAymNED54yBsu
tXzcwhy8J9QaEOYHGCjnx7x+0wv57am3kMadIayfwNL4faXDpbOl+v0OqivrnQo+myp9b6i9aRRJ
cR5q6kaGba8L43mfGxZsVTzxpJoCDruA93MmcDa40GlMngzK+Kcz7KLbhqMYEnX1/9EfU6C+Hw3y
o/Cxob4QDkO3wY9V6096v4asiIT84tvcpNc2QdeUH+LKHu+XEHb2ZVAkfrvjrG4y2fpLVZVS1EOl
3dr8IcuQJtM2+AkfE1CW5jvAaEHQ5MBkvsBBwcmtWuprNyd5vKLGiCsHGnLIqstAdoV/Ri1bX/iD
0sQV+Wb1vS6Ic6OHwE1Ikrq9V7/wvsVT0MHolRtyvG9LSua+yUEnLc5qzvs+y7SzFTQhLgg/RQCW
DTGNX96v+y0Bpsox/MOj3mlw9kQLQWLoDZTXAjQ+FfZb+xVMsOwYeQQn7IJtGTZEKEJHO7QO4BIJ
BDpCoZTkYqHEPGuET9jSdHbunHPn0yHKrI9wqZ+ntmIc7JYgg2huiUuQgy3e1eqYUPsVwVBNjF9o
jAKFTE3ocwqX8tQdvvx5sOoe9CZTyRQfFyrOywjr7dYJyfSp7dmFvtvehxpypMywILlo5kONoQ8r
Rg5kR5z1rFq2V10ThNHYWmBt2H6gHBmaAzOZQaVk63njQQklNfQImLWjLqMrrC2yGw8fDeCoANMk
kSIRGRqJ3ExaRSJ6d1Sf4R9fUAvhBLkT8V2VgAziQFXsNIexwMMqztjA3e2fb1brDu1tn+M71ONr
VMdmE1DMHDjqtg99WH/qrH2TnFc03BD/VeoR3RCL2R3Kupacb+/Hc0nibtzETiZdlhMHcwXSMQpt
uD6K1qhG0g14PyxzJQdmkezfOKmskRML+iRD29SCdTWf/CQA301gCSwCYY5In2vS9fUAJ0xEG8OZ
a81thEfpcw+lOPYhWkAQ5xt9NiXBBkhcfRlNdLtUayuhHV4V+WP0vjyo/+my40ecApHEpJYUJqHF
IXYcxa73N9qtvnPfAAJHb7RpnmFtSlmwyf1o7uYXdEhV+4VhXpEwUDU68j3lLzeIDaHBRSpOus73
0pgglB29tev7jOpQZNu8OaDgv0qQcGomwPCQ0zfzVDopi3oR9edqqTWfHpDdmJQDSQc8C3Y6o1+B
ATW2LXyCLvpragTYBK7rYT53oXJtGetKjvGNNW1qgLlCyBg09rcQBUcS53Dy5jQLp0hjfahREnUu
WzYkoVC47W4ddYfeSJLZ+jOj22MlpMxMoZe75OGHA9C00LZvaduEXVdgcghd+c46R5wf87zk0GXY
iPcoXcQusFo59W2TXwx0hSwDcZngswrDx90XQbpUksoZHii5kAg/CDd2QI4dStwgluKcN2yXljAe
QGCuEJVrYcLlhJgdciSbCj60VXo09ivkVZuuQ17Kx2UVEeSLUMwd0YDcOqvwRQgKVhIYfxEDR3+r
gdHs9zRb+Gea9ORx0NFiG+l2wrwYy7WvGRkjbkXl2dyjNIxe3G8v4d/Cu3777xV/pvCMq1VxVPj7
5oAcKmAQt9cjka9z+AxrQtQ5X6iOq24iOFLB/Ef/7CMg1gYnmJyGsxxQID45mUx2wCMr/kVj2XpQ
xNm2e73NWVQeHIhQHIQW/9/jnLOGLSrkOOOlwJ0hs0rKk+PTazfZz7UoID4mbERvKwhA5KKQEZi/
q7s88OHV1mEUHTtFAb76cKpaJsUPo8iwnSXkm+eDtGwsGfbdEN03K1LFDs883x9tfCkTHhDoAVgn
jz3FJMaG5ZiU9seuU9aK61rWvVTi178eCcWRoYe4sxxCHZ3NtjIHzM07LVWq50F4xURIcjrHGmsV
Y5hJN+fESa9gmd6/vTwqsblTXtx/MbI+YOMsHyHiVtqLql9HBhRZ7XDIvVP4g6WAHukQcpLqYXso
ZPt12jFiKt1Z/5n+A6t5lHkq3jsCCg3p+f+IAWE4ULEncsGgCCkG5K1Y+w0dWfuYYvHh7Py2ptpm
rDUGt2AhhhI+qWe48TjtJ3mu5WnCY5tFQyshM6VsW6hrcXXbTs/3uzA6ALRWiO5TUTlf6NPJZe7q
QT3mc46egf4Nl0jMeCRnK8gTPGYoscNqMUGqNj9oNfkq6wjodYh7hjpLfxVh5GOxLQ5xTZBfhoC6
nGtjGZfPtzQrwUchBHbcXtRM/wZ8KKP/k2Q5SaWTvBOVAeJSp1lYkdE/mCik/ZyVTKJreOR2S1Dc
ibRy/8eluRS9sKjEGdpDLVXlC1iQGHA154dVKBxZ6DJ+1DkpsBnpvKZdJFVRKxYfL3PPz1YUqLII
dhinl415P7GM94XV+TZfulvaKFbaGPBqYvLDTCbAX3FyQLek2HTlD+LFC0Bx61LX5q1bPXKrhyxW
7eldCE9nzQbISKNOn+pDJF+0RpujBMO8ohqhZDhQjQ9KtuHnhtEuplEQdOmdl+LqvuXcZW+al7ee
OnPcQXCKCiDlDEfAXJz1nP7jlp0MFEHQX/P02+7ZUoVpQ5ty1tDBa56QzTaRuEXSblFgfmT80I7j
9u+0RDsF7/oGWbPIwKmvBow2iNk9M/q50WHCGhOZibG1TakB6g+cL9erGargUABRvcPh6UbTAM+G
iEHScfEjXcGHvLZCrHKQndiDGZ3145qV0WU4lfQVGBJR/e7k/6jdWNRbik7OFR+fNHU8rlPT1E9Y
fEkNM0NY63QVJVsz6GZH0zADmmLVXGo8ZqXaBFd+ykfwthCCiRMjNQ2JtfGhUK5ioOeZJ3I8YVbq
fBRnKXGeEvzKrtoiDT2Zj7KNKRGpAORUxenQtAN/AhF/nNaukhcxH0Vnb+mnSJ7SvJqH7yyV0BDs
6XE5y0nK3sF2GljOyQtn/MQNLoZ49wyGh8z5uCX9uIb/IpZHUwld+9THZff+ckAcOy0shh+HAqPl
vYQsQyeHtUR7Ll0Bjt9xkyjPkQO5Y3UEzlIxw5epKT1oSG4sdVErpcVb4P7dui7QAtFbO7Yhlgy8
TxQp1PuQj1hKRYrI1GP+SeogNvpQ/NWqscSn7eIicce+WxGY4JGxdOpFG96iscSzrjZbMc/ZkW4b
F2ykfklUWycf93Aq0iKZuUkkvcxmUGUe61vu0ByGau7JHnDc6ndfe//FImuKn+ft3TT8E3Sv+F73
y5BjEWU1sb4FqygPvH0ipKPWtfcnSa4IfoLo9Km8gIxjUBXKBb/z2PvVgQhTnAyKiT7nRoi6DhJl
K/uoflliQ4VuII9AS4oufGddWBYPS7VDX85XEPh6uvyP7R9ZoLjkkslbdOAFpFerX/Mskl5xz7zB
aXCN2Gfv622hqutAwHojPiR+sJDckX5p6A7p6aNfqbPXSIgWunCsjAe5LfFbaw1MvV7S3LE9eKX0
m5cM6y9cqLDB13eN/B3rm7aKvTkHwfMSLYyE3BoIk3oMQMTv9BcO5GZiclPjkN27rwy+GCIchwoP
HGw3FUYAd7jQJKwgTM7H38kzvOnXlYR2brbSXulCAydAa3bJ1eT/0wt6GCfPulPUFry1heBuGNOK
WljQu23eGGKK5DSHmKmjvZENoiTd4xavs9AnovPP0GuM0n1WzrpiHoGFcgXIRuEyg8tNxYEB7Y6N
M82aQ5P75WSrJviGaw7mdEer9qn1bPMWvDEWuCXZzLxFN2jvMtsoNTWMVow5n3f9E0NawLvCCMPy
DNYt+sXFqyAW7eX8IUJO/VTwirlZl1BRCB6lOPXGAj0NdkZ8Kto/gV/8SqkONQGnZydANwxjYmLg
0YyL9PZBgsmdrr2BnqjIF0lnjJSTNOXYlT1z/vULVwEYGaqTKZkgb55665O7dKA35AE1EXV6U/nn
K6WZpbjA+DA1GeF3G4TQZrJHtNZg9zFNyK7JS2kH6Pmunq4ahK2oEKHTizJ4fr8HelSbAKGelioY
4kcv9cr+26kgDMjAWSNaQU0x0KMTjT1CwMkbu7Ml6D1MjkkPiWqC+CBJe2O5rWWITflMmqcswv6c
KI4wXSTz/kkwD9M0vDaCtyrmXVbZ3LZ5IuL9G2WNQMHKmfg7/NryyPH0fXfhtLVkbV2yskUIPsBp
YSUaoPezx0tTv0QYqXd3CFshXLBTFGeji9cQoO0s/gHepoPDsu9VhVLvK8Z7ApTDpSkJ/7vKOmmR
uGHvoc+hjX/i3J8Uote66fT6/WP5RTjXTZeGj1Zzegx7IjvueWsJFbTxMzN7COQW70/fB4wS7fZr
yednqcAHmVRuH+GDG2WGusHO43CVlZzvmWKONgK4YMgk8cuqmSYBTBueeuUqh5HhSbShAFHZ2pnJ
IkObiaQpU3q1sz9zb/xK7yvJRcMNFWTxQJDsBK9phvbOci36o7hZBYrJoMhHDvWMW1xoDoZ73egf
p5a4N6YnzdbSy5+vPC1+1wnuSX58cUQ6KrPqy3oJcnshtFpWrY3p7W6/SOgJHzjwmvJqoIhjR22u
IxqidvA3pziic8Rf9BVH+4I0Sedcz+yijxJbOgDag5CKTbBr3ZTWwUjn00kt7rPZWnf7w6rmQ0VG
N4kQqAyfwkQvxO40+7DmpXbhDMtHeJmecgYLJAMC/VcIAYmgbVLjHaak4PP8BR5+bnFXYa92eK9c
kYTOHGEJboOOB21MZ5gRpyi7kP3jv9Or1JlD/mxGeR5l/Z3v0GXE+KLJ9InzjV6YWIN9KOH6g1J2
qhjNfPcWwvvXX7AzDK+MK22w8S3lT9O8W4zI/lUycLnHlCAi84cZXZpfIFymntSng+57hy202tNi
aKAfp6et5/fWYo8wjCrvcmTaL+8kqt9pRVtRZLldsizoDmpAGualMl8awUdlrj7W2JsAnlk5tOa+
TNwLRX2UKlgPXsoZm4ktrF5P9s4U6t7yXCjsxPqWybLJ8ylsseqTrepHDsVOWpyx8IIq91ozJU4Y
05qhgku13YArD0stgO+OoWd3Xn6ZhRGenpptXXo9WiLSrGu4yqBE7BMsFj4oEOKtcrOb1Lq6Lqzp
QZQhPZUiAQumR8cNH1Vo4zgsinbAu94nzbqGP2BoMM87gxJPUh/JLmW/M8t5mlYCwKjR5oWlt8/f
qi2+mUXXqllNsfnk2vLd5gOdUjtve2MmfbwBzV26Rdt8Armi+cBz8006BnB/jXtrXAl+XQZIvkgV
2MDE32vDXxAFvZqsMC7CLQYivapIbA8NlnQjlRKv8wdLfdsjRZwu14igguIN3oN+IGAYVhch9wZ1
NADeVqzpWjJTvpHMzsezL8AqWNOaO7T4jQN/e/2ZjixCKtjJFUp0bZ1GrhAddMzSYpAcSlMXWx9U
kiGMWJwVISsYMvR5Or8EUubJ21wIybqu88u2D3XQBq/PuQqDInkTyeFeeUfv5bQaL0EFsCmipbMR
pFJSc7Rjc9gEKjGHtuLyi4/veYRM0IxpErjH5/4EsxezTc9fSKqoE2Zc2meEIDorefnSyDD9hczp
k9g3EQvj97DrqFCTGVioRbd4lBNxgq3YylkJsJ+SiGYSIWtrP5ovr89icjqE4t76V4yZeDXtvUTM
HqBti2J12ccS3amylrb4ZyG2+Wjm6tPvtazHJH8SXvs7u/ANwL5GV18inXrpuRC1EOd81TsPuNEe
rx7SF4Wd4QKgugt4I3c6XxthH0iAmKfC9JieFWENuKBXQ730BAsxu9lSFtDAYYPra6CUg4B7TbSQ
MrQ5qt+1tHS+k0rHIDB0k+TAxEj/GZ16YQiGjQFAOh6kFE+LXTwhjuk4krr68wcs2Z2lCMQE0JDb
PLub77a46iFc+lXng88A2TAK12AuDdlJAeXk51ta15h50BnSYRBgZVy7O5UN7Tb1H9g+44Mu7hLR
hKHxrpQsl9JHoQASu/VBKS0yroo+DvTzX2zfdh7A7kG1r/kXV2Ti/bHhK/HiU7khMd7BXEfnA/15
seydeMiaGnCCsPaM8xwryfU2h6vjnHnyA6bjmpDJgCEiU+dYQfU2isWXMFEe8JiH8sBna2sp77Rj
81hkReHjbZdIxJjmueKDkVhtGV9TjCAtfWUGvp4fgJgn4E2F/+9SPDah+260TXUF+qxNSh/ZkfSt
kzna+5NIhuCEM1n/70H6Ud222RfnEw9LiOtYe4cGv4qpGMM9//JDIDRspTTpRy/d4DmoAv28543a
VZsmyR6rVTMuebCSA+SOXuhjCWyFs/69anFhv6zGuzRh3aHW998Mgoweqp4HJR7sKN1yi0Ku8T8o
RK8MtbELBtn3cz9Rax+85deCMNeKtcGKTiJSVOhC1HeIjoQEVk3sO1o0lFVG52nQchst6ub995dB
xzdB3oZUxh+gvORHUe4aj8vvBu+9L4N+9Q3vQ9MRahj2sKdQ5JUP/3vEiYeUewj6chuXWM6sY0uO
FPG2OCYHCx9o8biy7FMIaPDVmBCHFEoyd9L40D7zbt5xo4YsTrlih4z4c728J7ZJNE81wHPXcGyt
kmZakVREFeIoIPVsuFlSXxT95efKZAP5BgILlS2VWuAqiD/nqm019w/jIf5CRHxc4mVS//pKQqVx
LPrROjU44xJCKCz3h3b9hpod+CnUejHm2X8G8D1F0V9mWEI2ho8odfy8KCiY6zrpjSTD6Mc1TTld
P+Jt3XLxTylH2A0jEGpPc6Nn/gJSnGSv5jMILAomO0PjbLYFenjsA4ZRDasdKu3dcpCHo4x0bggH
dgRB0Mt2UrJg9adp8s2pJvHHt/zMOeVMLxZv6yj0HVEjdUhtfO65fURKKNzfHfr6ajCRr81IH46j
TIcdYNwG9kIpDS8BSMXZDsTr5xQVLMVq2KAURnllvr1lquW3TRO6YcDJg48jLwCFEG2OF2hRHRjP
A4vqPvTDCcxTuHvE/aTLW4EokuhWOGz6kuWIwgTeZ2cXIZmqxpgSOl5VixD0SgufArgJyfG5TxbH
Ev6sWKQo0iwbYn8dqLZ8EZZjlaPSIZFhckKbA0PacAReIcwE1e9BsCYFEt9UX78Ibs+RmQln1CNc
fhreYQmzKcxGhPYZbML4bCJ8TH2uzR1pfkieVFNe/4kF5P7/Ui5tbYRAgvNXWnBXYg3C/hzLwwcJ
UFn8NEqIE77Gkll36MntulVxTyEsf1F6EyBlLSLwMbQPrxSnhl3wD9j0yM5QFjx5QD5maKJ54gul
SSi/rQridRWmmvciHPyg32ZU2l7GzQ5eDgQRXBfpx39ippm93yewhAyTBCaRmm27hJq829TAKrRa
c3mF+QIHcAgp7FeGGadzn5Ep/38rx7FlwLjXwtGY/pLk/xAzu8o9xXNlVXnvIk9Og/OqDPyVI8J4
b2gG61aXEvK4vo3K2XvQc2P5O47VqdnTkCM8AOUasrhmUIvgeJhxKswDoPej4i2SxZMHBkmBHQy1
HODbBnRl/Cpq/uMmeFF2XGAmgJ8iTaFoRE+5/BVpxbJe5TxSDjyQYPfRWRgfHGuyNLw2QhFJgr0R
fUafA3ckmKh0YwJI0DZZskxPq4zZYSaKLngrA6hOWfqi78ns9imzkhhtaup3mcNlKbILkQAOKEw9
nl/ptvOgpmr4CtfWGPxSDQ38Er/plkakYtrFTyigoqUajmr0jJ6Q/RQLVAuQVBZmP7vIP4O6tbYe
qhjt+ValZ6W/UBIlSyIgkMXAijeSodvyF51Am9Rc/a+W2CgvuYuam/FBMmOVbrrzi5iCSVh5yde6
kMry6FR+ItxzCJ2egk5BaQGIrhB7dIL2+R0bSdsLeCxz36vXrFIuqR2U6/0pFH5KCe4EC8c6isx5
MZ+94wA7wA75DNET5BwcmUrGGscBlGl43hwp6aLgo3hsJiF3te9LMmfMM9Si066XbwYyLwrrYH1t
wPyyO5ir74B1aa21cZX7apKjVyNtRKo3OHyY5x2cUm0wIGSoBw1RN/fP7k8WBLcLAz7TUOSG3pxK
HDEjV/Y+CVSFWUgqHrg42s5IZ54jmT1zuDiZ5Coh2Ok6EnM+xnOk4LqavUfK1U+BPQrgRe4qy43r
vn8ib90/Bszin9suH1y2ifcXCpCU5mv3gVtdxyj5ZBIcqh8ATuWLPv8vgW2pguVQxfjJr6uBNgv7
jFb9wXhFSRZnGoY5SG6jhgI6oDxIvVUzARTrtq5PdgUvi7hs/NWiAANtbPANZKknMb7juBuiL4hN
TLC458hygbLdhT+rgM51w8QpJTiOoNVihinVGv2Gt9PacqqTYwuKS2L8nWheX5+NGZytCqId8heh
hj+Thhs3BdNGwGnir08xFI5Ktb2oCjebY0F7GdFX9EMxGAO+L5SkNv3iXpQNW7ritC7kS7T4L/yc
Dl5ch3EuEMbTJE4hmbG+s1MUzhpxyvhLlFRTA6oCRguSAtz7a2163ZvfeIDpRxHJ1wPlu19hBn7E
db716ztiNrehp9CsXjGaHIuwiTjWyYVaYTh9lVTqdjZg2wQiosEAzM/gg9y78htqmJ9La7CzogHC
xaT2J4xp9y2byncI8NXPAHCVg+NfMSHAJ5bCUv6ldrZdFfgNpaNgjwS3Gi3ySanIs/Lx2b7/3cbD
OtjPePTuyqNcEGuc3zciqWo1qbb2Arul4lxMLa8RmryUP1p0OZgbwEmjaw5bWEiDeKhWVn7pCMmB
f7y24ktAS1cQiIxTV/HiDTmNKyubfQm+eRXoEFkBP6j9pQ0fOINdZwkGynHdqz/Et84vrEqfF1Ip
yTmgi48JLkHbttCW49MTjvR5dR9DdPWKtDU4QweYiMPNoPvFHoF0rCSRSq1Qctu+kbRArAAH+Iad
MPPz+o120cSV1UcTlwh+BmLMIw/Vfutoubqg9xfs9tLvbaQE6fnt4E/mJFh61N707nBpTH0k9x//
08X21I/jYH2QKUQccIJ3/L3XZP0oE0osAUgMBUPOrZxFDJZn9Al+xyK/UlGXohpmOfukv0Nhi6wM
kI4xrDmEavrfeP+mDgHKO7U5mZioa8f/YqnaWEAvZnnq5ePuRbZGfKY4K1Cn2R0GmYRVzRHwOoQE
07KLjOTMnSUALolTu4B+NGD//nSfDq7OSti0bhzOtvZHpqDUy3epJAKRaQIAwNCssrH/YxayCIKv
HVIG9fZtgUIOkwdbTjhZH4swq8/wafzUa5hk58meTpNDlih6Je0AlqSyKysLpIyJRenWvq/cPQX+
nZRd+xvt2DEZvGpm7mkDyWi4hm4pNavU3XKjvqQ31V4kUNV5Dv7l2zAOwFh+KW+/E9K2oXuAAJBX
TlSBNKVODlm6LN1ymVquP0AkbD5afCInPzBdNTffH2e6XABRU+eXcesYfklOZQegpNxeYtl6F0cb
iI4utmSrhgYNhqij0WLKpb9hf3oR8vAmiazjZBEY2pm3x1TAa+RpEcUVDy3DyzgvCdMx/AFHEDHd
9p2gcR8vXpJ62wM0gmUbzIk77Zkp8Mj4tpDhuPUIkFQsHx0gLzH0cgY6z0Yg2K10w7nuPgtVZeEw
GWltCZl5M0ZZ9A9Uj9sBnhKp999sqORSp+vtT+zb50bjP2hsew6tas0vNn+nXE4lZEim3ad+Y0R9
iHtEtEOePW/YSwHnrdhjYHTvTQCZGxOGgFI8azlPa4tXpnFKeNmAgFP+Y4NHeiHdxIRA6knSBJ3Z
PEWiA7QrZDx1q7/sC59yMf7GfjMQEJ2UL02OJKHMk1+8Nf+lY5Of39ij4JiKpNMMdj/qHzGRRv6x
Ta14yi2Rd6c0iYwYrtuSac08MZl965PH/NamS0W0GUXOV3TNfQUnL/jeqpJzFJUQIzY/7eI6FsBr
QPktWZrwew/Je40D1/j+HX9e74LK2kcTg9/nyTSqM+OozoFupHCj7g+0rW0aSTOI/IXmRu/C3FUb
8y4ojRAd55QQy1SpxqALXkywQJVZpz6gn1AfA/hiFCmQrB3cuikP9s4vQYFWcwd8R3/Z5oPPIiRe
kN7G6b8rB1QeawhU11+Di+XBzkLVeNB3og1+7RIYUGnlFnmNx4G9nVndadg10qNtx+C4Z8s0TI32
TZyEh93I4dfIk/bONpH498pEro8dUrK0B92UEQWQt46z59Tctl/ET1oJNsjH9Qwq9hKtSN41qrnp
Hk1004yYBlPtdhpfgvSD4k9EXdVHVKgu3lGP3zOfT5iTIrJjRkfzMBAkviuq35HIhG4vFzaq721Y
T+Yc9wTBwjaMAM1xZ8t0BzkK7M0zxhdnLkxdksOdVN1e+eLSTdlkn7kBbNSMaOD/fEAbsLuJ4Viv
YgglKe7yFADbTnk9YHNeerOjmgOFswWDFBawyfMtIAte/5Nlp0bqHqXXMkwbsmqjISx4LjSPlHnB
X+mgZ4Ij9bPwW2e858WkFlf64dtDK2hrjftyB9047Ennqp5o9PGPoRWFLsq0FkgUfzq6TmVbzBsE
PuKFz8qRno5ZuptWWr84obgvbvX7Z5WBkBNsnbv5vZNzuHozjpPEmj391kZXj3XUbcReSlRJb4rT
06PPAYequWrCN3Xx8AZvpfk6Y2htkPJkvX7vg4SXVscFgUPjLWJJE8XaJP+ydoVK0d8OwVlYLFQf
js/LGDS3U6QNGBZAUVY5eEzZcC9LHqniTah49WHOit1T1ARADh+3/XmZ80w+TvDyh+sNNnB73N9a
+e7pgIL2OAiTBureDFozlQK0LLaIZgtS6xVMode6GiSk9/ws+zu1x3FvAjCI84w+R6nqaheS/CNu
ZLRdeBNXviuTDMSeWkd2q0KMKr76zJ0Rnvm6Kdunl4g8zKGVAYH+GyaIpEILi7F3E6WlaK9ZJ4Kl
OXmcuElO4qQKGmafdQbsGMR48wQgoOP7ERjpoNIfiEH/d08agskFbM789r4Wq0/grfo9yIglEh81
O5d02uo6dYKW97aZQuTwpOH0s1uH5HwpOOiX/Qn4hhqZ7jYOcYLfKddGiwNZ40s0f3pVlv4VSvMw
tNr4GYJjkXMEZjhFTr0XasOXqH1tX3jj9jZoXGuKjcM5rl82VevXM0+IsZ90yc5Y+HbaYKsdFDM2
eIXYOYI4m2WBQ8F+uSzb3eZl6FaGusF1adhhiEc55DIECVQFCIwJEbsDbvKniaozRXokCaBpf/UF
wXAElhbvZ/1nP4kPg//OAfqxFRKD2xsUXVT6WGyQx8WimSG3Sp5Uc/BBM33O+SvX44e9+fFTu38l
OQu9kY/GdZoiCiYFVxAVJmmfM3Q5d5BxuLEdL6mJhwLthlv4C6gh/O7d5pFJmiu1Q/cFjZLMxpzM
/8VHuCnkB0P1NIKstLZQkYNumWm4y3fDRtZrrrkfwYk7m4xKTpLY9k3JCIHm37kwh0eQIBhnthzN
JYqjoPNOsIkfZ2h/bAF+15l1g6KE3V/g69Aj0iQkxclxDdE+QjvGZLaR5CEc0oDtxCjPZsoYkiba
GsxubAX7XVWLmwySw/1GizI2eYdSEmuuGrk5w3dsQ1z3wC8j/KSoT30C7K+lkG/ZWe75mm/IE5pd
cEyeFhcOZ0qiVTxgTUSfDnkGPWZ8mPiNwH8+1qYqGec/CuXV0fIKUioJoUBPsKY5XWWSqs6T9nJo
rVzKZn2One2SlBiB+DmJREQSByfMwMFZhnFw5ulP9ZQR62A1y8Ru60WzknSm7zl8vj5w5QoxgVjk
9r5ytppqU7KLOSl5Jd6CQTIGFTIJiPZplxqIJ9aIwbndeCNsehnLKJ8a2JxR8zIRiGvxn7nH9k30
ukJXWBe8RS92TLjnnEaVMbia8i6Gms0iu4d1pkDBM4dMLckmDj7NrozH/+0vG2ZNyTLEvavT45gp
J8q/cCiISgzBSOoMBc/l/QuucCCBEKoidU9LsN1aBBZqa0xCQmTV3UfZxjEGgFs/2c3ppRqR59UZ
ulyx5rBa8cguHIlYM/I/TMNY0KOJvCX326IyDTb9EliwG3ASpud+WZQ54zpVeNni0kHVHpKoz3kJ
yZHFOb9MV6bZZ0GZVaGj5GuC5N+42iVIIhN32stQkkvoaCTVMgpGTIReBYnp2EodmPbsolLbLaLn
ThewWx+WcC0lPTkL7g4jowt0FXbcwdpE1jEfAPr7+ChDV+iddLxruR1I1Fh0CHSum7o3rESw5qL5
ojkatLa76VSIZRhnrF3BpXur+gzVeABFjB+du4rgy/r/INghVuQlOXxvbwNqsWNeXtLkgTz6Ydoo
JZ5QewFb+9Emi32noHQLdEXDzNae40b8cKgham5scmAZE+z5dstVj453tlfWeW8kYvy9QEJhU4al
LBeiy3zgl5vUKflroc2KbLZZCqgR2PCJNZhVaDPRQJc8Po3Z2EH25YRH4AQFZjk9pxutA2rEHwkV
5rpXeja1tu/H6H4lWjexVtdhUFAXiTnQMivBOiGdIv5T059Qw2Qxs0+B4KxHLCVz5Lwc4ase2QJH
DQ5HsjhJy8ZFll3aFfTQTmvDFfXNtsX27KwHRHSmCm1lxjd6IkSxBpHd+Iv2tUiv+K/w/Fiybzk4
XQ5vQYVGkPkPHaNF4KPvtONzzy1Y1Z3gfuO1lkuj/R2oGc5eV59xdSH4zR08YJ5Ij5XGpPQszvnC
RrRRPExAnSbTYN3Sq2QV38/t/6DeeMHYRgi4wQPE6cnO3f3jsFbEXuObOKdJAksylMvDP65LrrMq
NhRF/VUAuOEpL93qgGt+C3eTN+WkjAJNjo/pdyv2F1wrYUjBWsXn1KTuZGo4pzoxDjLtHk/QwzEu
6oh0ifAxCKMgRQ7IfFwoCd4dfAYvVAmbtOXSvmWg/hrwZ1FqGTJQBi+OvU2+Hm8wqECNaQ7bTUa+
NZF5a/1aveVKD2AP7UBeXDTpYq6ZhYmMIWam86aWzY9gFtBpKNsBl2uSK6wq1tL6lba9O4fu2tNo
7u5Tglt71AWvwjOYOBDHpdtKDhOFYZmENDF3ugi3FCJioHsIKo+3o/6mD85gR/VazqYlCSwYmVhA
Ir562fsWBvjFvCq8ZMn7zowB8EDpLEv+QNgZVlSJixw3/7wd/uED+91jyjak+UiKzQYJUYrQdaIb
yeyrg3iik9UVtUQHL+g+Re72jHrUhJQOGqsWzC/c06HA2hEBblK2ny6oOUEv7Vgabp9WkZQngJvR
ODGIXOgsnCE89Ktne7AfsEsfcnXHtwv7TptJYgXRxy20V4Uqln5IaTGU5whjz4AaeDCdTD8MJN7H
4kAyFAzxN07zTiZou7qrlWaOv6er2GpRkEJGt3ljtOZM+Kzm3Ghvhlntht8DuUUkTXmx8hcoKeDb
VXwr0WCxQt/DiVoK3vFnixVANNPdZ6NPEUDauwJBflIjyVdhaa8+UJ7RkkxDETN5EYY0rinD04pD
g3uSNodzFNuqbK1dGwI6ivm5rD1N6u8YuWJhoFxdGWp+/eoLypNnXlojf7ozfEG6hO9L9QiApvU4
f26TgFzWi3bYlyyC3Siwsd3BU4CwwJaLioUx5+MORFZHxqWjF3OLI+ga6YoeawF1fAA66Gu/TVxP
bZIl3eb7By3Y4aDzWiE4X0YK0n8fIHvp+320fbscjtfsJMdywXwkRQfZ3Ij4ISO5Ce3Im06VRaZ5
cFm/YjnoDfDeWglAh2XSv99yjMx9EUKGRdl7NYrKGOUeJf08ZAikOORe6/dH/7bI4uoRQWaJIWmk
O8Qz3yuCb9Ni7f2IjZivUogXKCqPPSUgcozcDABJOoPqFnC6Ra89ouBQFNDm5mqvWaf4m9yC/LE/
tEZCpGeZ5pCdJoHykFOSwKKMKEgcbuJ39aL6d65Btc/xL161+h6dvX8Q8AjzWY3VXWbktaz05/7/
VCbIgooCXvo+mJ3YtBN0MAxEkcA6PYCAfjl7AYHf4urFhhjDQz0GUwHPmOQXmzigJF3jTJCKBHlM
P3oLw5ciq1Yt64JxtFq7YxPdXhnJ9qRVan+4wM74uIqWz2hsnp5wjfKcBa4sc1VDTYuUckIf6dq5
32Gl1+86Da7VkKs8Qns4WpPS4bkrIhAJ6axGyUUmYxzkc3VXCR74C0t5yUTBCYd3UrfcH0fN2L50
2sQWbOxxIGXQWPWspYm9BYw2lmNxG8jEqIH6UBwQFHyjzyJD4+LYHZUepbXbK9XKniwFpVs5gUbg
s0k0CBMYi0yEytkrSRZu52sFl/vLU2HAuA2/FWRE15Dp1c6l48tB5sSx96W/MzD/2MrdQN37AoTU
z74ETfOnZbG9Of6lIz4bqsv4KukcY4cu/P8jxDct6ptyy+aurjDzPzt7oBKA7T65USKB6snJtgzZ
I8JDrnd0yo2RjNqL+USeog6OQI6g62JRI++GBnUy1xmuVf+DpmijYqv1Slklm1O3PCU+fRUFh9Tg
HjaCn1s9O9L4rOL4zZ/KwWA4vhmizIiK5wFKb9MOTQgzEHk18Ap0FAKv0EUfxr9WMlgshFihTB8k
Co9CWyP6K4fRpLGhoE5S80xlTigHE68TquEHVhF5H7Lm6hjAspqHADr1+S/TZSp3Ovcg6DyyxBaS
ONi+K+1Cc5re0V+4hQF5tgiz8GeMLtmtWuMbYuP5kkOXzN/9R3yCgj64qlBIEeAZqLq+vADaUMGj
OZzY4PGBVhjnsCQMkTT0oIfzUqTEg9EhwW0cjpeGP0/7y/3fJQMsndfEOIJgECKWcY5n8lybPZG+
VuNgqoKFUaudAVYzIfj95dwC3ZxAKGdrQYcH1yQ+Sqvmfo7a0q7fbCzIdlKAJTEXgulvefprNE+W
VlrEzxp7pQ2TFi24HdqtTcnaK5DHBsDVzprT5synEIJJwp9jtUTIyBb0sbD/haLQU4JCYgYrFsKj
plyvR2gGxWQS0q6Nc1r1ic2EqAivGBSMd2V8l0EX7O2i9wV0W5AwowJkH33Q7eIqknXk23zPYZZ5
GkJQSObVYhDKRptkUOPGju953efNO/na1O84ox1N3etk3N6I93a8virpPtykYHpmHvi/PkGTtSxJ
Brtn5PyB7Q2pGWaN2cAgToMpaVEuq28QrIDdkOq1LqZOjJl+bkC8NDzHHQjJX8Asrysxt8GVx5Uu
CcI8HrQClTWzPsimQ28rW055GxoSCCxeTaSp3JOVZlTu/8pvo5IIXVPLUHpfzPY/t2vRLmtvD4vp
xVIE9YWboWlKdVMWfw7Ozt7pDidqR85+UyRo0I+ZM2yCDlQnnls+orfL9RnbJttBhlWXT8wHVD46
0K38fbHackgfardP0BZBBI2d0N7JF9muIp+7H0+IT4jabP+4cWAOgbGSkS0Vp8rlihSflW/OTPIc
3WyneUlKnyj8geMgwnUfQMjG6DYwdseG9uYyiEXA79dI5y/p597QYYLyS6E22hbffd8fS6HKFq+n
o2wCrGmZltXra7wQ8kI2iSjlvNGtKjmH6wbpfZ9T1AXfwyWYzAnVlSr5nQYjYjVugpQVfPbYt0Wn
MgApu9gNder9HGbB8/77nmCgmVhwh8k95u6VXX9bhrghSGlep8Aeu8/osWkNaYcZsSWd+bMapszR
5xfrfvY1tizs8VQeKEeJR/hwGka83LZUIX9PNs0Ilees9vs14SlYM61c0KBoWbcuBXXthluRqLfR
6c+2J7jLZtIm3RyJws9TQvP6+2Zk/E7N7HxzDah37JYXDwrK+8QgjOxeQz9jk1B/THnBBjtbwKT+
QKOMx/i3EZxmPjlVAOuyOGuDiA8/QKdmuQ4MBlNxgVoY+bD3qPsRlmU8B6jppZzzj6D5YoTNboUW
exyA1TkYRxwD6afwNxrO9zyYtKVEBxZ9EF6CbfT7MRHYmm16c12mj+5SOpLSSV4MMCjBM/6qvKGp
gwasXq5lP1uh0V4+28DCpEny6qxYbQN+ncTSQevcOpHSDAKDEFwtT9EVCK/3KIvLloBGMoVtd+ND
PDAmJTis58w26UwkHQfxAwYDZvV10Bz++NeBHkOccvemvZ8vPFi8mpP2gDSKlkP69cNsB2Z5g4Ui
4hCRVLzrfG7jF1TL+HyMkyYj7Fu0XXqYfujoMS9c7Z+92BU+4qLgtQkx57ygLO4GSjEQiyJ+wmmn
Iugot4mQtVwLRMehFOYTBy74BwPfvZ0bsP/7z2zbdCpjhgi+yzhPNcSQWLHUcGnzZNR7IwGtWjhm
DYrCymiHp+mBn4q6KvFMB7R+f+tHMyGsBkPMl3BcqOF9DZsE3x81rvASCMqN46Mc9ximIjHYuHQd
itJuKa5nuPm5HC5FmNCCSLOoXMLnTUVpWSJ5e8URqFanUAaMCiv3whASSy1f79qgFCzP7kI0bGSy
UZmXMiEicUBftUI+D7FXZvy9k8mwBlNbhKxuYAJ5RSI0n3AbX4oLlK0bsD1ZxZ2ZOeLsIGP/iQqk
6CqyM7O7gKOIFs+x23XavQYqwu1sqIiTNHp3w0B76XC9g03vaOiHu+Pv/G+WJA9I720lKipeouZ+
368zfgCCoylGFRhYmD03f2mIZab6FIuW6Q8qGh7tTkXmqnZPLda7KJZQQcUZaGSFXKwOxZq3OaZG
Q15G+S2F3iJ9UPIS8IscvipuAhf7AhQJMWEcK9KwRE2aD33f/fCxnGpvamWhhwxxjFU+pFU0GQeb
fvFpPlPzidLRyWfuKlsIp7Ou0DwCTa9qEQHKKIfLOVibmKWSIEOsGRfcEfoZ0S2UMh6GWAPbsTVc
sQNJAZ56C/0FX1HCjtBI+CWKMSi8disqFLx2Y2BZBTS6lPEai0yDjTOF4VRKdlVj5vUt6OfZwy9z
D8jOxoz4mHepAyCvfYitAoTzvyyCHfOEQ6rzdZPxS3rR0Vt096cPM7AozqXJXcvrCTjsAQZQGy0a
vJ75oVEjjz64JSU+/jo/Ditw32PdnJEo/+sfJVLbRl3ZD4Qq8qQmeL+LKmk0Kl7G8ufzW0Nc/Wee
H7cD00Lmqwts9KwCWsmgYKxm1RvU+JGKZxL9MEwbsVqhTq42iuMvgLtySBA4JfAaKAq62HruIFor
pkDyhJx4azDKRLGhHxlR7Gx58O9kFv35afcBFyZ/z4ThQ4iKV+jCS4osWpz/FZh7Xdkl0jokE5bj
vEYP1lktoU0O0yEDZ95prL7tA9X/Tc4dQVXMMF4rdMirJUmN/6uqTWv96zJMouUAtZXtUtSSpWiV
P+ScAtSet3NvghAHX2llV4R1L52FVmj80K1tYv+N9XIzMzkgYOJ1CZzRKrahwEwqb3Ij7R1VP3XD
PqcUC5B/p25kXiYJL0geFzlnDsey+m6cmBharcTSmd4E2K2c1pr1I+tolxws+pHb0DwRf8ppwQNL
MqHeO4d3foP7D7ZdrlqgxJ4xWDeG0rZnrZeEHMBw30ryP243f/MFzyHI/yXTxC+dc7uH9INotPIW
jXotxCzz7UwSbpxGd3KBirjwM7z7xJZnrErP0Kpq1k5QuI+4dcUt1eTghCNRHUzN4atG6XWzL0JZ
Sfonn+FMYZPMg2mgEdhPkh8BdL9W+uVkS9WudsE1ACuSc7ie75JThEu5wg+osConZPQmClLt8oLN
HZo0hg/vgX8P7dyuShrMZhS7GwrhAXU3nbJ5hoBP4xugzcTInhvfWpk6BDprZ8vu8gpysoiC4Ivo
MYYP29a8nkHRc80iQnpXxVAvv5iK3r9D0EqtZqEir18srFJnNptVbnJySHqaH/YV3St2+EfD4Yq5
SltWMH0o70O/r/kF8T0lCqeCzh9bCg2EibqNYrQhy+4UU0thvck7inYZEVZ64NUjNZEnZvQktI+1
b17NPcV5U7Te3UESlTiIXDR7aFrFltMYUcjlcB9rI9BFIxHe+jZ1cEJ2SRD5nzTzDJlC+tngw51I
2WeKkgT8kEq9kD/GhnlAO/pKStdyF6UN/+OUgtbijXqKKS/k14jc/pLuVzhiKFp2DRuTU7LB54hL
ZXxVhK2kQnuoP9sdC0w5tBgzSDeBWcibqNkCpK8IeFg5WHvd/DCJeNVTLZ/WBkaku9uDC/A3Ammi
K/1cItTswoUBLPGNAknItj866LRu2xkwTi83wGywXKVLuh01xl6K/AFEzFEQhhPSLbUJAAXpUA16
c/sZGs4XA7zApZbd+L0Yg/orVKi8QQddR34GmwztGSmQiYeewfBkjCxPnqRqqi2o0/pVMGVeckbO
zvJkWj4GrPirFOKmmX0NvT72AS6WlcttgNZaxla8wHTvyW5f6omPfsDnGkdPbniy9ShMFtNSJEcC
mIO91PtDGZgqIOxf5xs+D3Y3dpZL0tprbzD5rVEiVcU0hebOe4J0fnwq6XSriIPNBTNCRcCqyb5u
f2sscOX3mxW76zVN2xxuJALw0LW+QQk86wvuQY9G5cMDSM6eQavsB/u+y8YZYiazbSVJ/Fi2SvgK
psu5Ns7jSqXDDwQKRoYQGCnB44Hnoz1QbNB08P4iiHsCDzjxITUAuocpDwaiz0AM/Z0MaQy/VuBz
auIBoYtSBxbmcPPAZ8pHYi5IoB6tYs04s2OORbsMt4Y4DLwcAHkyqI+QNDnOhHGKY6hVNX8j4yqf
DaIhikOIuIcbU7pbbS7IBqLuPqrZUugK/xgZzHmdGI8d77bwIsFTnd+zbrU0uhWAsNZ2dC/KHbEZ
uRlNdq8zM2Q6wpXA5qgETeVEN9qqAItUUA1o+cU7mYmzcDAG/JFS8rDAzlpydLxQ21bpNIA11p2Z
MxEdPwndYTkimMmNjudxDk+M72p9PcUAJT+nCTKXWZBVLmStrp+J4u93MkQIWFCtNweo0HCJiWdE
e5Dvb4HlljY1X/vJ3CfWVyFF1LUHKXszJ/dnu9XZzCajNPUG6K9o4e2MOk2FAUKxUKRsu8/FzrKP
Jt730s1BJys+0Znrz/j/77jcfqNP2RePgNLrs21t+xs69a5Qpm/QozRNEaNn7Q/eIu7CTpNvnRSu
eCshi8nfCjP4ZovPdJhBDOEzQ/npko4Q4ulY84UXLd9vVsGrtJqJCswoi2ivJ2D3Y8agrL5iNeUu
5K7AJZRZGBg5rcCYf+ZZ8xg7KdaxTRrjkiQ6rZg4bcmklWI4IPn/Lz0J2SRc/+JPPhyOWiuOWReN
rCWTqaw85mpphfF/SldS6BjxXmM0oHizIYqHZQkjzzGDZHuePGJt8/NYO9Zivgq2DV7kyZzkeJYn
Bg1HB7bTe7yQhRq53AxxjsxmbaMcTFL8mJdE9cdvd9XEaYYDy88RH2yGNwhNNtfB3TwTzqYxVu0G
JkZZWod3/xjx8da9ct2whwM+c+K7fEnlBoAqxo62KQH+P4DBMJIG43qsndRri6kQOtM594Q/F992
XiKpzr1L2gOIuE3SoRl8w5jmN1ZRvO3+Y9c67UwAJ5O/ioWwVVM37RRY2J9qwAsM4g/nc2LTWruf
EfDSl33UAxsCL/hnALGAV6KIVl+u36+z8b8aJquBH05jcj5Xmg/0tGdky+H6BpHQjgxIM59jPC/u
nn7dFoSoRew1RpcHaw/Ob9NIfpPPbRbRk28/cD055q1ZYc6cIk+XprjBCoR2LKTGTTTxR4C903u0
cbkifAvANpCjnwfBlJJIKU2LZ0j5Pe13dxaDnxIEa98Bd8PFMvd49z2EUz0HcaoxrNvqParqI2fN
ZVXM/oRpqFcFGkwtS+BYurhP3nS5xWbxqZ7JcJ+M2xD6B2weJEIlDbKOffmOZwa4ixLJBlLl64Du
V+syfg4JVkNPLM2zjaFIh1vFReWkr9kURYEatN3IflKph7H/eEAf04hq4NW48ptgiSpCFoF+dKDe
fD49m8K0zp+yES6+TXqsCAYcIiHETNmHN4hE6SxHBKcKM4Km5O02jkT6rLmJaEVMP5iYTAopnmPC
j0D59D+l/IJunVTJ2U5jn9OIbw/OVXIIyyFJeNMYRfGtsAjMeKFypBZyE7PqlQxl0svG0U/Wu7XT
ppiEei790+tvsiHXPb4ZZHPtm687py08EWzS3gaLvlRVfhZzubMkm+qdhA1/3TuUrUfhvVlJ+9F8
ZYBM7nUBs0yQsH/Uh3rgLPWYtirdWWU5GkPYCRLLKacUz1kLJmlGl5sJQnIY5jeSm1NDrQkT2Kb6
fpnidzTxhrEo2ckPMMpNkn8HG/Ox+uJCaL+k3j5KxrnkVOtKNAb+zj44/410MwlaQCweNG9Y2CT0
xAdsNFxBVYYMU2F63jMjFXO0BWu5G4CUD2K3IK/NZ93flLh4FiTMEVSShdvI2nDes3M+R1aLS0p2
snCfmorLFKIhO7UvDREdBqNOR1K3nDeiT7eGETXPTytU6RdhnMmG8EMQG8TLir+JN9EPr55fYRxf
QyFnsy4ekolFd6K9EQS6iYcU/e/obeAWBPHnaLpnncvjNnq1q1dYNbqK8QTTB+MaNVdOkc6/bniC
TvQsnL3rZ65TyGyB9nChPDNxMejy9fcZTH4bFAlDVNcJeGNa9a4enTRV6ADc207R32dqp1bs16NA
tKRTzVn+NdxJ3JzTcxsKFKaBDM4gCuW6RFXdeAFiiWOuAdD6zS23mP465c9tmcK/uY0tAYyFfvfV
T8GJkXsgcsoAMtbUPrmF9yaOJMU33+wZmJBMZ1A7dNhiQe+Nj/cJLpJJAh0d63AP2p/S4F1J4a1d
9s0PP/gnCO+HINS272kCM/6HyLTCLyL7fqkUHS4y3jq9sXiDE2w/ZMS1XHUzNlR95qiTNyOCKO+3
vG5UlwkBN0/LGmNXaSUSsVbtNE2kNcDl94B9LLRaKuQTZow9ZIhnXo8rvI9u/arVe5Lgnx7/Bnmf
LJbO00WHEMtzFLYOD+2pleLGfIFzwpsHQQD/EArL3rgpk9jEHSOMKWJDwad3s7YuFVeFOnfgxihw
cqiMg83LkpotGmzVrFbFv+NGFg8XCC9g9lrU8qckSwG1pAqMcTU5yH42cfKvt5Pvxu3aS50AdM4a
Qqwz+LmQvU/o1LNslEiBGeY787FET5fqu6ZGAtT1R36HmpyvKvSPXZt5uaviVhGYurbmyTI4Qx0j
bj0GTkKOXzuhks4L+or7OOupuapZbitm0mhdAJbbunhXMJm2iyZrUSUS7RuZA8bz5sFNXVsA91Ka
I3FUgXYKcMCwZ2es8O74diDr0cRy6ZfHuf8KAHzWuwk7GOoo4vDvLwEBuVlFkspWTEKDMGC4hJcj
l6d80HSNYYWqyWdGBkFEmP+ywYmuSwWSuWpG78rc21d6+Rz1n2zxjZ1PjtkxEQa0XYn60LiqZDs0
SqBg7gs7JO6oMJ7ECsLOoxetpTf6xt8Q5M4wyuUM5Pmh0HTke7LNPCTI0vXe/qSLowv09aEDADVr
LqyoSK8j75eQlOS+aAtZXFMFHz4wlbwGCH0cYzMU7f2q1X+WO3c41n+Ltg+1bKXOk5dTVgzks+ah
YqSoV/UmbM8ReAuVBt45GSNkl/bCX7AHyvvYRvNgCOj0uoDm7h3oHEHnacH8phjKPHDNkyYXTvfe
piJg32g7MmTm3Z0050dpCZNCxrFyc6xSfswRuH5yR6R1r2LK8abm0D3iF3OWaumOTbkY+VGAKppj
kSOSKF3zteuMPbMA76GXIYOFgubBVICc0Fd57Zo7DKmpqld2vz9Ejw4H/bSv7QpWgP0Vo51AiPsS
MxSJdEWJGaz8ROlYPtnV9uedSU5i4nzeot/aGk+2L8IqJLTZaRMyWPszfQ+j/4dfQ4F1ACY8eyVV
SKtP0XwsTIidu3hpV1s5chVuKzTH+iayEBfElF37zytOcO11s3dMhJbA617IxksIbvm9oqGCyDuQ
rH2yzIcGxTp1+gs/bhg0u0UCmsypjzLDUojZrG92qEkJjBLVeq8k+ZZQ2R8/gpGwiB5stl897C0K
37JZBA+M8ayznGlc4+sCXWY2bDtt/9DEivGNPDjO05a42af/rHX6ilDEntXgM2oekDAoOtDiLvxY
kAbB6cQcekZdejQ/qJe4dYga47bVsOj+fGJ42YNZzsxzBzDfXIKxrtb34AIK2Z6nsD0j73m3VMV9
ymexW8If7pBu/cMM0QTdq3sp35GGY6s99p4uMUCCiEasq1VNqejbpgKidTpp4r9C8HesXDBYOYdx
fVarArauI3fWN2uNx6fLNeIxgPgW6Uh16mTm9UrJk55HBE3SRFf5jbmZNHelV5QTCbL0PvL18RjI
kl1jyIQuh5khhO9niPCtUBD1AxwknZcnJumX00knw/0MI9VOVA/TEkuzowSDhsfwlDw4aK/jyRDG
um1nv0pr3vMQDRfLF4cLX/bs0nzAkXWmzXe+LtQy8Gl+vTafDLTaJJiJIuEG5HaROJT2JwgDyo88
+j6V28WeXN3uyjGVY0Tf96FWACDB38eI+oed3aUSow4NMQcXHF2pPqpO4m1rmINOhnjspnGPzmSC
WOsnP+pa4KMEfrw9MLVt4/tWp92R9/9C9xexYU/v2Up8fMln/DZKiq7MXe5TWQlWx5KSzq/AO2yr
dUbsw7e1sISBzIsF6/HBIbmuLhW7ERV79EnYJOR80BXbqfyM66vJkQ3ZFrqSvpc1DSWHM19gxI2u
Tf+/+w+NmbD6pSytGyDKkDvm+ihgO8hpSwIY2/a64gaF/xTrtd962BzEcPjR3GZhzxa4kKdbL1Y/
5lrJl2p6glpdcw5vqf7sRTn5fF/SWhxcAL8OyFmgC2BGqxjTPTPhuZ3JyIoR7A/uJTg1OlbEiHCS
1RCHAM0snVTls2jQHs3UTfZLrmXL1eU5iaBkVZciDkB0mEDLr1qQzwW58Ilh9W4nj+OjHi4d8dgq
fnqkO4YmT/hQcFEkNdAJ9QOgAPP1LCTCPEsz04KAF68r5nPLWueNAMwXyvAorJFYiS4tLFTbYDCE
vtJ0R2HC8joo+WVzcD17hnmBrwHSnMYXtVVbY2iVSlvn1VsfCo3MxWHaL2UBbWdAaRn3x70FdSvR
EokfBZiY1/BjLjq8vxudOaF0mIoYwtzasqThSdrJeMTOBUdEe609GPNU60v4V4Q7oAw2dK2capvf
i34yzIrLzKQfay7lDxL8tT2v88bUQ6xNEDfvSRQV0/tODqUp53KFSv3pjHKcbTxNwWsem1SPqWRW
RSUaulZQSRnq3RVdXFwMN6GY/ArDmv8HQaY+RUOLKso1rmIOJ3C83MNT37RLI8rm5X5YxGsZkfoX
wAq0S76eMGKYtSdDX/3+i6IGh6VgUHOt1swAFGzcrrHKXwMy9i8Y6AF+tBQCEe/r8OZLOwvu2x92
wKpmhMGcuADsJqIFc3J4/H/rt9jJ8PpHyFKBtjb5Bqu6bMgEKy3P0WNhTak2sMF9brDukRPFcW25
0lFRlvimfcu6uL4fY/jW9BJD5Z7WY9XVhDMFs5l2yY2SD3O5m4NNCXkiWOsK7D1Ifp8M6H+NJwxD
WR22CBSNfZnr2FEObDXHp6cyGXJ/EjKnY7nrsz9xE3WnHwrME03ATxNX1MSQy7lP0XK0eiMzBxvv
Dnbbm+SIfQbFH1QvpdcdyeywUw0MLKJnBMMxX2ItrhEnF5Fx8UZVqmafx0oUXHQNeEoq9PNxw2q5
Crl/esaGiwDp5LUNhauxceDrnlosEGCEvzz7uC4SnL8N6+dxfSuaYBt9GZq/zqlbBTqnGhFRvEAD
lv3IlFzA2njTu20hsOBhjWop87aH4sjVFfYnoXD7uhEgyECpnNF0tfs0PaeL/x2q4RazyWAUesUn
lPUL6Ypcs36GyH46qMMPgdB/eg1+DZdyuLTY/fynzvgC0n2lXcD5ACcKmhhm9YIHl5Ib6w06RSkK
9UIffVY/E2KnLwklyxsfaKjsJpI2I1gdKAoc9MqAm+qqy7VBlyva/18mKIPEpIGWW+6IAxGGwros
w2FPQb6ZAWvFYsIQlRMxdejszaJGGt7shQQN8jEdnmeicIoLpryMVz6gOD/taWCdgacTuZrbxhgc
7v9Vcacv3ma9+ket7+ls9cRiuAQIAFz/Zo6E0gAUHcjZfUpMgo6pa5r8dfvU2Diqcn9jQLSR0fsu
LiYn97k7kKUMq18bPro0dF2hJgwPm24DXLVugUhwZExpvgGRhqS6U1aAbse/zmbUqp0cDlyN8qCG
JRxVP/ZAYwQaZnQjm/QCx14Vcn5PR1YytXwu752dPWBfSd+q2w1URCUdl9qcw//xHjqJ5fS+u63h
gq/ykB8kZ7AWWpyzlL6EMz/DVJjBXIODfYkjYOfefZtN6mFdI1JcaYTV//Uueqme2FmNXK8HBlUG
7GWpE+7z8rD2iYk5PFWQzWn2ThiSnpcPHnoSNfQzr0Ijhv7U3ay5nqqMrpDRG9hwBgHn1z46GVRO
nFvVMwStpitc6vYhVDZZ0Ss79z4+iRGsXoq6lUfasExxccsxwq5p3lNM7zZsg6hlCpUjaONCpvt1
OvLzY+G3dD4P7ot3WEKiLBd8JZ2O5VX+lS/bPAEiG+r0N5Qa5iYF0LfcPN8ANEn2NgYnPDJofmjS
rKtHe5TsyGhdFStK1IFoyQstY+iWIiR0EhT/3PldCdJeXHg/lMuoXNMpMvlETJbyNOZOORf/0j9J
O0qQy1f7JT8uCd+QCMXp3bwgUjuld9kBpXR+bD9jDy3NgIJpviaFpMaojpowGe16kvW9QxN4Dht/
o1GJpUy8XsVaqpxBe3FOZF/Q8nOuhQi5POPnvS/Ks6g+cVJY/9R9pL0+OpfTQesqlIrMxadynaPb
VPj17SgJ9GaZd0auE6yx31/4CqiiZLXH8p518WC+XLQ6z+BduIQGNPMh1yORzYiMlZMKUbp4nVSt
KWYxcL41V+PeHSRfOTLJhp1laiYRpuHol93VrQKCvka5CQhHLdc+5n2f0RZU7XWG2Lc5wAqv3TtW
GUSPQHTT0AJgQ/KjiZsvrXeTicwynrPGISP4kFTpMlgGIpQ7G8WD8cbBC615xZqdSS4a/AqOKEw1
pd88rehYo9ODRRRR9Kh8BrMFNyz5hq8weR2HLnXAA1IsgXi9z71FbWT56DG6VCxdqaBphhJ7MMga
++khcX06LYUrYGTAVRYbCKV8ZzmmEyPQ83PNVkHkdhXlO0oiiwxRlL6wjvudYk4qOjm2cfktWE9Q
X+aWs8CbQslHsFyZt+2bLTyCjaCMA2ZD/ub+qxF10rzVA/t1D8WauBxLaXMoSFClDEUtWL9lHhtT
H4tvDwPRcKsyWNQ4JAPi9lg+Y4zfwabsFL95Uqp/lQWIz7BNSFO541HCuLpKsXpdQksWp5DsIB1S
GD8qVCj+8YSlNoIuwDQYksiKTP+nL8LujHdaoqj9SvCllJcw05P9Sc914FmqIC/PytQHi4/ErY1e
cN9+kAyky3ch/p0/00b65R9mOAuw3Sj1zQRr5ERfmSkvkWY/H3mAb++nSUXZIaBB/DnBI/CSfDNa
PTT5624lF9ZLYzpqA9lFtlvflf9xI4aUOo2jQdR8z2twigo7bef/K0Zn857DL46v6PDVMti6te01
9t3muSVerBm29AnAMh5E1ZybH9AT66je4v1tjebY1v/vOhBpoqwW8w65tFDQrnDN2rU6l0MosrC/
0GjvUYwuD8PH8bxgqgiinUNz51ybG52GiNFhDfsxSIaegcMqk3mrfetgS1cWEwfMVydwnx1eaST2
AkOO+jE0rPu1eSe2/SgXkeB9RiPh7/qvbujQI9kcL4/+sy55WtAMNCf1e8RQgfMpdEecMeQGG4wZ
YF2r1S2QwvgIXQSAOfG3Xq1xK2FKhRH3EL6kfHBjpq/TDYw1g0ZD06F23tKnjvXZDDKJYKYA27nM
fJ+aLZbJv9qXkkm6oe+2bhXNLjoiwgyaaukimFEimUD8mfLrSeMILgAccbpSAc/yD4r1STQ2WVRT
Pk6UqdlA8A6rxds3vrdSx++shCH1GhN9zXaJ8MZaLUUa1LOuHHcr10ym7ssVgeVgscMspmSJWH/v
YBDuwfpC8nvK0xaFOzffXwluD5vw/plHeP6CaaqmvKFZRY30166SCtwV6OC/IvwUlJXBWiF19DMH
CwocBgjLzg4uxv+igJR3DWnLGqCX1tR1XcDHPiUAtLB72yOScdZ+NaIMOtCh8rqdy1C9i2MZ1Ria
Mhvpn79IVPtG+or2PzvaViJRZik/bBhqJFawieL+pm19YBdnPTmzYR5DFWRC7WDdlkAw7CfYYVKU
dSE7egpOKcGRDiclZYk4NGsPW1355Fcz3v8GiXnTD9dG6v+1Q2ME7/W7aBsfp28DPcoo5Snm53oH
4k6LuKHILK26WEmFq4zYmEEkM+YKinPDnFl01aHjHfhDe58UoHTWhYnRIt6qrukGJfpfWPV0RrQj
jm+PVT/UAaM4BzvxZCjMcEOl/pQHfOQqtmtHTes7mGGgdaBeHg3vgPIKjghfbPOYFrAdWEFwix36
RjNQJEdoAuyviFzhRzV85GPilsvzcGdVTtXSPg1jUJvzX1INPZ+bQo6c2cRjFe/qXEQwGXciuWuO
fqR9asTs9AJImyTNetekdAaSRkiuxfXErDHfuudrMRqNGGkMaYjpqC1NQLlWo9waGaFhEx4LLPfX
XYhyKp80JadPZ9+v8q60SNBxgTgdZfC/TtmftxYWowOeNwqU/zDtTiJxbX71I13kGVhI+a7O2+1M
yDshnsQkjJde9qCOYywSyiIfa4mR5Q5a5OIg/iV0bSDNYpDWtudYxPPVJv9VHSsZoTaefaiK2a8e
oKm4tKgRXnIqJEE7HtfedpUKZ+YVdn+C5NWIIh5Csz97Y0u28QYuv99wwD4nEL4bSbdqmvOSiDuC
1LJ5WPHtL6b2FlQ+O09Y3jU40imaEOZJGLJOUG5cBxSwKd4SvLoQC1dfYCvFtPL5/wfychRaKIwr
h+nsIwuDSQ4bEpQp6uG1nqc6OzfHP5a4IXKEklseIwZCfTaiIGuLadoStNNQ4nRVy0nntgIrGKu1
6g1fqpQdH6jJk2SLTNp2RMpQbWLk1nwz43a09I4VhfceD5QzFvFGcniwSNWD/59IPqLQa2JH11Gm
aWsNfiXBIK5V7pSwL/K+Q9hY5NpGYXrmlEusb9Ehi92X1YhsGLX8ba6Qi1b1A6hz2PMwbQqV2z0L
tkaM93zH5LO7yYwxMSaXvtSCHLe5qzLOTj3u6slUzj1CndzbMhHnuqydeG80osHTeRBftD1tuP0/
3UuCPr23HiqrS7CD5C9wtwxgpoytYFAN1YqOTnVUKC/2/BzwUP8X3fNADmxMVe5CbJurt9Wy34ka
T1O6XnXqR5q4PfXEYzChFbPvqZKNUYfbm4miQXtCxV8yCeyj3F7YSGlDNRgo/KCs1RwEV7MANyC4
OAObLsyuRFPHRhD0/GxfBFAIkeoStl64VzmVPw8/k3TSXHX7tSeB4zFJ3wVUGPPDoO/y7b7p3fux
uU4yBh8K4vjyRCBlJOSA0k/mHv1vxbrqmT8bFuga8KOG60xdvUa6D5z8VtJ+Yo2/a4+15aL/GrI7
G9KTeBI3cPqVsXav6bZ2cp3OTrJW/tcO63e5N55pt200zbP6k4t+1L9tn7U9BGjWMkgE5GpXX6j1
RB+1SwF0D3kmseZts8fFrOyZpnA0ej2SlzeA48RWX9rQBkXPleiG0IAh726EUsNPmMYcGmRFn4X7
E+c4ZwGlIOtFiqGE2s+jUJ/GCNfLkSUSS1w9mHiQLWKGvB/5sWD4yS2XNBB5M56+T9opRgVTpVla
jlcXk/U8FT27G2XAlGgfcUoXzhjfNzTa5z/kzHR5fBd91xa9AIm3ItRLi3EBwxcZMK9Ha/69sSk+
qwnvBZ4zMAZS/NpUHe17KBJBdFXJirKMpPfnb6tM9kZf+slFP4O+tr9c3+wz5+4D3FIhRClUCeiS
eXCgreB67FJM+spksxvFu8fvSIuZHeNwBYVurfnvm+L93SwpPtBe7T7fcU/XUu0gP5jHKEUIS+nN
FcOZU026GIsafU0WANuD/lQRRAqqTvg6jm7UiCAi0blPkINEZdDmtIx1NCncq81GZYnLyXj0nsiq
UC53R5yE82PY2i0lZIlH01RhhDi7QnDzYzZ9QCqg4FK4OySalfgTV7G7VI9hNhGikdNKfxtYdrgz
XDVxleN5jyUiyCqPiaXHAWnY10GPupwa6vJWZaSFcY2FVCCsZwCX48nrH3KH9UuJ8K/r+wb/tnSE
uljrSTpZS89UbQxP0EUCC/gSFXSI7XO9BjRrUpzW2S33l8J5+OjbA8Jt2tiUq4BmKKNhTmrVMDFH
0IhGNVdGMsARaQZJqnt6uq9mu1XVF5lvQ8cqIhfXeAipmnOROD75M3wJqNIJQXFglVQVTphasCZ4
9Wtf+AoouST3QfwHQhVHSHPOKvVXiCwoSiRd6gpeR9bDIZ1mxlm2vGRyssNAU4e+A2+YI+/V+pC8
7dgMcadWFi13QOIiGXm0Lan7RbhseMlUDtEPkpIZA/khcI1NxvlQfRlGJ2bFAb8qZlC7HNir4gep
pPUHsRHgWz/WlyWeB9lNrwQG84sCO1bFpiIxAMrya1jdrzMFWC30zo3pNrUaDfb3k5v066DNtmt2
1u3Sb5zROiFzfD4FWOf6ueadiZ2BoukhoeUwMtfGbqSXO6LtLAdxdhN+bJIMJXGADWFm7BiQmtIL
2p7FQV2LNhnq/DWoLqJXKm9iMe93VJ3rUf0fx1gVrhIhwqn3WAptpf8zouU20U36/JGEz6qYTFYo
Sqyj8YNUsTLRFB5bHcjBPH3qf+Fg0vLr676nAv+Ag9dP5XQeZ6Tlly8AWwuZ5MfZcLtZOlnE3Dwb
yuF1Y0OR+SqV925jsl2HF36xWpH/buEwxszGK76zBXPQrwhcEsgg8A7xw7hLJzHUNwsanEYyVtKF
IymGUWYItbvvH1sEhNnVNaWFa1kpurixYpBFx9z6l88AZ15r5uaKFfZeaCJGxD71sZ7/Qtypl9ui
Siu1l5K26E90GXFMQYAc/oH+D5ObEaQHwA8ucKT70D020hAu77sjJkKUSc2qtpo76h3tXrqDgMId
OshigGBaRg+RXfJvVPXvQnBpuT3YjBpseLSB4hxji573AeAQ//8OKsMFTOnf/AQ0zI/PFbaTczu0
Urp01shvlTIfciXGKNDnWbWsSO1feBrUgo5k1GiEmDcY1mWlE/0Ef7Il/2DE2Iz0ZNVEuEoDjgBT
7v8tN1I/0twlaluQ87hwrBS/sh4qm6NkLqoC9a//XXxLVOT9u33s0fxm6ukagKxba8b3lLelackY
ygD1FrgKVNLfkrHKzqdYOlVhd1YxgWqSYAGKjsCndX+pB949nmWXCO8fbGwJC4ozBiLURHSWQM8m
CPNJqI8yxLDX6/esRVRKOk5crd/5H7DZq9KQXkZ1o96mqCWt3Q3QvrrNLUMcJ3/N9OIcSQv4hxVx
WSWezELkiZj7pZDNXGlbvkZHbZ4SWVKQYSwO7kPRT01sm6eNQo9iZpVD91IJ9c4IKyi+2ry27O68
HpU/d9oRJFWkxHJzOEFIFxKugLTSrXFm8fIoShFeCKjNWNyukXk2WRWBN4Oj/r7+toAOya3rXkbs
vNfC8vDP/cAY/0rU1wrb4Kz42a9H72t7bQt4qYDnuNL1JuLwHLLbfuMBMbE0HaqArfuwmaSwFoCW
y1Rx+tYh6O4Fe01gm4lYFUF0JhPpSmv4lu+dA80nMCXipIGgm+Zp9fbgIaUOJbO2o4b+ssGDb8HZ
0AdT3i5WawJgh1FsQ4bkdRCnat44FLt71c/O2dWPS3nZVL8xm/XZSgZ40lzevmmw7xMSEyuRC3gN
Z3mQi9rZzU4e9PkK6GIsIxscEXpnCl6CXIlZtA0t84No19Wshjoexso3zisd18P1ik/SjNE6kvqk
Xqh5gl/9j+qmWQOEY3bQ4XdXlfAAtd+G69CoDg3cEd9QovlGncWQIrDLyYzyY/Kzi/YHBV2Oq6Qs
dkLeHmYOBXA4HvdZ1X6SPmdnrjKLgMaVKRzGfBtzPG5R+Af32acscKB4R0IuixUS7wA0EeNjnfzR
RjpqVYi3+z+ci8w8DzApLWF/OCuoySVuS8nS2nG19wXSMzk7r9NRy3DqgJPu8CZnpnzSl8bu1sdn
aVMUT6B8DCvHA5L9kOtZSbccj4OknwEP0giovekCXvZxjPgXnVCpW9Z5tvO1RVTgxkeBhf5db/Zk
01SlLVzEPNuhGTyKfAgboOFEkNkDxOzk8KykUJUeWmhfG+l6sR17uFlky4wLaiCmit79qtnMQsba
x9/IoFDNWvNC3xDdnPbhsxn59AX/vYmF52d1VKm9F36Biprjeg8iAeMExkbfzIoSrldHqFx2Y54N
c6Z+OScxOTFY2Hfg0ubZW93PM2jq65Anpi3u2zk++PM1WgFgCOOhjjEQfE8uLHpeQJfF4lfAkx+Q
FKUF6EGCNduuvabsAZE+Cbw2kOz48lwc+YpuRdNlsjMCjzLA5v0ysxnnDcSV/XAuceLJMAB8LMwZ
2VxtF9L5ALnNnawyFcLPZRF+k6ZjSFbUWVZykGZJ7ge5SITfnMXwmzlThHPcFLAEXl74/zDpcEZz
t5GnBXVjiOWE+vh2wB/QYFYqxRORwpnzN/cb/imQYD7cP+j5D64hdMihQJvsek/S+ACrVnYZ1HrW
TWGHgZDJ56AHdJqRcZHLuzuyha+6AUpRx3f4aTSczgPJu/9cq/49TWGL4xbFlZZLGJmseVE0b0H9
UPHP5DysGfQA4dNIQDMBEMmFJgljpMMAkTgbBee353PLq1OWUgDdTHry62DPPh9yc3JMngm3N/pp
tei+tB+fyCBCDcLUkYwTZ89YHDOKs1znzGz+N7HOm+r1KTe+jn56agWjtGtKY0wiOtTbbqIxgsMi
C5tjJlQrfPfk61KcoZNoZxN1h+gizW+gcrhXJzg9ecRGrN/OKXLhNd8AerP8x2q4++GZHKv1sRXr
3Po2uUIVfhaVMtoYBOwLch2oAIpTmt/3wIb2z/k5gRuV21iOGaTF9hq4/r84SPpL9EUCev+QWn+i
5Iv0UxGwv+GapCPhJ17vIvaV47GHA/UEHpDzLv4sF+OliR6ZJOfOrXrNFWh6+Q/6QlDYToFGD/ps
qS8bkztQ+4uZf3ytcV6oTPg1seNMUxQAzyoCgvcEurNo9KnJU6KFvOKqUeAoT3/tOC5s3BepEJJ3
8iNJgwNXl/h40iwt/rAB1sV+Vvb4w+Q9kh6Ik86/Bng02xY9GJDSyd828OBv6SYnpi9SJ0IfwW5q
EaIykcOz+tcwtbaJGxkrLqN37neCpGqiQ6tZe1eT1SmUCmbpgADJdd7xdmRCNmggJ5tF+RIHPdco
9hodLNqrE60waDuZZZ82pl3OKKwItGwtmHH1rhI/fDVShH6CKYz4Hvy8Wu7JtHC20d0g20ANCEyI
ek1JGPM7+pERrq/GuA6IfHUKhUjWUJaoPVIlcDr8BQ607cSxePjgXO1aHHeGewRbdRdQ8Z03izCv
bKfRppg6+vLxgeygfDLsmMhNGLkYAG5Hn4SKwjKglnnmz0tr489XYOO9yW9NJReuXGg0SdOVaXWm
WPXQ9Se2sTTNo1OVILZzG8g0ZKzmdjqM1PIwRrXXMn1n2EOa31dqYKS6lcssBu60C72yOlNHFZmT
KfpGaoxdayFRNSLuqA+VZhrUdzYRBeupGgoSczmz2WOqY5zsqa8sp3d0YGp8zfHIHAONejBzM4Db
VSRO2uhnhSula5kKO3uIMR3BOwuW9TIDs23iPb9olriKi2PT549A5yuBV9G5FD10883zJDUVTv0v
GRwL8nm27g9mwtY5GgOqmsml5YH+lLoPehHmDlHsSC7hkbPp+Xs+rhRyTMV7fJZ0SGwBx+o7Crxc
FHc12DGq43r8oz2/3wHO9YCq9n2De/xV4j3rK2aEKP/8szyBxeCHwh/RE0PI1tybpKyFFY66eaEN
eTmsX/jFGX5rhUtGRZk8jwPhLALQ/QoaHt0V4dhsoBrhUk9c/CAC5ppPeTuWcLzfJH/bHBrzbXO6
BCXwEMbg+SQ8KFUBwkqP2AAsug9BFTY/aLrPGfWhWri+ySGhJp/m0cD5PztpUn28ZWrMazhFdKSC
ak0WVnQfGgS7nWQZDBsCUXNz9EalqEbIXS21ITp3VCUvw1vrsjXzVWRZl8AVPgA4xRQOVPOvAQpH
6hCNwVihQy6Mpi7dBzcivZdHc+rQGDvdwO04GG7OlKWQnjbR1aflxe9HdRkcNQkud/yp5Vo6me6s
CbTHt7FZrfrjDah8Zyz66C2Urq4WApK2+t+vBOrN6lRzWbFfZ0dK2pGL+Tqa6Hh1BqZCJWNcWjXE
0GTVE9yg64v3HdTjgp1Hivlw7Ti43jLK4IAu/8fJln5Mo8Zq1ejVReUhv9CvEkczJpBsr4zcTolp
vdwDyMluX7BrbVxIzwk8ybJCrWdjGgTfDIgfrub3RavZ5KNdZvwzcRmHdB5vpuEg+QSqcOWz2sub
zjBJfB8x8G4HngjaUBiJsmHmb28DznTXT3oUEI1mt63dVc1teYcNUUXwTMhl3VpSRihNGBMWmawf
SB5B3rqdPkWK1lKEgGvtSV4kTtxXi4/OKZj2vP9tPKnis9RJxffP2H+OOT0U1KPLMcWIur5KgqeE
okH4O7Jit0IlWdZMlYyF2pSsIoO+PgEC2cC9P42CvYQnOwDblrQWZykzafgsNNcb4v8LJpiIAK17
ljF5AEdolR7i/KZuXSYs5BjRb4IZJg65L2SHzuHE0jXUsNcJEgrDrtoKHbhDNTs2dWUJVYGEC4eW
pgL10dID0h00vkK6PtfONOJWfUUfKebUAytf3uWM4VDttWdjw9+wFr6coSzEmE0Ql5cC1wwlEKge
Nz15rXx4ALsigEYKYJfEnp+3RXtCfDFmz2j2+Mz7CETNJXjV0rqwcu5LrLqcOg7ye60vf3U2GZys
f+eH6UC1/4iV/lg8aPd46u4w13ucb4rYLNdQUQjb1iS6c3mvMpUgw3vuDa3+998+FmbtoBFDJl/s
ai0vrNulMS5JuC/83Fnv/g/zcehqf1hM1C9N/GC6WhyEVvVRtBD+G4D3iHbcSKMzgy4fT7Vu9SjL
5viBvH9TYVPD19JXT/3eCzqWO9o4nbkd3FhkEe+kQBUcrgJm/vuqMeathSV8VaQ1H4l1J4KQO+Ww
HBiD0R5Pt+G0zRLhRH8BMEtzuNEqT+7EKPBpQglTwPISe4B44wSCPvG+cDy9cfZf6iqffg3FFhKA
mKQCnPDchhZvtOGOcqIYxchU5czg4jY5DxBbYn8158NF6MqUmJpyBR2PrVnNRiAaPl1rSzySmYW+
3gyKEb8z6PwdX/HEiuDoTpa3p/KHfHxRJ8yDH2G99PToHzUm6eNLYsr1bOPcZ9+CR4ksJyr2s+Uz
A21Wb90zEg7gTSXoh3A9g5FBIt+tpl2tAEGd0OjFz0CNijcnLlPXDphsuoBjsU0xQDhpOPaEc62I
aT6S+dcfFEViQ0zZQ0uLoVoVpjDBo/SQcxVSYlUCBiiec6hc8UaaWIR4u8cReQ9EKOk7rfAbNAWb
3Su4UTtR6HzK7qQvwrfYOpfZfstJUFxKwzFlPpR1NzOTtdl4p2eVbv7okiqD5I2svaoA4i7VgSMb
zW872zpZJl4VEBA0G3ZlDL2vqKRm0sESzB1pCePxGnyQMLmCw0FaW5cjqyiNAN0fkLMTf39HGvYm
vwgBru7fx/2EPx4W1YKXYVFztkFQLlOKSRS3PxFO+NLhsoJmQIkbEHVqJzZ3H3ydgDQHrqfDBDif
ufnJPcteDlV8FqK/ZoKC77soHqepuLFlqERFxHx6cftxtKcie5+EmqCfhBq+8x+fj1TO9tjZulO6
GgkfiQ1Ze4p7/1/DB4grGx5X0BamwGp0PqizXXnhViZA7GBAhdAWy1K5qhIYzQgq4ZnPQOSPEEDH
3XIX5udcmPG4D4t74nMRltixD+Wb4IWsjIF3ltX6GPlGd1kZw+JnQ2SQWbA7xjveYmDK1uExBu8t
Gpzx89ZBWRiPK1FYmSwQhOsgjWpq8YrCmCJAIRKsfUBHwYPasZNH0przSR3aDsLy7Lm+LZxcTMQT
tJq5c8/Xk4sBAqsvsaCus4oaYEjN4rSyWM44g9xlfSHhXO75w3bZbh14g5lREF488gq7niPTS1NF
iNUG6zlnM7mFp+PcGzYYoMZyfgj2IouqYTmzwGprXiUBlW7dUaCIR3eDSeJ7YsTxzF6ZBUSyr+Vi
E/0kwKrhk7qP12t0WTUt796NZ3cYwuu6mK8nPo8jLivI4kZhsTEfGYvDPZxEmcKAt7IIM8eViB26
X5m6+z07Enq58RsuUacs9l/UIp5h04Q8CD8EMwywmd1JXeCiVij9AEL5Shml5f9xuhus101JuCul
1EZolaZVcMTo1Jb0ms7G879vlIKg8dHpG5J33zJqlm3LBBA4kNcBUr+cBkUjJ4IPpQ8Qa6EwC1BW
W46rCjj41uSeUpzY+5tQlAAfrXhoxG6DmK1VpoaNb8QnGy9fKAXJEAifQaAwUvtMgARpzWr3p0b2
mcXgC2Zy5T7MEcnbY5hY0xd7INo5o5/iO2FeYJaURVBGPmHHLs005gxXB189a5DsUp66GDLRJroR
h0+bzqhRb7yWp0kuU8IRttH9d9E2A3oiT7pdM1TSaRJ8HLDF06dFFuMTS2c//VSY9OGet1v++4rq
Wzr0lEBmmcdY9wmPNcJFVD8vqivaVkHvr2ECDOUd4PfgTKzo+3/j9lNZ3Z1K5LswgIn9Waqsz05x
KFD9/RUTVLSyQxnCQCDqHy8qll9V/zO4oR54cpsHvPtZ6hvRQmTAbZN8/enzNFL7CRGjFySCsFVp
sLY/eLJBhHGKz5kBp3xlaiqt5o2x2lQgsCxXN1nWsDe8XbGUz6DHgsnA5mTH/2Gwm/7WMNsuTG9W
xVEu9O8D7INqfDv9xxTqWSBK/Y3fUXxHstwdX4fAxGqqvRkQs31vfmLOhzjAZSkTwdDYEJLMzexg
wOWkU5ccfSBgCGc2Z2p7YzZdopgEmj/E2tUYdLsyNsnhTTEr1Zks8aXowPx3Qen3T/PMKq7wfq9L
kaDSB5GGdniqzjatJLXw1Nfjx6jTn6P0FuJ2IryGYgrFz6nDxPRAp//NXrbModo64ZxS6Dcmd6gE
c4w09pnXLxt4j6dJqmo/v/wwMQl3IWOdpSO3wSzviMMQpwBEbfUpNvtM54DyKv4Vf6fRvxKItCC1
cQghL1eb16MeZvxtyxDrC9OpnAEuA7SJ4Xfv4NE973+KuqgmQnKBa8KUGalqcmKgaZQjBwVrKz7u
CkaNhJZGIlq2U89zVlZ5Cy3ZBlfOR1nCOtv/aImkL7LuZMhNk2RYcQuuBnCNpryeb9SniLtYn7kJ
Jy6fTQpw5H8n1tX2gITALRkBXwTqRih5QpCTXKY9zmQzmZc4wUtt0VerRXoZ4O5zmSiyLsTnQB+Q
oV8hJWDjzf5W1O53Q+gZIJCqcexivxmnulsTM8CPP+UJwuoFXAq7XtcwwdOSbq9AXAdA0jkmIx/c
noXp2X0sUTNblQYb7fVdaGv47Me8hftp4pNjgn+QnAZmQTeez1W5V3jyS8Zmk6VTw7pMiqAOb5jk
bYslrDbwNRlnXK3DyCjjNIQHZ347Z2qCJ0On2zkWOoqiuiMXfDqnyC2g/CP2OJhn0MlPWIs3dgY6
EAph0GzHXljFLHCrZXY5pWgFOqLxftL1jDtOsUvu35zl//iG81jXj79cWuZ8cw2ehd6i+zVqUpum
MIkaLDJ/SAOyg0Zbk/0gp84jUg3+n6XWe75lXB3PkJRIVWHmnuG9yqtyo/RftoivW5k09PLstJPf
gKTjybyhY9zy21k/xbxPq4Zj6QCChycpa/lmS5C6ub8TRRFp9B0zvV3OOFJoal2nbGfED9hjYmYg
OVXN+MKMS5gcCukmmBNEUa1QOmSo5UQY6+OEPdZjGbV6m7ZNpOvY0icGozqGlrYsm6oCtQ1mFFiN
BSSPdgOd/k1eRspmCRmWspyLrnHeibD5OH665kb86era4YjYteeMyuBpzdLs2rLykEJRTdP2S64V
CAws/gBo4OS9UTBaHznMoY6mlh39mmJhjikd1eL6JjvyM3rk+W4nJG1Srpaeqfnb7zTrX9mOxbdE
nU5tTS34kqWdu+EJ8tUx3XN4f7COZoOObctNVgn5vGW2Icp0hJQW3DVKS2m8og1EmCK4vmXy+OCp
BN/AxgdnXwzjCYyuKn3C8ofyfqnwAoKbXbmqt4VTdeQ4+tzPIBGawCXHlp+1t4/nO/cdnWmgaw29
DAl1M5Egt6i9RM1JtRbPy+wcPSbRxPTv4hhVi151HbkBiSF6+2y8OUBXhEmQCCXsYYYRl6tRBt/3
1A7I+BOypU9YLo0aN2p6o7Yeo3rbMF4js5UYZ4rL6RaqcKbljNI729dhiRFOP63yyEgkOLBGLVuJ
3qM2+Z/OMldgIGOaO2V1O2rEWic3TuhTPj1nNtE9f1JfLzXGF6Kxn+yPV1N0u/OukJC4rEmfAUkQ
7RZHHDPsFTDN/5lWUz1SrC+f/uT1KpUcZCq7J1F15tu0q75VsyFyPCGosWHatY+9rKG7eLbXE+RU
01KcdH1Q/odND8joRmCbCAXIvgzli4UYt3dRVPtRKYTd0S2W0Yi+lfVWqS8hMyeWHjVqDqfsxM4V
8ZPSLiPdbKcYPjh7qsKv3SENugLE2NTzP5ZTguW3G9NYegukuQOXzy3iAWKh3guvSUpwf+cZ569J
Q/r04e019TjH4lEgIr0lGG6/lW+GzC75KpFUsIg7tLbgPgKNH/cfMtbXV2ef62vrGuW++egm+H5M
V3pthQ+gu++dqxxdZSkijLDxC18viYBJ9bRSAYfua+0SeUOHJXBp5DItm1YSGLSmIFHsN5KjMwqF
6GgHkx0ivpWKphhErIJyBC7heLUOhuSJtevGAQIJzc++u92Uo3H/0ZJHfFM7OeUEwf2mWcIdamcW
Q+KTgBVrJZl1AlxEz0KWvloXfvvyFerI4P3O3IeX0OMI2+iL7gnan6QxCa811XZ+lzfPj/oj/gB+
WX0/Mea6/QDwLMRQ+nfxTtAMc6fNvjqod3qGKW5CHsYLuXPyv5CxKTAymzjMN4rSdU470Ug9l3pq
HoiKSPSqUUf6Lf9y/ewJdlm0qudKw4V04BvLv4/NM72My7SyQtfwJAbgwmg+uJeMoHBjzjGo+qEu
SyeGoSMlvPKNPTgnNJ552avI0uxApz+sanUCWBEOgo9P95bp/uAetxh3AU3zy9KwQoSgbKFOulim
aYrqaDsnnXoDSJgfAsGrtez5bymKW9hCnrP8zRYrWtCiGBAL42vV+msmV60QJjewzIoNp7ggjkpk
C6j4tqilwo0t0w3K/WgWAvEVOs3rpzAzASanKTQZs352wMy4ncs1scoaYx+OAPZvcEwLnbs05MCP
VccBw+nYc6R+R6Vkl3VC3KGDwM2beEOlWKDOhix3TBf5h7oAsdna44s1G2KAfC5FhlAcTR9DOu99
fj4UP+vcUjptZqCvK4rDVR+kesF7JfOT5UilEFhS7SvHhXnkH3GnG5cc9QutbiouU9NTL3csW81M
UCTv5Ggbqp75tLCeuu63xIaba/2otg0ZfFAfu9fSkuC9FyBacasyU7eMivJLruk/CAX5wMdAz4Zb
vnYefVmSmMJEgOM1SVJX51tWutiBFi+SACgTfeAfMtF/T6CuLoatswSoZoL21F3lPg3bE7Z9HDLs
Oh5z2e0vpJWhrHljP1UrbdL4/MTwJWv3sg3h16bmksNUREa7+0K99SUVWP6XU9ssNe7pwuf9GFPw
LFUIx/XHdZQbBqjbDzTjElCnjYGGUkrBzQwUNpOIu1ZzrEg6UC9F8AHkg+ItFMmPpnVCpH6O05FA
+8NVdembI+RC0kKaqtWkOjXYV3UfSkCESISKrgzcrWuIMRHEeVwLG4tDfzVfWVAitMldctA6MQNB
A20dZf17PmChXb301cLqduZCCGts+gC8WrT9P23lTAh7eH586mwG+WcYcrJTfF+FTvbGbExYIF1a
CXga7SFzrgfIuXSmir9NkksD6vOw5fBfiu1iU83sSj+HY8XHkyAbLIPtqgfd83Rn7qox8R9nxetT
eZI8tu3fC3fDh/IluDW/qQ4g6iLErPuk3rnPKqbVcfK/pEf8+oAWcuz0rim0/7yuKm6ghbg4yYnQ
vNuW8JtdZayrpJTqQHqkO6FeRcCghnjGXEaIPkdHMntOyBpRQOZKOQSM/WpKM0kcMz7X/mSLvzK5
hEzrwQpQe50B7yDLAJJdXwn42KQG7psBKaptGo3va8BWJ+S2i6lQLjHPIqn2q5OCoXP37A2h/uF7
dv/tSiyJ/vWEOAkfiODeNLaahbdCj38TwwGzAAadmLjtMQQQt1k2T4kfJw76/JJk5cy/jRMkqAO0
CI+qfVH3YdePlSj1tNVNC8zmKyNXnVINfwp+hLWMuEqG8fzt+EZV9zGjjgx0xNmlIAggGx55M1Zl
jkRtfP8j2rwy7mUacrUnhXA7joGIAsxG1dFTW3RZ9//SlE4NyrvBtvoPEeq0NyV+HsFn3jY6H6l5
YdrZsbMUw6VxITh5OCB9OEPnkvLpwuV/lp7FX1h07aO3ZFd6pLrcDE5PyaLru148m7EeH8tBuiXI
IA2nLDxmRbgCtvu9Nvw8bWlrKv81RGMXiULcSNkgh79vsDFgAffVSvIy3KPXXIinL0lnHb3QJ0wt
fm5MwSiZkorArx3Cgt+IENmmnKXyektlhAoohJviWTOM+shoCK4FNRl7/EYPlxcGM/XUODFxvpFq
i276SIc3dG5j3N07k3Q8GI+PaMaZkTp72WAyuKCIFdkFFIXHDPrFFeqUH+FgxUNA1YknyZTkjH7g
N2txtEq2rZfYEuBcTw0v/dLHzsFv8Y+p674+WcOV7hKVsDJscEHBvo8UNqKSLTJnPFwzZIKJvILQ
pIYzFBdyZq8t5H93k37re6CEpPJpb662EX02w3PROmZ+rBSngZV6+X6lAzv+bLR9yp1MOUYb0eGJ
MZSC3kTvWHIr1Oyl2SOcdG90VnwcANwOwwxrWzOF0ry9RS3ADgVAyVtUCJ9YRSa8N/w/gAkr+HpQ
+H3wcUukGcIA+LTB9DR18PH5VORTR3OABOOkyd0YRov+axYXDKGP7RMFP7ImW+ONu+/8CSsEhwbE
92NCJ0SOtuEVmQYHUB5PId+KZERWzGspG0Hctxkdq8bX9AxkkW2i/g/1jH+byDbMzJHXyr/q9QwX
pcCBMsBpeMQGiMoogcwT1zdii7RKwCLGY/N/v3L7mA7Qlt/ZEQyIcDNWdI3/XxjSvU3QXUwi7JRw
R+lmwAIXWDXAczcWxzrvSmtVZPoqaBI1lDFabLbcshaLt+IYM6m3LC9kZOmo1Y+PzuvVr/xDIMDR
gKKUHRn4uQSY6IIAYqywZEbby3Dj2KQ+CfKYtQF0j9PU+I3x8GnR40h0Rod1RxsXB46ipLoP4X3R
AYc7YbZWfS0ptbDwh58tM+lcBgMfQD7iGm6BhBrKOfXEL2HwZ9sBtyT/cQxWRxY3PIW/XAQzN+be
S+xyCY8K/u3eclPUMNlDXD5bKr0FW43WTplxu27G/JcY56ubyM5i2rUU9HpCDnj5Tzxzu7JlF+iW
LtYltgCOw7uqU6NUZkoTBuZ877JyiBLCErbyApOZ/AURPuBd6MVcWKYjmGIHKWq+pra4Hamyuc22
raU1/2Iwb2FYkpa814SEkTbgAvLCtqAvTFDnHcyjXIcPvdgqWBEMB2I5cZxjso5udVaClc9zhcuK
PhDDp3jhyj8pyoH2z7+BKcAku2MQhw2cLXTeBaqaq4qngZ5z0K+SdS9l8nvY4nZ3+X05Rvx1q7/F
ZFz2MVED4tuM8RWzfYWc93DvKlos8lG1bNfV8HbqaksNqc7BnVaMEgAcpQDSGtCnWlfDA7WbWLZ/
2VnPRzP6by3cojv+PGS7/jWYheTyDt9nfB8I5NodYdluLvcP5pP+ixW7z/5Lsxt+59ADQtXGhs97
aDY15dh5LJbOYI3E/reUXM2nPGAXk6mbNTPNfdybwXa1Kl+kmiMHHyLTClWo0UUSnYqMtfAIwP7P
nRXaz0YVeezwuaZf+b5nSkCHvfo8JaO6JgvYsNxSVLbaxrYM+2Gx3y0D6byE1lBMCkQDSG71pBLN
CNem7aKvHAAcNZPlfgLf/uFKMoovlhHGvsa3zQgLJGN/7fAu6sSakUz6yhrcLH4QwJYYqTV51Yr7
EqbIRAn4npfNDX/CdcvOmdpi6teDIsdepXTmpG29y8nUpR4ExCBmn24vPi9cjO57Udlf3gLdaKox
Dv00xjnWNPeLh0Es052oH2Xikl8jGijYAX23jGaaFOtwYupIXR03SkZQZ8aDyZZk7/q+7ADfjZLq
lb4Yk84h+7DWh3zuZkSYPZfCr8DKsQAzanD2gANJZ9YHPBSjlE3RTmKZRBnqJAxm1UPoI/ZpxQpP
Vhfk0Z+/CuplQPivXGUIuALEx5+37Fo88gPd5SiXu9hTDUVn86M8QIePzcd0V0tpYB5gf3KSqqGO
LMzbcxQynFpwNKXjtbdiKeBhFQ7h89PcWLGaajGPXDqtP3KAhsmqTa1YQZdZACprEhgvAuESEG7L
u7ANfx3xBEC1qR2f0XEbiQ3cVaPWqF5RZ+uTTVAwucNaduDk51LaIWxtUFqJnXpm6auoblHa7HGh
Qk9OrYQRw8Jjf32GsMkZYrsM6eB/7c70mmYCUuPvTHTRY7A7K1GRlaOTy4l/JG1gGpWR0g0R0TJo
qxPY8tExv/u2/wlfWPhNZDy3E8v9NHN0nMANA8FC3qRZFw6Ea9Sb5eep3nnRkFV1/ObKSHvUNXWb
xWNQXrt323QM6AM+CAlvGEOYnBwcFYNcqN4HgWjaEJoiCZcRSzMzbdooFM4HHjC9QMl2g/PKAmgY
dKLvx+ojNXRMtjAqvHGTlkR360Z/aiY2icDo7pTo5pRj4TO0Gf5Ll4QRT93Y/2OCCTLfd0jnX6p2
kknARMNG2jcWg2QZL6XIajres6no0hJKcWtKQQIe3bBmZ1kmKAeAOK/i7KFWR2aaTh6EJZJI+V4Q
GAWiwjM2wdcz3BZmC4iKHp/j1duoQ8S7FLHIwX6o8BhUuX8eA2El2ryo3LTmyJkN8KjvA5WbMyzL
DBqGPBA4sZz58yc6i7HVMN3ae08oieN+TlNsVWOFhOz3iyLyp/IYmn1J+o6kRZgEFgdHaOpmLbyI
8rrwODdnUmbOwBOG6/XfCaCx1vNTc6RtOqhaErHLrAtnGFXT+gNGZ1HrRTa+f1Pn7In1V4g+lqhv
I1oETZdjsYgdeQZoNkthjqoWOdSlzfulM9jkO8PuM1PnCqhOav6sgv6dTiHO9lMbzeDs30S/d69t
bulGAEdBjtcqzRO7vyK5sTBYF4rq9fq+3AL970WAGsAJ+/vMeX3kRxHnrBIS6Q3PaqqYCDJ+GNTt
deHGZk6n0s7itsqskjNNx4n22MHENGfiwdbItoZgJpGoOubpcD/esf72DTNNoeKKaC4wx1dHj3MF
sTFR02ToAgHkRYzvmIhufiAmApcxzOnb74lJdyNtbEFAdscC8i+b1lnEs0tBKuyCWvG8lGIlaSmd
WC0iT/MfxHg1aTDBOKQOsLg4JcdzfBgRrQtQZHYOSH4754X2ZAclAr03EJ0B/oI3uadUa8Ocvhmv
KRfWlsYy1nOoLqfSxPGxraHW8HunblWt8xahvhH9rlzTuDMtfMv5S23iBCZCs7wzmBbkSF1GANnw
We+ckMfvg6EgaGKImZcRpt6D7Fj56k81ZJP8QaKEUPPmeUvE0VG/k+VoqOUK4r5NhyXwgm6a7Yn1
rw9qEAp3FvGQPmGlDg5wMG21pbEqAbvFdhr3KUzQgJXdvc8JHKiz/JgkcF0mHaj5ZmMoZy9v4lt+
CNpzK0GlXaS75CQe7eJdAcw9YeNsxy2Um0uHnqcQk9Vq4kD9Xh+9sIPQlAeEvuGR6GkGEsSFFfBF
p0ASDEcTBstYP1FVr9YFU2sb807ier5DuNjVxeN9Rgw46YYz+p2Id4dEEUPh40w6ac+fihHXDJz1
MrNZYz/ekeTZEdGKt/Eas1OOYdFEWNDM/ToK81osT9cBcMgwAkf3VlzikvLhcN6H3xxhODm+xStz
Ws8wOKqrG4HK3eLff/2T7s50N+EWZWBx2kibD43fZ0De8U6UnZTE7CdGjxx+7dsbTlKTSWr9XtP6
W88Qq5LsEaQrNAg/vIRawnIsDyNVkb7UCEor7gfq16B/1Il7hyysTSyLS3rNXECjprfKpxKr5Yav
THiI3xCjAYkdwuzYfdMpMBT/GnausrL2lPF64FkSc6OdLSrLZ3vBrAxLO6KqFItgMxF9XnR21vJu
5GG0BSdZbk+lrTYFuIIlhV2d3lXB1rtGveaEzOpJ6QpXBn9+mrhxjrpYbw4Kk0OqFlF+ZNxLcIKz
5YRS7i4Q8pfdZgAHFBkTo2yElQ4HsVx1oyr0BkOlFukRiS/Q3P096y1AZ7YZ18ZmCW3lfemVO4J+
i8pRSyY2WZnbDuJ7M9Hcn66TiEO8v6lCblLsV4W3X4qvcV4yKkH67vRNtXHseEvnE+ktRgQ5i372
tNSJ4gs+NQqqHfC69My+f8dxY0JTx+6XaEUCGix2aSqATOp3YbdDCG3BWda0kC44oSyMFCxTQ1y0
fzKsz15rGgw5PvTEeQqQyZHwcq4NCKupncCwA+oRVaSxXDJ3eFu7zCDfjbvRYTUZB3d3DRc9Sk7H
/mCT332e7tOiDACYrFeU6JYtAdBqhMfCorzM4xc5F0C4UoTBcmat3CH/WuMvEMSwkrk7Gp9FzM6p
x9cq2lFTr8guqgnVy/JtM86VAdjcK77wcd2WQl82SL3ReFrXgCPLSNAa9KWer+jezU4+fF2RV5kL
xYRzmpKRBBpkv23y+yI+mTHotUZb1x5sqKLXne16+BsRs9OzwAncWxwDulbsgQnPETZFJM+px5/8
N2+rX23baEET9RdIfSHGHYmfTI0niQaO0zAXM2xMSDuBrFmGYAohP1Oco74NDmingZaCte5q4ICG
Ibx24ubooasJ9SsZulT9iJoqh6SVu5oi13jElnopfIROj9Tyy/arjLvHL/Ql3nsI+sTWvTvAnt0D
xPDsny9M4yZyIZLa7KfUq135lzHUX7vK4q0mWr60Xl3HskNbLmgXQ9mTmneF+ZygyWmOzeB6dV53
uirfgDcpL7RoGGd+xGGD/ewEwJNkDvrVYLFFjD5+lzLfRFjJnt5W3/7F170kGMdpHTEo9CmyFABI
9b3TBgZbTkFov/W0TwIeHWJWIR8BB1g2ja/Ay0r3n5dCzaCSAgpbrS1aSMNt0y5rDAob4PCQxjij
jdP24yukKz4PiCo/u3VLuh0FjXVdM6Lqlc4EwyC1mL01z9NStC7v6nCvz0CL/VzWaPiChx6xNqVU
2/AWwEGEtzzE9hyHBFdSkvJgVQNBaSl5gVvXiME0l0jCw7+UQVNqvFQbsMo2tHioHP3W+jzCN8x4
hW4cyD9onvBV9t70ShJbLAcnGvVKiVTPvnfXGnnrTAf7rj8wOseyOVKhCfH41f4CaRTpCYvX/bgj
3Q64f0O6MsN/qJsX12H8nFRdTwredXxKSM1wAPA25pFUY7VFnH+P4TEcdtJy/QlmQjW/jZ5SxpNL
BjstfzihJZwTLiisNYsfqMDxrJAUSGnBzVVBbPG+7HIRGIsb82W6iVZV27NeTsTcN9gIoAluILZ7
S/R7YJh4q0ndvBX+52RkOSetf5nEvf3W35cCXTlkRI2Dxf2dLke3pulzvId174rxGOv27kQL1kBE
HfeUm0WFzKYx4b20ke6F1GWSxIgugOvGmkczfBdyke7t3Vo+Cg8tpu+P89IGccTRd7+o5jKU8drH
kHWdUUDQr0YNlTpLmHd7+5qjRblgoGHUn96B00fPPneG5qei+JAIFr1xsm5+FUg+ppYKG16Vgb5e
/8fCTZ+fPxMU1EPV43IZplhtNcyDP5HzoM2nwv6z0CpVtUSducbHL8vtitS4t71v/Wrkh8MLSs+e
FcjaIiWZIXlMCBgBRLgtPAWKS7vXcS9mPt9Z+9GzvppJkZ0S9RGiXSvtkrVnC673JObC3RZ5DFIO
/4pgM3SO8BwiJ8wUtBT5o5HZj50Obyesj/Kw3OKi9ps5w9wSK2O/pUUeRfXDm2fAjcF9Km+pohi7
PZqMnddYK9nUBzQaEbAhRvkxuBCht6bkeTC19LAKlOWFYyuJNo8wGwu1pTZN3xR9bBrpGleXbTxD
ZMLCqA6Sjh4CEPol0xXVyl/nYdfXPeX8fijSuFjcf1TxlC8hIafZBviOXDCj1xufrdbZUX4rbEqf
VjsmY1g1EaTXoJJX1bkTxwkTMshouqq14rDjOyTjQtGkJS+8YoC9tFqO5CI1n0Db5C3hB9B4FJSD
oihNWNNy++eKsTb1ywyopTl+hZOdCmsxCjkY4F1lqk0SW6cJTlWYSiCQQf7OAD+y7QJUMUtvpBji
EVNirTjiKUpMM8Vsnn9VVc2rV4PptaUKwRxkliRVAlXll84rWO7juP/gIkbRILJox8B6AVTOMfGv
uIpV/vSkEkTDLju2G1YhnFHCZ1Q/A1CGsTeI0Xh2/QlFqnsthtUL5IWSPSRinvcmRn5+BN73VByW
0NpeXXGpP/LJVc/i//K5Ul3lUxbYEE9MCiYhCJcgZpuh/0zEfbwEncC42iu/IRMmyIbbTNzKeXb9
V1Z+cPaWIUxH9uSfNBclpJKF9SwGOOyzx4QJB0qSuimUOCOeYHAWZZnWKQTQNhrkrYE8l78JrmCu
ChAY3OYA9Ea3XjrkeycEohCVkIjqHtUi1OcSmYenIds3E41+//ihWeWPk1cfFs1eIGmQTfNDG5WT
LOUca+mMC//fjx9rExaW+SuWTJUu2IZrX4+vA/RyFkFiJccq6kO7NS9mbcs8Sh66MqyMHYv/M6rl
ZcU+plUTWQRZDaCuGedwtehv3rf6K9Jlt7plgvhZBKWcEjIdONdfxyYzew1cHRGO0A8elXqWAcH2
RKZl99kpxtIjdLjP4pp9qYDGK5tJcj9kArET7kKD63NLC/SCOtBB5BP2e2JAECgQ8kw+vwdfCphX
gCourCryKzvTUqU+N0HJouk5e/a/7tOs9bs/0EkjCoBVi0kbMPOtlx1XY0NsRe3a/9nlW8TGASJo
TbtOJdnZgdoO3r/GxIkdHhQhgb5i+0XSJ9+CqfQhrY+CjofvfOOUFN0JAkQK8WfmI5hEuSXhMSLx
RLyFV3apz2oSOQLTMZdyTJTnclVuk7CTp3o6fTIDNIXwK7YI9HjYGNs+x0EYXYLqtKPKeRJCFhvO
/FI4ZZhbEY1vtdM9aWuXFZSfZ2lsEUx/zBkptTJgw/PVCdafe0dKHKcncp7A2/sRPOEH9Vxz48Fs
VKcsd8560V6klRaqb9hf0jJAH1gBnR8/d8X5cFu4r9UpiPUBaQveq8zT4zljlO/5ateF53SYO+sX
woZr9/KHMj4kyZ3HA7JrNrO0OqCUj4fe2HUe2SPdbNBppJDoyx5fhwJWrkAspPK6JmOH7X9i5wgc
ldlvEoYTYLJSUWg2n2AHBRuI7lyVNTUWrF9bwxbdoJ4rBeSModoi6hcYgOcR+Sw5LQEyZZ/F3u0G
kkxOwSKeQNDbDse84b5PoRD5tWocK6qJv1V+eqNKfmBVZGfeRs4CLE+2aMq3ovSclogwgTqF5WuM
FxDWxs8iRjsGcCdvHsDaWZgRRR55a9A0wyVSwpBf1yYQJC8DRcuPGIbarLH9le438NAPSpcn/S9Z
f+FEVac6B0rAw05IATyTG7Mzg+z7JgeCtj6PhcyOkRxHx4hUT0mraqXtInujxLXUtxymWO3vVrDr
Cr3rTsbuttDltzq2xojtNA/l0rotpaSgdtE8olb2XPqbmc2lI4th1nMl8SR3L7lb4NWrMfR2FAwf
Sbvt7nPCLaaxmTGZ3xUVj8tRXwa102qXd0gcC1MfVm1ct+9TJj2v5v15FRmC9wazeaInzdcl3u9J
hZjtdP2LaEIA9bNtGMqutXkFomrCrjtV1XBEzoHPnNIajAQNnUCFyBUl7rF1KHyayFVqebNvwQYM
MWFRhfepuYsdXQ2dcGK6Q1bJcgPiikZSBba1iCkixxLyXVW3ZJMyXfUpUvalAvc6kmB3bdDjNLYC
9yavRyjjAxw0cql65eyKnd4wm5SoML7TAEEt4lQWch9S3A95dHDrR6BwZ0beIOC33hZ9vG7dfDpt
20+cCwwDghUVwLjHt3OVyIQTeYPXfMLGHjIpUhFFWDbtHGgHuYgTA9OU1MiAoBpRJsOr/2+DcQyj
EVSypaBZ7Hz9J2+RCyWtHFBGWktjOKpFhxtPI9E4Amsgd2ciJsjmO+ZFuigZ9EE4zsHMPqM4kzso
DRSndnJWJhBXOjFc0ZvOWYuczPmX7CHByV9EA5kjmGqzaYGmj6a63/VdghPCs05dVVGXbd3osVIu
rgohPFGCLWD2wrtHWIMGZMJHiGzpAhWotE1O76OBuXtuzmvlhM87OT7c+xN7EUhx2fwepCikFuhX
d5xlr9haBnur2s4t2MkWSu0qJEAgXBlxo5+0NXZM05wsSBqjiFzMuc/+GofBj1uYDg/dcdRr26gk
X0SyXLav/OLjktRCXFZwptEeK7qWhB7skOyN+mBcqPhrzDA0SIDBx692rfWPs43qPgqRZPSs5wyf
qS7XLtjapymLRWYoxRYD+GnVrZbqUoOAmk967WBRh7uL4s36UCSBYqvR/Wgf0ESJej8QBetG/3Um
tr6F4x11YzkwVvMSYo8kj5DSFLYWCgPGnyI25CVg5ywjldecZt9r547z73a7nL0o3lhcR+TApolC
U9BxNVlxkUcX4vetK6/1RNH4PxZwDOrQ3tnLSv/G1hhzpKq9DmcLnTKtn1RVZX4eTlrTbDpKsBDl
7Jl7p7PerYYE3a7fuoQt/BTscQzlk1n1M/jeVnPLym5VV8tqeYci+hHqFJicggGAGzCBRQlHamz4
HBI4a6SmD0pA7iVS8Z7nLbL+tz2iHwj2P6JM0EIayM6rjeNm9CL0D9nFzNNT66wwoyT4ygepBEKj
rvk2GcSPZVCjRJ0vAsxA2145NElTw5SgeYq4mF8YHyhLZaZNjXTGh9ioS4T/2sE1PL17v/jJPqHN
ohwhbeZhXe5E4rTgEVH8GER1fy6xp5ETGbz/kT9rLYd/ghBBYU+IjD7gn6H8fD6M1ja1JkJAd+Eg
uKlBzGZC04iVtPiqtHrJCEoDUGItqQQr82m3f/SxiJJcD98TBTjDZ4YIa+fBxOCf3XdDU+mgsqzf
lPHK1d+Tgt11JRdJWFfmu0LyfjkAgXOcpuVvAz0Ec4OtT3mHpk4+dCMqvDRZam0O47UMWIVs7awt
m3ql4xlC4Tz8+2k7v2tFsLV5zIQHutrCaY0EDSaHYolIUzVJ45GhQvgGc6ozb8Ost2tgbP5nIpHX
fYuU77y0JEHP+F0J0vk5I42eFf3I3U4JO9uAWhsIpxIK9ouF5OHC0kGCd64fuyYai95YvI+ByMwp
GvY0CyKMlBSaqu7zA30rayi6qcBYBVOjjeInoUiMWbhmAZ9skjE9TP1M9bmepmSqfUsgAlAmrGvh
sW95ajlbTjP36zfwsmAXW3JRul+csMlZlnvH+MXTANy7ejVsyZI3J1rXZ5yVCzreg2XBuXFhIJJK
zHEx9qwavXVzAxuxi83P/uHFZkgXek6kxV0pS/Q8ZEGjWq5ZzQpfsFCtRkJtKWKFOxRKWg4VH7ii
GxDFGJG6WBBf7T7H1MeYYmDRbUAMaeSk3WWuHRS+bJ1AakOJwzwMIwzz0muB0wbZtRHcwcDp+jd7
bz4yx2H6LUWFeRePBQAX1IItIaCw+5RJb+y6kIZ9qWhCMD/K9wx7WxaDsb+9irsp8MWfDLFsQWsO
PaPL/XPTillz7XY8gFgzIYXB83/iRPaJARei0ZvdphvSkRIDgDUcflnAfHgkjYIgr73WfTBtFvQD
FhnfF+YuTVYq1mttmHgKkCwedWAYREJIz4HjV0sJ2pMXIuJiyVwLt9V3zNPd8oP9z3Rh6hITlSGl
Mcy4mB0hoNQ78+OIE9H6/rc3tBnvfV7OdOLc8XTh3QyKu56jfeIXUV/EPBlVRMcRcVXOJQH1P5B5
r7iqs9vhVh98rAwVIbpJ4CNWdBwWDJJipTD6+GjtiVb7l2tUaGlrEDyy9Bsye3z/6G2SDuhsQ/VQ
Qpa3IVyJX20YLHWunn5eudhSaT39KkvShPFLcYAUpyX0O5O0vKV3TUZ7fQ2INTdinXZHEdnVGp29
nGP0r5l9G7A4NgOpu+c2l76TV+G1djLxqXOb9PkuBUEbSepm8DeHL5oik6rPcGlAnfyDEi4RV4/R
7mWqb8zzsRS0O5c1dLKPoKzzRBEgf3+Lf9vEdhEiXaDm+jfcxq1Uy6U57iuY8GvVVx2DC4pQHgqI
xIcY0WTs076u1bqlTlvQ6gOZgvZ9oDwPHRxfaJxwPU3uCUaNZ7ImeLPyXKk8VtWWIFHSvsRYUHaD
eu/u8S9aBIoYQB74iDFSYEBQRZnc9MhuSaBIr6H1UQGypb3ov+mZqpopAkZGgWBmZEh8ez+3MY4t
yeE4SxuER24B45TGQBN6HVSqIfn8gg0GexPGqJQMTae6q+hMDa9wNqEiy4xhWqzsYGst6+rbxtIN
/qfA7wEE8fdply1CPkSoUvWMAlY4pPLNt1vNTeXVgukH9HlsnuLcIQwce6ZhJNmY+NyOd2somCQT
EAlMsgXquy1yQmjUGTFa/3z3BUVza0v5Mdi91F410tHPDdXG06YaSrm5Jv73+nFSAIA2CLAOhHWp
Rqf3h1Q2svsCBMpuqzvUfz8XuV/JBYziUNatDc24vy60GWcUP+joYRTeHJLTN+kOXqSQG1ypoLrq
54mYFOf4+EYX9NcorTs+7RWRo/AzsPobFG97VsLYei9UcSvNmuKaqgRvwViTvP+IheTkBHEpOjzK
kNZMDl7oBDwmE2kdQyE7G7+S7fT90RM5STqxcIR49dn2eXJdDobCJmPg1xPVUf4nBfHa0mqLxXMT
DlDoyd0TDqJfdYDztD7jC8dB2uPVD0Aguks4gJUvupBZa41NPrrQ4uDCvveTeE7OF1TVWG+K9eSb
vhydR1DaPu43+uZxq8icm5uF8UUmaBeV6USYl3zgufF2dKgAa1++aoTTb8fOc6HrDmzd62fAIDvF
KPom+9nrZQE03krF89R9eTV1Yakg267xMacVNEwCmUWxcgjOJksnnPfktEc1uLjpK3H7VJZVQJru
e+UonfrYbD297Pek9p8ktoTDwXpeREOZ91O0nIRG0MNPHLa9wUFxFeBzEt2VbF8dje1GyyApAr3x
uWsjUd4Y7TY+91qDFy5mLGghPwktc/qNcAZ65cviqEem9dleTXDmcYzlzaJrt7jMW9gucQzMUGvA
7MvDVZuD3+COdqeVYJPC159+A7NXi/yqJrIs9KVsBEUsp+FARwiEUgeKwQ0zRM2fFz5MavVIZfRb
9rvkagUlSU2Xh6RZ5vdajDfJRjeoPI87G1mE9XhsbWqqBXYIlgInm3B3fIE95pYL4ymKJLcvGUxO
6Cb8KYlUazs2hcpxzzMGPP3kKHnd52C647m7BzSMnatEEO8RYuUtRxaLYxzZYlWXcXZqDN9C4KwN
2wxox15jHm8RUYgzl5alHl0/Hf+UPmPRRQ1DNhjS8vKs3JrGdo2VdFahIsFE1oCm76XsiIvxiaS5
hpdYGEbk3pPUvbRCqGVmHNtlzjl4D+Fw9rjilNVKzxmpp+XuRq3v5pRapxcgazXI7/nNAeSvBbxC
YW1iPqGnMpJS4P612v3Cht24tEZDr64ZzVkEg4cqnyHyyvQsYNzRo8pqFcGqkjjblDNxDaMHD8Xz
o7v9MFbDlGD/vENwxqm+/XCIKoGziBkDDkeo5YlUqlAL5zsTe5dbgVaRI8zHfkIqQpCk7z8qie0b
+hSU67ulG7FSpnBDXx9Zm/svpmFYMzsqIIGOx12YKA1D+FHiShwbaQpciYs9dn/lIZriR/Cp26/r
3ypk9BV43mgzzuTv6m9xrSAoLbP3+6LqHUFwuQiAXO1o9nppxZSr7462wsJH2JRRoERkjk/V1hpB
3pxBW3NiLK9GeLzLatyzXM/GKgnZRE8aeGjJFMFbGinVAjiJsnhVM1ck/YFQ0ci8Hh5fNuSSHc5V
gJp4p46v0jRvzHEGwx0a+UCmXu0o9HvjAbadRUTuWTQxa+e7pkPVZ+NrmlfZjpu0SDMe/fgoIdEd
sdunzUEOOu97IpAM9UzItxU/hNbP8KekuFIO5XkaS17CrGRnjYr+8549NcsO7U2JNKGK/DHzCbqx
sM7PW2qZPDFM0OqPkjlWiML/n8F5ka2x82eM/94YFwZPhnSzY5DXeOsTi43p7j3+jd1k2tgKNfR0
k7DUsE3Du72ElYTmfoi5eQkwPvtaPtqZIqBGmwVaZzjOKU/fofCsAPTeKl6xJU4KDtl+wU1Vm05c
ay4a9hZ3ZxStlHw9Vem/jmMJ1SmtEw1De442/DIalMBdWhMfi9ZN4J0AZs4Y9tqc2mTJk4k3hUTi
l42HsMZ8ybcgNVb9eUDAAELGGARLnRhLSNjGYUzoii/jFS+jo6azhQ+iEYcfwksqdzwVJiML4qBv
K1lY9o7bu/l+AyZ61aLi+4wMhXD3mvNBbEh36U5xelqzjsCD57/qZ46/cmry/Wf/KLc6k4YdcQCe
EJQr41Hhp/4db2SPWvLRgQNOLEmp08vhTUMlqrfjWvPeoN7Dtd92Vcy2iq1coiJQaUmp4Gs5y/Vm
QvECjclcAb4Uc0IWKInjD0pGeWLkAl5OsiFHdZACMpfKp5kUGC4JnWQ8BRt7eCJM9D8apCrO2Gl4
dh9jhqQOPkjgGCrdMpEh2fVGQLOMiMkMLPgOJr3PTg2FR/zfJD6TEO5W3HRahYiMoCqH7ChXKbRB
FOSyy1CEryetQ10pDDx+D9sbJCKeDvuDqrvQJuU6zM7Ihbq6oymUKUnIpwWHjM39IpvlFrNa0lOq
AJNwo8dAZGo6vQmByGN0/dEr2RdE7FF9PwWB+GZ0CxNXDq1gVUVurVgzG/YcLLuA157dItSinOn4
M24ki40dquNh92KQvtRFenAV6VaxJfm8/QnNzVz1jLSwP3LsqjQJpUTjmV5jZaDbHeBkQvl9LPMA
wKnHB2U93Oj/wqySnDrJ+MhF6YPqPX9HUtn3bgxQ2OSnMjnJM7dB1eVDI9uNImcmDZmqG6MDajJh
/6Pzus4YfpdBIK7gOwQDHLFiXyUmqC7qfp2/QcPmCKBQZauIvrBkJ5fD/+RGySh/ss4ARKHYRWSo
36t9Wb4OzkEm7GH2Lng1vZkOi7JVQm/bD5IsAKsUJ4QEWTGtfzsneinfzbeB4DtuBCigN3y0bEQL
IM+Ox9aVzSItvcPqls9mtTAXP/Ski99WRKOi3Zjp4+WGwQGDtRWeJIMvB5RsCmt5KE/vZELzyo6r
uT5jDZUH4Rk4/F3jSbrAi++s9JLICdH8Fdc+1HQTi5bZSgHpbh3XyfekgzX3KASD3m74DlGFx5dc
I3WbQTkp4L/N26nFtgRCgMiENjxl2L/BkNC4HZ32pah9CEfeotDhywdlnTHnJUx1OSQvzjHlWmDR
NcJfn0yVX410Mk1HRjyY4au4JKZJ0PZHK6iYsVFQmw70rOppW84zGsvgq3s33HyjD9WRKVK04ud7
6q1WOcS92TggKkF8yalmwOu++UlJWdU41X3ZL1B7m3pnrqIe1yoi/PWTQ4BwnZj+4WXELoYR5ZO3
1Gfn+M67KodoprRiD8pDRFlN0jZ4qrQtgHWiuyw+4V/OXd+lRkMbW8LZ/Crp+OenLHF/69L9S1Wr
rX9O9+rWjclpzZ8P/3LLtJjw7BBUm/HlmA8t1iqdISKlwfKMBV7OadtdxiMiCJU+rbIdg0auTaZu
DnbYLwGV2Uf1f1VsbAYj7o4HHBaEEqQcHs4QgoOMQQVEmLqz3MVA1keY6i+AKPc/gS5d6cAF3fNo
ojOzFRKfgladtZwThAG7DYA9hZp+77K76+FgDsia8juNwU7JtylT89XZjUDSoRv+Qc8UQTNO+6wr
yEgctzeEdn6xCapgKXd/xogjzcm8wHMgCQtLq0uRnISJQ1tND10N5xlg/dSbdYe8HoXn/MbELwdu
kPMUb/1WN+JwikOQsxYqt9LJWsB6T0lzBke3ULTHlL0IAPdj/LyRkNWyy6/RCUelDeh1sAx2OQZD
zo2OL0aUBl/tGO2fFfijucrkD72oFfS0Z4W6v2zWBwGL+v6uUZg2SrQXON+xB5OIhOgyk4ryLvAV
zaOhXBfa8s1LUXQOwVoTHc1pi1x8bWX4oEyUYxyrJRsUXXqrE8KeMvqQ7GxLDq4VRt/jAo5bB4LX
Y3jngW0x7hd09SnkIkFqL0AUYguT56sVxbtjpk/TLlIM91ZeDJt66FphrXNPLe72ghlEoA/fjNGE
ipfhWBg+X7eMAJeBSWepBas+Vei4gprTyMsNcBoLjHPrDuqPY6b9FTmUm5Xd8Xhm55Pgf5wLBmqj
+fgQi/RfhlDkqZDKQp76S48S3Ax33H7y56KfWgAmEPxkpDj1ca48ytUXaddyKf1PEd4UtixKWxop
i11orOfkEXg1H0cj2+ex50jde/aZ4Xroa90+nodTc4CROcrox4Ry0mjyIZ+DnYKZcdehmk2GEh4m
dpknlHPyH6Y8iEEQlmAAlmY/e2Sg3eQe2cCO1BF6jIiV944qzoDS7y0uOp3XPU+ruKqnB7fbwJff
GjSUenf2FBgjzZWATeaWj8IffS65Cy2znMP3/6gb5wiy5O33/qFLCtMtUIFEru2WdlhA4aFwfjiN
oarjZ+qBlMa8NTsnr8+RQKAY7QpwmQd9J0i+5LpWvPAHcska9zr13iIs5KdiOOZBJj4w9AZ+lbr6
sLNHInlBW5o4srJVc7m/qhTU0/8qMm5nwGqIhu+/pcnPi1B9DhcEASdkyZRarOZKuOC+QyP3VWVz
fLrW03/mOylSx/EZ9bOVxrho6RjBOMXOqwlGy8sivJ5X899qEnYLzIe73FLA5zbi7/xHnXypOSlu
oko2JZlNm4Qy3U97AdOJ+lw7gIjQsaEgecD52fTxq70gM0X1Wnvrd0gfl2A56BbY9s/iOvp7E9Z/
JubTcHYdynkfCWdj7ZhuQF4rnw2j3MW1wgI2sosJuFZ1QKUYEdfBCILse2hTe/r9F1aEVqQv75Hz
wVHIirWA/ZGpI6gn+gDoccIKnW44zQcwCp00cNlxrf0fQ6utJrD5UIuqITr0dmnlIJMzlOEdtPf4
YU6y09EjCQJ35nCe/t1XkzXa4M0/ZzHbrLqHrcsqqAMHMdc7LzWFIaJnP0B4nElB1+3pcGRbcCoE
XQwa/MauozuI6V/vmrrbiDvg419u9YWSE/98zHyRLMDB6YYxodCjEh/fish8mgcwlytK0kvcsbnz
5fNm1GiWm+eb3jtjBZsJelJ2wDo5oq4Py1rRRr7wBalRNmLLkCWakY4wy//ll0OT7J7yAWQP2C4L
cFulZDyTIaQdj89xspjNKz5nCPuuOZ74hASyXM4uQLCh5TVswDzfSJ3Klv4ZBJeQqXNVhO8NpODU
Ab1TdQy+5bvgCK6B2r8eVz6X9t3EqErTbKXVRwGyBTMuroh7EgR+SLQQoRLhP9pMhCjHrwIUrZir
5pYpZk/bsocLOc+HwB5J4MybkyyM9xZpfjtiW0TDknoJqTw1I7t3jW3Oe8sXnZEfT+6pwhv1WiT6
o2PCkj/ec5OE62OI59PDb/uujq3Y7wbxfD3OwMHbu94WMDEz7ghAhslLdAusBxPAy4E1GXMekiIq
NR/OtovnjEmCJIqtE/ZI5GSuxZWuSavEI6e3jbC1z+1uVHUXnSbU/CQZj6C0pEMORK+I2ypK4DPm
1/toZHe8UQa4FduuUAoMfgQWop/+sCdyxNovAzkXdHQiqWIipWxFjJ0cE+nMQ5AEsINe0kXsJI0D
8v+TxJGvGc+qKP2SDwpWBGTL3B0RDcHZso9QT1HCQD7x4syP+eJn1YXcKNXarkOgfOqwb4gUXDKD
lyAb3ZuWGS/MBiCLd+ZYhE5tWb0jsckKr4wSgigjna51tRcZC5DTU2q1NnSG1yIJWDg3gs9Kd6tU
FUi6N+Fr0H708ZwDgRkVLFyY/Q7Z5zH7X8zzXxy/a/nitbL/N8fTgVxtDBYHaWrRU80wzrHoc1O0
NUrPn0pP5T5rLSSBIXdjCfhqvu7a6/YXon7zrWMJ/nAU7I0+iB2awDP1fc0SQGvb34E3FZ4eu9Ly
L9DfKb2v/5uP7x8Gv6QMi6ft4AVf+BgMWRZAEFYFo34XyazDkSoo3qTMIcngOEUtm0hd9c24XVu/
HvXGN3KcYW3g69PLNiLLvvAbLftgsGn7kA7MmnxCEsfVFjMloCTeg7qgvJt1Kh/VoGA721/PWmEB
/GcPxfG1/1RKREGYZ36bTfDYGcaZv9HjBIxlK7FmKBdnZlmzmmx5WkHaZqzPBwavqX09fETl+7ut
ZtibxrmEn3XHu6JV6AN0s6cXz4I5ERG0pyVG3/PHXRDIVguUjc5cgzwdEGnMsB32K5XmknEZ7qR9
KBU6oii8Tb/Fhew1WW9xigkGfc6ekJdUEEAmxZEvqM4RMjafEWFBoLpXePsh1x9o5s97NJUFCC3R
ZSXuA0U5808eYlw+ko8X6GEDZKHoen48pozETBGbs7rV3MPyuq585nywhAupsHGrzoVhzop2rNDo
shn7/ed26YVgb/MwjlM2k/B3VOXIxV+k5JXe8zbarGUoQNi20zfslyNMt1AF4NErlPcDve9CSDRR
FSooweCOCmckg2s4PlN1M8IjJrqbO6AnIhahuBkcas2tHj86pPIAWbZxoZ0vo/x5k8eRrJe1AJXe
2GsOqwrvUqFXK2epOHrV7wQsJ9fvYvGNzczTvnD56ip/NZQgLYECUdu5r9QqRsb6rNLzJxesso7C
02ekfMhyzlN+oYsg6GDw+xjN1CYa34M9VtvLkgeKdfdfrBq+zFjcdKnAQaitDmPMBsJ7mBbbvB7n
kEReI76/aZgSjD8qw9mBqdTgfLLTBJx/atkkPFQRGzkSogejoRQ5XvcMYD7mn0GTnWYlBEkbPa/Y
oHvHU4cDYfvbUxijmNE2w9JHeumRJkQQIZ27etVSIpY9M3cWfwguen4alC0wrMRPM2QDwqFDzGOC
QetewSBLM5kPErjGVV2MHkBejMUgKljJ6m6DgCsGgBIl+8bmFDlgb6ZHxkpq9B2F1ylxIdBkRZBl
Z8RJmjtkSJdU1rBkCDRMf/yCu4FYbNmi+4alWMDEAo5W9UO00nbrqDAUh6dCda9nTUZr47bADJQi
D6rbsH6zX2xDf+ChM3uXOREeXkTjCQeSJehLiOkpW1etRvcjCbqh+cs+l4aVl7fcZ8V85QD6pc6c
a2Mvox8mixGJkSzqR62fAxgTWzNhmbypXRNXPxVmKHkU0InjXXnhsfQtKHrE8+UgBvztyfczw/WR
x9YkgHuUCvQBVTfGUhdZjJcUrpaJmMv7m9w3hfuBdhyItje9rcaUVGzOozQXlG7j+zpT+e2o8MnB
qLNyrhYFCJLKkOQzewcv6dMgzqa4hWzpUkOQYhS93Tk8gqr//bjFtyr876XsHyLmDX5q8PW5QMoV
VoiTaOgvWh+k2keqBw4LRh5imXHf1r4PknLCJqT2x1tctd/gy5tATxmqwHwVtZX9iC3CWUoFii+b
ZuVfBlA8Ud2X2VIV2idZxXLzxRSlGMqm10twfOM9xEN8ONpHCIwSwPofcOb3bwJFJo6G7/oz30DS
MR7srqM4F2nGPqnZl6laJUNRzoNggnlhUy87SKP0rW2DzrhaEeLVmO9dqTSxY6AbkFvKhhf5JlwE
WHyseXA4ozLf6Nj7L31J1knz55jYAJFPL4GGLN60mdC9gdT9aSVazVJ7Yfdb6XV16MPQacbAOQWN
VeEWQcyFltOqudsUWg7vEDqaeQXJg6aQ5ox7XhtDhZh1gO+8T1qFcGkdY9Xfg0lzk3bMshjdqFPQ
YnMTbC8lpDn7IzCIvB/JZy7jz0y3K8xuM5bIE0FmLIsMCetOB5X3fVzdNXnqJE8Q1LgmdrtvxCyv
KHldhfX+7BosX7vaNgM+8iFSJ74lKpmHkJRJmf1akiVJ5JTXt0T+4eSME+atnaAdZFaVKx1iWa6z
tfl7GykLjcoq2B4ROycAdqaWNMZI1fdRiAHuUbKsceS0L6h+9/v7CIfTZ87qcwf1Ap5MEHUbA+Kb
JAA/9eMvHbrQc+VSdLzwQHuQnfVCTorS9HZezWz6hDNABEzJLjpy9zDgBhgYyHix0z8AUiHq3MAg
2meiSr7P00gWDiUC+4ewy7Ab9P5laeFlh1iFrXG4TrMteSuHLEes+N5fUkXpuc/mRIEmcmyttg9c
7UA/urO0RgXQSguaFTtNHm2Ve0/Jg/AhnyrVDipOQMN/XdTLFnoPVwRt80zvMPJW8+GYJK9xfYrO
dGb7+3MzqG939bWrO2b+2x7gQvbtTGj0LsAvJJmzx5a3u/Y88saYHlZUfmSyNvL3xiehXklhohOd
fcS12iPIyZJmZK9Fakj3tUMKjPfqFCZk04cwNv+sNAghjp8EQLIzQAtIMqNWSP2IFUVFTDf9r+BM
UVnbTZ0YJcgIZGQz+EPntrDBfY59ExM5/iu2mL7FjuJZ+ShdLER6Pmh6pMUSN7DSULEhj6qSYSFa
clQ37M7c3WFQJFD8JpD3jFkX2tDUC17pJeBf17H2B06N2ug0mJfxRYuS5KCTKmYULz0bI7PyuUjX
oMjHipkvtX/HBqyxIGI2jZYZzWf/lILDisN9K+n3p7+YUtA3czqEEO4EurOkrF555dHc5MrGvPzV
XpiqhOx26u6VicVrpOCNTiMVN3irdCrFsmvNJChbIG3rGfw0UCsNCheERLXU66WOfwrkyU2IrrNf
xccAwclxrkw3t/ti2ciykgqMFuPjb2mgdo8pyu1z5FeB+K5lG/QpaWKAII+FNPA3SiDGdVi1CeuV
lCu9m6ZgFQY1gorB/Biu0uWy6HbHoxqkQWpBnA8yc3tGwsqD2D24BgVlLb3MwGGYTBFlt/t/5R6P
spMRe7zVDNkgAXAMxmvw/wJiXhN2sJ3rff9Fa4aF8J3pnBPYRcLqZJ/mBA/zmhHo1HnEKQgIeju8
xbpbGCmINNDTzur1y/EjBwXhevcRBo6US/1ahBgWWfjKZQXaP15fcdR/JXZqw+RsAfGlIB+eNI0A
LNkpx9IYTP7bnoV/fVXVOoGha1143exSigvV8lRMZRZ1a0igEMmQgb316iSZeMguWUqpJ1aBXmLN
zoZ4dZQAHsCmTh+V6U3XG4zejfrmFA5uBduB+5OHqcMIW1akECuEO1nfotg4P0O0BnDMBygz4Xts
FGzN3QdHTAwpMq58rwWXlqOkWRNQ9PpP1N7Tb5qWtbVeB5r20pP905otHQ+7+LxapgxHhF3NfNM5
Kf+NCgftMfYOycH2vi4IDU9jPLQKCR7yO+HEVETVs/iCTXEmAWGSgg8gLMSmKG4hvTOPY5UW86jG
3HzYUunrMn2QpcBmvO8M+xYfcHNY0J8eTzfnpkbhvaIPVdiil5LRA4qpc9mKGnAkaBpOJxfAgSt6
Y8PMeeNJ39t6lgf/68T+cgMZe6dln6UFYlm7MTWjhQhDpS1ZTm15/0AcqYliusrnED6e9SBGJY+S
XQ5Gp+XFjLSL0z1ip8vvi9gbxQqMjvX6L7DcxUcJ9nyfK9Aou7nXcuRIX4zsaSV5hUu65P+27xWK
toZCHf+Na3u5n5wNMqSRO+cxO9qtnA4CWTj29lwexKblXkjeXh/JcCJKhLhNxSAOg+SCcQ9Pshjr
1FRJlB4tRyaQtTkca9rgE/RuON2GzF/ef1Bq1hxsvsu1jdGz48nAA1KgvN7UQZbJGy0g6k8/MuWt
dtWwD30kuHMIZg5WyuyFklMjQmkp72iTrNyn+Mqr0YORMEPmcEwz37Zu9Gabw5wO/ffvxfLNbPdV
zp2+YyVTTkGg0ctOj5Q/F3YgBBN0SY/EBfUB6yq078MuAab8Fi2w4YvFjqc31+Xkc68WeS7Kv2Ae
+3kgKHK4og/RPloffheP/dtqZ87uVZP5CGG3cdWWaH430hcXVG7k1kqCmr6R7oXKFnus9+tkr7dl
mIvwAjrm7QSQLMa1ynwOij2BNh3xUATXQLAHIAOSvqbazjpgWkMlsiSBJOM9+CVfx/CaPJZZ03Ak
QP5eHaDyiJ+Xh3JTNfA4qyEWockwkg8dJP65eXydWLtJqU04uJHPqIv/68UX4w3zD7heu+DFoq2P
hzt+gsxfAZVVpKfZxpnfVdELj+RTxbVOSwytcVhxsXbnCDYI2Ge31TJ6gDZlRyu5DDra/esri8hE
4TEvEWSz6yT/MmV/pInktD1SfoAU/OdEFb0cmHqQkAnpxT4ghlTo8SV8rLNSIe+/Ka/2khET9N0P
kK+C3tRDXkNg3ocjqKTfWbw0tFjGuwfHSaO5OpsVyKoGegsh3U6zzP/TV03GUsYgfdZ1A1fwdKyZ
+6R7CvOnwOg4rCy1maQlUCWGdnKSKAd8SVLufWs/9DqvC9SJPNEDMUXFev6S3NE40lkejrPDk05/
KfvAjW3/Q/iqYeD5re1WX4uccMVquGkqOAz7df4wdwcG7e/5JVd/u4EGqnOhBTMyS6F+0v8ROw/J
Kmiescgrzha8+4EDse+DgvRuhfegX2e1LKWv9VNqESX7Ee+UgQOYj28wNRF5x2O/N9AhSJMDVNRb
2xL/MOMi3917QZ2VKJoEcoudfq8B0edtmAncodIulY7NKNx3uK1dhf1f+ByaYvNzX9AmxwffR5MZ
i2DgNjuMoZbeYHWgfA9LAD2t/V86bkkWdPYtbSfPYgn0idugNHhnjZYTTcvNOzu+bS9I9Qwl4tdj
uiEMyBL6f+HthXfWLKdkKrU04DQhH791ZImUu8zIks77wGCGAO6mYpvzUbDuUldLQNqWgiAGI58r
y+LpmvcR1LWn4D71nX+N8fAEWjr9RpNq8REm/CqG8o/jb0TfXWqgV6glQcIgLe8kXNa60MfZWtYF
OoCiw6lilpNAOt2iSCzkF5ferRmjnml1+oiGzKE+t2fju2hZqZ/u8d+l5rsa5bcr0+XBqBN/hn6Z
zPR89mNWwjp3PW7UJI64Pb7nvRYX3e5ZRpsuGknfXstlNiHBErpPn2WUZxOH8mIGn4V8B/n2up9K
6ut8LuPt/wr6Nl+vf8JSLHMBzKGL/tnSf71RexKPIN4jXr8LSNAu4L1+EgAnZNZh4EPaQeKrabgp
Dk7VdAkUTVieB35tKGL4EdsGIdTxsPViz5WCk/f89JyGBSDz5KqPDVkixFVVPXT6uWSBck6tpCzp
2l6U6E0y6kQZNUO4k58GhHk/pQAbZ3f3DA0Q4btmzBZc85d3p+Nlsc4R1T/rfBwe+vATzhDKpbnj
OXeeEAiLUw1jlQD5Pxag5de2vhW3WJu77fMKKXcYL0jVTppILQ/RcMDfpio4wKC7kC9hE0wpeSYv
lNp5ZgTgY2f8fMoWfB4+u0WKg/Hg4R6NyrF/13ICHRKik/RJd/MgJZX+EZLuYBBwVmtcUVcQxJx8
FC+6ZdTr7orldm0GFDF1Rv+3C0Q1petexkpSEczCMzO2hdY0YrHzf0Kndekaxz1RaWIElZ+mvUmk
pZ79g9K/d7nwN5Ur2O97BjbKW5EH1aqHL/Dtx6jEmN7aEhOTkQC2GFrC4ft4X6yrbS1epd9ZGAp9
hNic20+MDlXJ6AYTs1M5MWcxai+Ukm64N/rAjc+aiVDMNzi46XI2z62Yu7GUpNzcOU3kci5JjvS8
QYYHOwPraxG6ELuWOPfO6i8drG5Ku9LkFV67XWHTri0DBAhdku/6B6mYQ0PGCRrqrGMPy/wi/FK3
i5gvrLKyzrNFc46GNtslK8p/LUohe+91jc1Vd5OxKeogAixtQ4FbWWk2NJUS8orwJryEvNgNrY+z
/ZkiRzEPYky0OhHxdIIbfX/9NgnbTdWS2VZvFwm3Guu2C9+bkmhD588fTzHLsmWB6K8iNtXHpF5s
8uUIJugbt3yg276M29VKBlRrSQdEZyxPU6fplrdduKQMEHPyrhsXF+bFEEkneJ662eCvyvDN+uvD
Kiw1OTXuGhPX6Auhso1NQMqhxrCl9IGTL8vg+6WtEZLyL+eo9ey/v742gCBI/q9Bg2YdI7sUmilq
EIC5kXl4v/oCghH3G1Tc93z11suxwhB2Zkr77nTax7BLO5c4oQ3mKk4+PJCpJdd4Ka4a3lVICyHB
IZqxNxhojqKIQPyDky56UQdpJcB7YAKVB0cjgAkS1n0MLjs6oTp3rDrQbkQSq6YQq19D6PUR0mxd
CPwuCqSbrO/1v1qGR9vMhbzylJR00BVJ8z6SBs5De6YFda8L30cFMlUucE3J+7Bj4P31CTWRowqC
8/q8PkoW+eXFK7BllV+v1GpL9G3qBnmTmLuKxwFZkvA7a+yAQzzCSn8geNPJVSYf0ecYRb+RhA1h
ucWrLuW57sOI1hy3NqbnJ1FPZd71ef9FPGuSoWI03rDsnCnmXAtex8shyimGrPMqJnVWe0wdzhVL
wy2EhufFIIysosTyk9cbZFiuvHIyQNX74tH29w7PmfyK4xdi/23XSJGppO/i1HKhv61g3Kmb0ato
BK93v86S1nypeZ7YLe+8/M1jv/wv1JgZdPFuIusJfP/NaOwA+E582e/UempWjDAvdjVOcDQjxn4Q
3UUs/2ZRGTYtJX5eqJl8Dd3Rh8beVFq37dUOZmLdtudaGzShlJH0xlCKOWvDPyiK3tUpOwmYFRsE
cbPhtbbs8tgwA7P+2oCvMd6o3HapDXDw56gPLcfyU5g3SIEKBYFSzQetyAj09sYBvkB8eEd+e605
+cw77E51LL8ZB/urS1o0OErldgUsr5xKu62pL89PweXmYfChCirw+mhbrqY3CILbddNxRWpZG6WJ
5Q5sSKsc0PIU6U8aGI1VMEwapQJDSwWFTcE9DS647BPOaoVVuhEUFVyh3aYuTa6DRGK1Cj/X5Qah
p0twd6d2XzjHPBGOLEILbGH2qljn9q/F+0sjmvb0J9OjBPkZ9Iwn4HuiBM16e+zA7/bDE/GAjvi7
yKFv1HPYkiDJIEubXQ70K4m3mm5Uc1gbYZZ8KIMvj0+9Z/T3j/+IbWKBwUcpLQh6KB0hhm9MHqX7
hR30MsggI0tZaUidBT8Q3qF1bpsWUdz5+5bFXtdKsLS8gvNCC2qvR1yeF3uhrXw8kOeqSFUOgTyj
Y9RvzBhnRxzn+MWsW9IamiwOsH2KaoZ23gs0GWv9mBZlIp59po++hfTFX3ZOxHM1a7jAcpiB6BBf
mSNCpBtwAOIhlRgivlCa8Y5Gol2WOp5GdFvh6QLqKuBiDwUpStGtQ/TyrNYeDGlyggffYjhxQBoB
Z4FteYeDBrMSbdPCfdVC9dRO1boWMfZGpgNHfTz1+gceae+9t83UTRi4hh6bvoDEOh86TWvjDuSJ
P4KHSGxpfyhcRidVeyqMBHcmHdmdIk0CWqlDKzDfZLmKtFyO7mGVi6AX0BRE9Hf81ynn7Y+6PGHe
URFrROcEkAi28BA5DK+6KR3HzUf6iWou+gwLpJMMEXLjfk3UJxH6P5e2R2J5fNgwPJ+mVtBtOBg/
wP9nsTSyUZjmQGcR2e5pLoJrV9i/kALESE92IMsmsM3MDkaaevS3TnFKqT//n9MVlZNO1u+O8CFc
Sef5a/IDBXIkkEJjCPWHIcqbg+FMKoKCboHad2cCY93VePk5UHbRfpUWWlBw3b1BJbtGecTq+tT5
7ZvCKZ2P/FhSaIJUsL3pXJFYLq3jGHicWk3mndJXbr153ZxJP2X8KcwiLptbsVfx8qEJVyV3TbWd
JgzXE/LbdN4QiV7qxCxTdnv/lV1YyznQsOoXAF/fAfg869//AlvPoy1XRZQzRZsfQj88avXBSHxi
4FMP//sChh6EckAsPNLtCSgfgBkLKKTOEdoTsxg1PyPZCEJTxENwYQ0utj6Yx7T106i6gI6U1Gj/
QhrHMIQDF8wUwjiN1F/RePwTAU4F9EFwQP+r0cEiHtZ6UDI4N0U1M49ljRKfM7L/HAEn0EJoBhFA
5a1HXNJd6YE2QATD0cvDqGG+N40N2qyTH911LB/w0qAbWxFDkNb2Kry92JPRPgaXY+i2yDeglHjN
Jfni6w2N4+uLOtJpa5Th8rMtkBmZdK/Y0p7tqcwguJsnfJ5nVTsR+MV0nj1QkiZM7pS+ut87W0nF
DiJND8/xHGifwkvDJZ6cDjM1wQaDYVjazg3t9bAiKDGuD4kZyhHmI51rt+cdiTILYnqKr54ZKlmv
SXkSVoaBiP9F4tJRYm/X+vZsUc48Qxb1kjPCAQXLFwUvX2l4BlmtFBmFPSCJmlhBaRQ2C8h0sZqY
0VZXG77kGZphzxzI/X1r5Y55z81q1Hn+kLsYjh2A1eg/cOfuA3ZZGlbfb32Go9NBbLLzIQWFUPkV
e/mc1Ki5P0nbdGkbG2y66K/lIrludeVqWQiniHIT21L+7wOS3qyRFoAnN2hebM9EMAJhyajdT+pf
5dWuNDlmBciZJKUdFn4P5SsCXO730t4/lRaV7D/DrvN6YuQpkRNM7TDxBky7k6d32qEx3JLbXZBd
M4cZGByk+zOQ1MiDL9AnVw36EJ14mTAfL1juxUvtif7/nZwjxBUG2+wX+AFIKf9dpzhwjPiuE5VF
2UhqdrH0FdpR7Yl95eLT+tZiI70ticrzscPB7E+KO6uleNgeCG/oiMy3hAYDp69acCpY+YKnInWF
UbGfriKAxGjUjHeX8sh8/pcVad2BWXpfhnBj/8AHkeR8Ulqq7rWZ0k6YqGubmWl+f6PxQMSSINh8
W6UQZyNz7DsDOq2EJO3Hxg8MxRLf6AAEvsAxnAnzJ8tC4cVNbC+JwllGw+REwJbW16Q2JukZMsmX
ERiDWdGD9PTWaWITa5Opc/AJfRYu97OwW0mE7F96ajx6S1npiyOAnA2y6inh5WKgTd8Ud6ydl70U
ks61a0+1pynP6EV4fJH/CDf4m3a2HyRAUPA9A9pY96nWQ9REVRy8NQVlB9rzLaJsMxVuWLvc+QO7
L9a/qSOmPfi0zJUw2ePY8R9be+Hw7eUrlr/6Z+NJWUW0nBw7JxsfIRaMBew23XeMH28AOk0RgTD5
NcPf4to6yYMKwMFq6IOSARs021WlEhjhqxmqmsq1KTNqIzEj0SqHp57mmYh6wyFk/kNhnczz3abr
oFoJu8AspY25nLrB/VWQ5dxxRcQtbOHLsDZLltSRCMv9IymhDoUdgk22Qbo1uD3qo3AnAk3MrK87
F1KA/HDO7vV5C9vDAAV5E4EWswDW7DNqN1Fu1zJfTbrDfVHhKuLPQLqgF3UW7uDmMxy/rkY3C3XX
n46pPyOmAZDqKhTfC2M9s87MR26muzecunqqmRIWQUisfvOZwKoKIV6nTByhO11i0wpUJBIP6qW8
1ewZqv8cRwIVfGi+zWKR+oZFnJCWQY2rn0/ua3brdMzru+gNEuhpMsSwJhB1Yt0G8c+Ph9Ccw2pX
dYfkpv1PrDjnXUJ9SrvdiPIx7Uu92wVhWrEsobKgQdXUPAA+h+VpTfljq3yvdnhxjmBx8X6HgXMF
PC/Qbe0cKeD9oq5vIHeZf9syI4bHAzp22/7TB4E3zKuNdzkAGZG6+Qs2kNZToNI6UDB5/xjhQrnX
8JTppqNuYDxhsnJMgSe1crbAYjEZoDuHSc6TPYuz3Gb047k/norjTSflgNec0VGCLLyNFGsw88s7
j26/9FlZgFhpIhtgT+fn6OSIWmehin/HeKh80Y/Mqk6OEPgMol4oQ8RAGY1lqi3Bka1u6LzUNkrz
4mQK2qQaEKtCbxnoGRw55SDmobJicHCpuyxM4SwsPfiaX3oF1+Qj0xjs2INPpapla2OMEXmBJkY0
uaOhxZmOsOtTmSwmthLKnggAGfkUL2QHgn7Q5pppim7QcnnFv8DFr/wF57bxhJ5M6CygD/i5mlA9
TiFm/2AC+BfBRNPv4KrV7VamWgCIRSeNJsltiTHOl8U+vKxsGlOK+lCbNIrPIgSVe9e3DzPF9JQX
NqiqMV5UZ1pX1Mlbu+FAs/TGwQJ/n38+BLts/IfQ26ImUtRgKWWtcE+z8cHxIX4I1XfxxoxexPfo
1Zl0GFgdpV3pMYga1zIf4eLTyp39R7y6yH2wP0NzGH30vqCVjW0NiFT9CI03EUv23uQnk79now+p
lbR3r7M48oRrMQ/syuHy+OPxUqwOnYrqJey3+oZxmYiPXdEOFuHcGJlqLRinEH4NvwGjvQdC49Kx
j449rf/yFE3ZjXbHc60G61k9i+iqcad7oLZcKEtyd3agfN6OrDGN/prRMW9+iUobWTuYrKz5wrRd
w+OVDHPM+0XMWAMNyqzUMU4nCQ8liZGdSFDOoNvWI4Nm4c9kbFDu/sFsQri5P751uhVXglm7C/wU
YpZf9fKkBfQOV7AeOIyuczs4oeG+24rYE5kXx+TDs8UZ6RPITcUMSnJPPnGespA13XO11S0T3fQY
540/j+2CtMo0R+ufVb2ifCMPZ9mckmLUQ6Iy3VCkBZFx4zARSwEs9Kv6+YyVU/dztFPCOrg0Ubav
NKv9/xGMne4KjtSPeEX05c+VfOdiJb84CLu1dW3Npn7FZd71pVLUKuHnYdKwYa/vycB423R0AXMz
iAG8AD12o71GhLEw4w7N/5oXvj4yQj0DnDowXuhRzdktAOzhN4lDPKVSWVcmhYvmqMXBgNwrfxZb
WRpverHD1XR03cLXt6+Ox3IYEKoMh6jYV1zKSzVqBlUoZZSAugCNcyQlyXA1R8Tew9TJw/jPzF0H
nVMztrhWlP8d/pywIGieYBkSk0ik9tPF6KQsFnyhAIEwrX8FXaQPkTKukzjFG50pZzbO72hKb0sI
Ohi0hCZ7ZBSgQJ/Jp+KVV/9LUF21makhnkYBfS9Q3iMh3lZvp2UEBSfev5nrKk7C3EOqJdkvLWyf
0fNXA9hrM+gS/nPWnL62YLLrSkfK5Pz8E1YS7IBaW7X9hf8pqUonBt08kEr5XsfxbPWSaK5YSkgX
Ja1tVvRLiIATjasyb5kVZCaI4YtjTRSC3kaSsGE6CferOBC+qaeFxcz2+i36atpGR/jHBPB7axeg
8W7ssWXikA3uYR8JWPgIzHOSm3ZbrPfSO6ji937qcFsoNa8OzAPt0Q2ezMSBxAk3pbz6y7OH/+J8
+wzkfohJl84/yGXrt/oK4xRp4g+w9a4hkQr0r/fikUawCDXNW01DHcZnGOQtTHw1KPXmmUpXFu1m
KKRbp340Bk653ZDNBL7+n9xSNibh2lTwFd+SyE/WrX4ul+QIOJjyiOCz/zXbI9hMAyd6M/o1iZY+
Vrp8j+Hf+CDCbTsGDHi5B/AqRG3gH9aEpk5GRWQvg5l5TM+j9xrFkF9wDjWALl94jP4SobqOT/O5
gjlaExKhQmLLX2R7qoNjBbMRLHuLrYiyAk4t+KwcrcduVM0Q2glbZq5rBu1Vs1R3IWI98DmDIfYy
4B3cjsyd4/9lUODEoVX3bEKsFkUzIVWkGVKasywN407xcS0JzY5SoXud11PDjdGbTNptMIq45OFf
0kxl269VMR7oKknCl+kIdbYz25ZmwGdgqYNg8bw9ahVP23V9ie6rZ4DgtQRMES6bPhB+iTAhtdDk
rdd2GNBjq4XK9vj/vcavdxNL6Y/tgU6kDlcKJTje13sULTvd9Lkh/3FNVYmrBybGOFzJjjg1qT/x
/FXyR1NvQfSGLxPQqDRMY7B/d2TVwnK7dZ2xty/avdqXYV+Lx8cBDCHt4JCMPcmhcgjo0EScwDoO
7Fst9r7t3d9sJTtwo7AbpffI1vmHXvhgG4I9qYtLH3mUT7Z3mvUPZz67pdkQaAS3GAit0mEm6U8g
P9bJ3cRmLAhmlgtaHc4nnKaQyhhh+p66F5Gvw/UlNDr1IAISIZn9pO/OhzHGCT8nRn0GfSq6pEBP
MhnyNJyf2KoQrd1lNH2rm9JaCZEPhiVJWnJghCeZjEcXi5A6wvqxsYjfbSvisTIzV1+RliwDUoh6
4kESdVb/n722su7lNfGOHapiu7h7CQCx8sH5QS33Pnt8tpiftK2YPWxv/zYvCTIQKtMmcFGvj7TX
BWk7BasEgvvQnojYlyP2hyDjggpwhzZEFc2Hk2BlhOh8fq6WIw74oKXplLHwONe+zCz5EZnUamms
nJzDjavGF69kGQ2yDyT41W3XqOIIRxqJ5Q1eGdhAe18FWMWviLjrDr0ZRmyMLR6sjldRt/N0eqqW
IRvpTpv53ylcpWIeUsuU/CqVk7uBQTMRug6zGO4DKkyG+A/+p0CDKm9BcB5GxXLKTZLWISud8TOJ
zHcvtQZHwZf9WnJwteGRzVJzv3ajq4AR0EPu2OxvdXCutkr64QKRI03uAFnsVepPQsgtaBYeFHrs
Ff6ITT3cjX5alVPgcG1DGZ7niMxNNe0XMQFGETNcJs9S8xBgjd6QAi2OVSNiI27ula9wjSEkMzZ9
+DXDFH42HQuLVFcqf8bLja5UKv4C+w86QW0+SSAIoVFDL00n8NQoSZMFXUTLhdmehLCcDjixxQu0
ZobbnVz0fuhKcdMcvWX0bth30hzhd0rthmVvx1Sq5MMyYijo7xA3/BdK9h/kHTxd4IaqTRK6gdMX
sESSHA2+8uv/R5E6ChPcL1Wkq947OJYuQWo5BFUl7AJFdvt4wpKZyTNKVqKAcL/w1s6OhohdTQ4C
sPE9KT2IqQgD5Ck5IM4eDQlWznYwg4+Y2zGKLz8UNL/Ll1Adws0fsyH0c0HGz7SVYd5mS1S0I1Ub
8OvhTgJrutcD7lI8u8pQWmPTwwe8lagujg0ZU1ybLYlsb7X0oSwcTgfPLnYkXJ/S3N0dy8UwEBuQ
X+sKi+z/lMSPO9GX1M9W8xZxD3I7WfgJ2X1fOzzZMdoZb/qL20nidCtjquiutZAkAyD0na+bfEIz
4Zu6vfN+SlxKhqImJ4HXkYKtIqB4uPqH0F5EclBTn2OIdg4C361HjJnNKjKURTmNBHBW2xRfFbrz
6sxNkfLdcPG0rUQIY7nVgieCvqUzxsNXrXB91vh/VHshojHpeh1JMdZJpxUrb35DtSKafW04cl3g
rVdZl9bVUw7J0WdvqQRB/ohhgbxxCPIg2x/nRs4ItpgU8F0QfimRs7PzhZPeJ27zHbau4w14o/Ca
Or4b8cdrV4MeYk9yvi+eP/m/pIb0Ealnka5+0fEPohu0yZNFFpgd6tHHU9XCT7MVKPkteah+tlLx
wylnV5Af5zkRm49ezI1+TsibAZhDx4RV82PLziFJf3fnLMShUOwn/t2AfNOvvM33qFlhc9ix7iU1
+nuH4sRn2xwNhQq60BejC4i6NmotLoTfMGn0Scr7hSeg1CH3hGdtM1fbAM4eKsP2rCRd9sBPMO/i
JuYpIOKQlKEA4aAIntGo4pYtfHaJuBBtUCJjwFQNrQ2aQ7VUKnOYLGSQR33tX8feIwvlMkCBi20+
HdjJ1wAgmBgMa3jepgQ6EYdXxJYBEQIu+eHVZK3r5hq1kl4xAgZW2dd1rUqtFfyYIJZGCDEjZmXF
k1ao3jKco1pvTvy93q+5SfPSONAAzy+QTJMgl89KG88pz65YnF36OX6n4MYb5v9bqzjF/uUp3EDF
BdKvwo26YIBE6kQfoWfvMMRSfW91BWXJSqUFJTE20Clml+F9QZRrFtK157057MK+6tbHTehSJKtx
v/WilsCHLNlPs0vtplaiAnlTbHOVvIyRoOTZMR98/YMTM+T/CHxqGWx1sKJTylkOoANRmSC2xZUP
CI+7w9uaym8cIYfD2TLEyb+XDLZ3Bqdprtxoz9VrUJuAfDPH3LrzAHEmExyz8VK3sCU5jozMoug1
lSR06lJeLmoaVavZ5kB1kWGi2d0vUibzNfz/sPkW2BhERyg7uFbHYZdAbvWlmZlikuNK+YdS9u8s
HbEYheyqs3SEO0Pd5IlrUovndf5XNtkmmO66iIsaB/kVoEgXe7wwdXbgYY+F/vMJksnQMLtTOdtz
no52NDVAhKPWb4i61F4v8gZD8H90nUj2Ynl7Klc5F2awRuOeJ0VTqNdSIrssL6WzWbaNkQmjk9Dj
9PSDBNOR3FlEL1r6Y8nzfNg6bdJB4d5aVk0DIbmoFkM0wQhgW3eCtIkgNeTvZ/XBnFKLXfz6uRTS
JHYcdBcF1PJOecXyEvYR/ExdlekFsESGIt4expeK5Uf3lEqs1mfC1WeA4EfWXpG5NEsG3lLaHsJM
YR1BSgPKjQgwMMHPTJcusyrTNLoAe6gixt1OQ16mRkyvr6pIndI6Gy4tnhyFgtb8NWNIpme7Vx0T
g5S8a+aDRBJnTrZg37ftIpwcNMIrspLMCqkrLHS8jE8MBEB0cGLdit8sxGgyzP0NHePirAyp3w4v
UFRNbBTk/7xRUa44IVegyosBmESv+6ON5tXAv8sGHbuZlMOEuJqyYT3BQERDQ+M46yRcaE+2sp2k
zvLfPjEt2sd/cmxkJ2wmwWADQKvFIPMWkC0Ky1WSPCtSOmKXAI0HXTiNh0vceX4shxF+2icMuTiJ
nu7htFdAEitzrOp1/3ecut31PEcabo70gvs/DhHA0MaTW8TubRZJlbYybOQLw0SZrvwut0rZNeZq
DUS9tB72MB8jXeyYp3bpMqtaOrJ4blTzWhaMUHWRP8ghAcayDVP+BXjt7IyuNLGHEPfe5lRs/wFh
r2vmjSeh2C+H/EBE19zT2C/5xL06hJSkm6saztgb3woFk2fAU2SrA9W7wkW5Xh/0cwdV9rBNeZLg
t8YXZFGGCag3hhJtZOcqRU2AwiteN197VzNhv98OdJEGMvm+QXD0Stjv1GlUtbubXR3jAa3H1qFT
pR0Guiv+GMHvQuXFBSl6vgg15Tc1TV0RvmgUFzzaX0H9ikdrqzU4TTjwsWeiSXIJSXFGvLH3BOLC
OadTXebKCCSEsVNq1Lv679QVVM71hnRLJyzLLAzPMZcdd0+keAyUap7KZeswkIGzYcMIcHETf1nm
4KqNG7C71VkmBCbKRMnMbFFBrVh6CshtDuYZS/WHkz5MxXzdiHa6Rmc3U/BdU2xCqzh6PF3TD1ia
CiUFylnKpUcXLHSl/DnLoIsdqPdMuANx99XFubNqELaR25LE9uhT0QcQKOdt4nE3TUKDOSYz9+YQ
SxHZcda1fKW8acY6iLAubmMKzQ4oZp9RMOiV+1inutbW+iG6vwVolF3qCPhwVhntO6dcSJ/pIFrZ
7CNybcBe0+jQ4AOw/+M1Sban/9pVY7fD9FQpyx0d5f8nCP6vpT7P/6dtP1amNIQmH7iiqiXaIav/
wCcOzaZzhFybix+yGLEucLK7A2fEemmJxyWoaJgUYmffzttUwLjmexi/ZYHthXZ6TGb1ZmMrF2H9
hfubBwCCC/C46sICSM0VhbwrOYXA4aB2tDSR3QE3ZSpuMZgRd02dTI6Swwwa5pM59YF05gW9iHVT
yTvxINcPV8NyBGl0upoCurZsUZRd3uPrKpJ1Vu4T4uUMMkmtqztULVQhAnfcV0SFlOOA+UbEyn6K
UFsHJu7oAIiTkSmWf8AQt+4Xl+STDaD7CFXuJdk6cooJ2Mek91jJk7bsdcWJO2uByfsgPwyyzAbi
M1fWYZ0pRKzvovY5KRQh+o8UsyDhd/9nVBIgDbZacurrhVyWouzDJHaKo7DYCaJrspYUXZ1qX+Hb
fKnzL/p9M/x2hjCc3buwKqm4voT2KRyldMaHaZUV4ZZuC+gBVGACjI2a1Jix0pkIuaYJ9MtgWMCb
0wgatIfNj1e5BNZN6zW/3DDv+WVKXZloPUqJy3HUU2xdwfId/WXMc80caj8fEMIh4X4h+v+MzoZM
uo0mUNp3uVvo5VPs1RhIpNSvlcz/YUmO1eKr3WtBIDjFH/rhnn3labdFIXlXqdJAX7b673GN7j7s
1f9mV7DU6ZjhjR2M6TNjWByQjSyWUNNgkQvmSUZDpCO50MBulqOO3Na4RIHD9cdN8YC0HHYb5Cbb
5t7WdmVcDfxget/Bh2DiWg8x0nxcS3XNGIPP5vZFQNe+nRI/lmZLBfvicDszFGCB+X9hApiQ/gmV
33npM4XSY5NfVI+rqq2YU1n3uj6AmCMuFViXw2wRGnvt8BLMIJQbmsUHarbVwJkmY2Hj4DD9xZ5C
/JiUzL69h+CWzP4z5kclqmyMarz3A3RBbff3aYN/yUk7o+3hOsViEnt2lGLlqS8lE18fTTlSvbqo
Cbj6n8I/jNsOCY9z58Ygw/p3LDLKHMOqqkzJ59zzGQ4yo2JzFfLQoxNTgggsE2bxrBAWPDN5D34h
fXEQGKr0tJrpAK6AaF9xCjLJ4IDvxOhgVpsltJgBWIq9Zjy8EbIXWsKRSWCSl73AaJAYDJDZndPP
t9Bjsw8KiDtL2n/9+uuzjcAQhRHGU4MnE6gjkHbarSwEE0BkD9AvOWKKU60lfEN/gnf2lTjw8S++
nWam5CXSfta7g9cPbbaa6/wa0fCaiRXLJcDjfsE6edbTIV1kxddQ5y2CgcvfkGAyn0ACc3H00WA3
8hZGQkalGOP/Jz0euaJuMnHZ8Ta6xuPjCk5rFpCLY9rWnFblQlmbWEl0x6sImwgraWowwmFAhZYm
tMx9S/jVAJ9tEp19axJjb4AhmFZ9rz0DfFath9lIrQP0mV0S62aKv/FcMH0cjPYbbOKWuSMnrpAw
/95AQileszapZy1HTF2W8qNMGu8Ad5GLpZ/noh+PEaDendRvkDVRPf4UUukphjbS2eetqSVIJTA/
jILOkrwKBSbjhVaQ2bdDqpn4gWesBxNhwfdsv7HwY2lHgqkZRAaja+y9rcT+4MW8iPnij+3b5XOl
HfVLeGxja+i07BMFWWPjolnjRuK2iwtUhipZqy5PEf+I1bCp8YT3GDScJimCmqOHhM/sgbtEKG22
m52apN6MT8inaX1hT+cPUmI1aj0R6Ed55KiqronoMTZloTcznBAKiuG0/a+p5f05RhwDr8CjR0rk
zrUZpJzNg3lqhsISpAXukab8CIYCHauaJWwyLsedhdHtYVXp1phtI5W10z9rYh4USh3rLd56Ngqx
fiLT0PT8mTtwt1YUcDbTWQPN2DzXk7V+Xe/kVg1dI1bZo0UkhX9NfXrVOTegLcBhvwAqsRnPxwc5
TiWFNcn57CYn0q7jG/r4CxaZFneeQiK1aL9T2H3CHdD3PGMsoh+W7mnJbmxmquoVAkNvdDAYAAr3
wxeCpOzatyKB3jAieC1JfQg197rQeHVfuYkM1+/a5fEmobINshrwFzvN1TEiCIraZV0YDKpEAYXz
H9wphJxaApVI0SUew+ZZ8ayub1BbSFAd0tvYRwJbefZfbpvXi9E8pcBsVJQH8vz0FX/dRMF3Lk3x
jWJwVwHie2EhMBdEB9Q+IXkP4oWQx4rURYkvnprOdIvRBxzwaQPFoV9lFiZBR8pQOCMHVrUUi9bM
WxcXhGZTAZemz2Ugk3dF7bpWNLEzEn9wMFHgW8QxpkRi5u/qBRJi01Q9lEwRkZnjKV/wj6wVLHPm
etfotR/ZFNczlo5DBmalvbXJTbIwcr3KfWk3ScYmstn7hgrN3Frl1Nnlf9u9Gr2HYVA3aetWP05I
GnVGKFzN4ZFB/MHnQoli36l2kW2cW/Zra8WyXhZsQ4d3UWaD9SWBavBTD5B+lB8OH2Ns9PB+dDHj
MXU0PAC7+mJI5fpyCWe64PjR0BquiSg+/fg6wgUZzTe+EPx135WDObRQTQ6l5Z+04uuzE8jCr6ja
pQLNia/OU63Vu+hSXuhNizJ30PRgK5sj5fjR8avIiuM+Pv11NVdVxKPLRKv69mfNSH25WAhK4KRr
bk4uHYVxQEOe0YWnu+XkMpctkOedY8eAGPCpOum1WDvGe35fbd8mPQSS3+qZv1aqLrMxzGh5bMiG
NU76I50dpcWi7dScdlVjWRmUN9bkcNnmR7S2DNHUc8xIs06OS/kfw190+49ebKWdOZ4gDocDdNLs
KDUj8F0elttBmsFx6vTVsd9pVMKqqmxTS1r/V26fB47iX6h/BfFlzy57QyTOQc7KUl/5DUIfTxjd
QvYIL4eTspBHD4d1R4p183if7YMKdXB59+MjaroO5mJgH09FIS52+MhhCT2UpTtr8A2N1yMOPEz9
BIe1nVCk4sZKF+FHrm4oibI1ph/i34km8t3BcumLaQf5ENU07htNzgsgphI+bagcBKGLyqapmkrv
1wzNW3h4AwOKIISEArK2y3FBPqRl1jUjKlRqMgkshn3H6IQWl+pOIEJTBPAjHvlrMlXIOxBY2gXn
lCz08rST4zZkooJXG8UEL/bOX9acpwq3nSVX/CrhO53a7ZrT8qjQWNcp5j2XVL/4dgOKf3VeglbH
awI3lJl5a8XwUWmRSV2l4Lro8JvwzkHXaYYS55A2sESiIbR7Nnm9lIzv7IFSLUR/BvpGTjYtJg14
pqm75mkdTQvLQvS+g/hV+iVdLtJZnPKld+XNbjISvU7nFyYX7ev8R8CTHEGrc2UuOi8wonj7uKfL
b5IujBLbhlBkEYQ02bO8cqi+zbH+M3qtnEBrH0toVQO3xMQ9oUNvHQWKE1WDJvAZ/3qjWWlnuPXr
xA51xNWpy6MbqRfM8CXIVht2HnTISfuqheU75QCZ7RTOGT1cEatR6U+2Y6POJ8AzSvoJABmqgkWu
vgFWPqUDaqVsjSLR7HKZstJRSC/GtyjecBf5K2htN/GERzVKCCntdTr4jmyBhTSvGJNlfWHcGxwM
k0UWrFjrsV5GyIgGL0JBoUd30hYRqH21U73SeiEDnsQvomxZmtiLg5GkQWMHDEz6OFTV2YRdtZwe
Qf4J96/EZ6GZDUQ/CxDTxTuVoFsi+fOuCWtHT9MgyzSwh7hkK0vo0PNIe8X2463qW5/8IlrSyjBX
O/K95UaEKA4RglUw2vWZG5/eqMeRcMek+YRUcDLA597nfnJkS1XQq1OA116HVzXQMW6AqCSwxPWX
3uN7gsTHjNTyOlGHt6Io6q38tn/Q/I+C/lClGCKqvcXZQjmWs5+/94AefEdWARFxDNoayUzN/UGW
Z4cUaWno98leUwGQN2LtxTKek3ajMiXljku/VYzKnTGFao31QRyKb0fvBDsWTiYd0OU7znMPaasI
yf5AnBXTZQ8nl8OP6OA8ADKA8Tr9w2FvGBC+L3u+CCoN+YJIc9JnrYNppuvjC9UpvqflIRu9s3eI
6ySI92oCh0uPL6WOi27ZpdOD7SqjzeGdo8hy3Ter+2fdn9a2G00Fh5an2JKRRKVGdBG4H7/FqySc
+slZvSZSwETx+JZbc5MbUEx7UX9Y43y+qNFFZwXv5heSBWbxGhnAwjOx5Te+fcll+1h/t+/n1HZ4
TALCrGGL8Cr+Xz2hn81MBUoilYE4/gr6PZcv9R1ywss6d48CaaD3rDPxMPVicVYT5okWhrzQ26b1
Z1y+Nm48cruMKN9xTJI0OepqGjsrWzUdHmgIzHfW4rQ5Ew6omeSVUBQXYUnfUEsu9HUYDSAm5E4m
gvAQt8FoTUbAZAWyQtelE5CacWWlkdSZrTSOprs79oNpsGK7ChWBqLfrP7bXOCMN5OBFKyfxOYcY
kKcgIa0VVJsXVXE6Sb1l4bOxSXcykChNywAnp5UX506sCUXYYovk9bfuV/U3YW3DjoGYv0SVmQft
CzECGOdxF03e0TvPE2M+ya1rBA0wZQy6nzCPvhH0mRu/hY/pKh9lwT0olE2yFBI56SG8llwYqwYw
BOqg9STWmOhimBtRms30EEj8TyUzPG/ou90e0GVFmgfntbh170bcoHXxy0usvo4Pt1G1AbXfwxfX
6NzCNEpumjKZLOe3urwy9mwkbb6BnzbOtvmVAN84qw6HOr5Ebm9Ju2SArA9SwLGGEzfvmdzbsi9h
CfsajXL/ZrbRVMjxUNU1vbTaOzctD06FCn2cGggL6P61wI7DvRUS4bRdYRmM7XYhH+VsofpOqyij
HWLRgRxCa7dcvWjMnJvK5/kI5SuzknlJQsXwkBolY1PU79qE7yiwnfBHjWVJJWY1bMSXfM0C1sO3
LL3/uRFmC/iOZf89M7NVQLnsgZGX+CW/4n5BVnUarkcV4kowevke4KQzgR0OeIVgbTmbDJPqMz+D
Zz8jTJ+smjna2oXNHIOpMho2OIP4C0Tk3YDaAAS1Ye2EqFiRecKTDr2/D52u89klLG2c7LihIfwE
QmkdsA3W1ML7zQXs1QOoUAWOVkV7gfgAzFf9aIArjZ5mhKmk0v0Ee5z4q8aXJNLMel9UmDzSPmPs
k7m8ABnpfTXgWK0O9Z+fWii06LjUDtx83K8RBwYuYWkIgiNnacPPKZc+AIHvTl31w7jrZjWFTmTE
bPkRp4OPnwJyvTL5UtJd/bKUIYBDgtO4ccjp/XHDJ+qYPbLTAMNp7SOVaXpEgD689QLRR2jopg9J
0S1t55xfHysIOa55PRcLHwwTLelFHXbSQ3sR2FZXvw4IE1kgz6WZ8emQ3n1+++DrKFn46TTXtPiZ
nzs2QDmoSVg5jAgcRBYSnZ22CF7aJ6HlusbzZQ9yP7a/eP73u2HLDeHwN6NhKx9QqgBwnij1zRuq
sB9mcDeRi30quX/YJ31oSXRlq/naacE3y+D6PomKF3HiPu9Zl28ftX05lNAt0xMiT4phwjwfqxKf
sqPNS/+bKwFjQ6XckRQYO/FCCIujpf1jGuEpeg6UVHNvlmOjpfzk5JJykrzIigqTo/fFL8TrWkzd
r9v9AmYUFtVLNTO75mxlUuGtWzZyoh3EfGJ0S6/nnFd9ITZcJdel2NJEmhnqJxt98OrE+1ZPSZHE
8ICHtFIYU5fHIeeqQz8zSFVh0pXLQJvWmy0sBs2r06aHxhTv5+ms3ZsAf5DY1TbJ5na5FBy4Ovks
0WVvJactz26/nPPvCm9e7fhYWcrqRfVaRf0ZENQoPIyJfErl8W4FF3daeKcNcBmzfhwr0j2NI4Cl
ZCyOt6DD9AzsOVbVKK5t29SRpgeZ/vnQVEUGWWQpC3yoEy4OGYsV/yaA1pTU0gKRY9GdbHe1t5dI
XyMFMDFiwkvDNQQxHKXguKCAHQggT8S1cHGRlqy9UbQ9zCWkRmD/tKPO3UXJlX5xk3BMe37udnPX
zqNDCPo1bTXvVTYZep0rubj+YQb4gD2OOdyUzBQ/K86ipd3pBi97SxdqhGinmGXCaCovd6lKKIQv
T0hpChuFgnmbf7IJ8A2Vb8W+ESxxnb7+waFg2SuEikSzFNLPT0clFNLVnhZVuTgrYk2iJ63pEQbQ
9bhxfEtBMVrMwfj0JLpke/iCSjJccwzGK4kdXYsagl9Lb0/5CGr5KgEhEEQ7pg5FThGMlfsleUHQ
YljBxXAUD8ufp/yd2tVkQHYz5U4Bue5TkUzCvOZQezjzELx0WxxAITr/VfbY8vdLHKLfuLtOHUpi
qDPyQBi4hg9qZufeSKvx3kT/YZKxCQzgVDLkp889qkbUaF+u5fudbucQWVZxjKUehV9GEIVHoeeq
VKq0Yib8gxemUdAmRuxbMco2KK3sXlQn0n1QsTQXdrmaE6BifVYqDZxVdnxi/nq62pdcbuwbK1pq
GBgfdU0cjfkZIxn/XdLXzuZ264hn6tiZDP9Nhj5Sufr3zxPj4Xw7ZCRgERmPfwDntkmxg7DKEo22
8SXrTyYNzdGI/QZAEdnl5KEDIq97Q1hqG+T1C/egg6X4MeAuKZPJyrjiNEN9HSCe9P8e3tX0dZA+
2+hhnrQJQSNK1uiXYUQmCY0Mem6WJaVh3Yp0zsdQHT9PEKFPOXKWp+Fn6hjjWuFNaFJckNNVxL0e
HPSZAlRTNRjXyrH78bq3oEeKIGQS5yQk7CxfxcWvZIyEuj+LAXdBr/B1dFPOEya59C2EfJSk2fDh
tt/xPbu40g908LbxeBnWStdLxSLTKRRt1xTQPZIj03FsxU+mA0xQEHq9R8D+vupK7jzU1Gw0fxXo
pSRmMiiniDFrZr2rSTyoIDVTc5DgKHojB2MG+NomUmmzJXqSGHSb7ZNAMCE+pBbcZRnh5sFLuQgO
4Nqc63CyeYeOOWS1gyV+EgNsvFIhVTwrXDufjr2UKDIM230/i5mJfyUHJ2KBy96vb9zHWFK8DRH7
IwooZkGMd6LImyEhZczXJnSoOLjYfMLEPZVUCnEBGGc5afWtkXOJgpCHQfZehW2oSP7JenGEv+LV
jMPOwx0EnxNx+K4V4r6174TPPhs1JR8ZmJLANMfXS8G3tSQWYh4bY/KTEcpYqVyMjIZtwsOzsHC8
KOp5p1gIqvgbLDRY0OEY8e5f/vNHze64LE4BCxuY3YWkYfzDTGKbhCluPiG8kHXTKdEUHqvf6AR6
Xcwnt9Me8PQ8NIw2mdnbsQi+/zhFghpiT5HNlY67VNG318dJOHmetrYNXpXYSqx2bfcsoZseLh6j
2mkWksk1BRnSJUrWGFBChp0oStQY9xTBzK7fK8VSz5crt6jxfssSrBh7vurQUeZ+gP4To1/Tv5Ff
k21CvIpsHFKt8yjF9J+f/2yslNFw0gbOsfv9anDhAWK35P+BZ/izaWG9P0MZRoGcXX4v4E+jYt0V
bDR0lczmGT1XloyoKASWRUMYj2LNknwB6vXfSxr1fWEmqtuyUbLgQygnxgm3CvZVPUUSAhVJlxbN
Di7Mhw3XiJjj24zjrQtOxbBhJWzDM0mwTk8QZujBfEOeoT1gIPgyW9IYAk+p/WgZRuk9InERr2kM
68qjk7Zz2qL9w6UaQt+hVVO1TlqdQL1WBxy+uz+bOcUCGtlS7X0DZmQFBCqCtmBunxsFTqJpunSY
LB2FJ9VH0V/yY1IbYzN8OMN/HwcvP8cXcs40fuIws606akblyFQDpX1kdZzVqZ6nmKVNcBlUs0eW
Gv8znnEGP6htFXJm2ZM1n86PrRdrk3dmpTe0hyzkoYiQn5RDbPPg7rtvqoCL23eTfIooCUqZucYJ
nuLTeUQZz9KxhEfQamDx89ZkUN/iMHU8Qufh2KSWmSIP6XsH3kx5owJ0dk1Hcow7IVIarOvM/LAf
MBRZqVku8InS3X/kwQw52wvhm/NXT8F9Fe0/0qLI9QmzsoGG14eHTGLz9vbFeJnJjXTMsvZuGgqG
2lLZI3tVTeRJK4Tuc9oDm64bp1yQQzZwj1gTNLLtrGpMrUMepAnnNoH2rKkxf8BINojJtRjRfUyN
Qbj/OUkKDEgHRlusDfLZKfMfzfPNiPUbq4CEeRdAklChYtmGrjgOJa4gR9R1+23vWzzUSccSipuJ
kDG2S7lQ86PjY0BPLqcXNcn5D5cvEtaaQYw2CRP9sSEke6iH89OSqYdWCSQNgQMpAEOewpVoDdyT
GogSi/7E+VSNrop/NWc5FuteYccjDLd0w1nNTdss/wQNzR0K7hqbYRf7q7zV6gEY5TGdhei6QWtU
M6xmAyxMjBK0XMVeFSRv02BpnkcYYtFJOxMN4v4d5DBr8miXJ+Fmhe6wtlZzggEPJKru/mvs48Nj
eaVxaVqqjONAvLm1YFHVqqQpFrvT2eiGEA1V9DWmO6I3D2BDgLNp/h80md9SdIL/awBoiOftGl4/
XBzba0OrfW0zbSPB0QJZkyB7In22OZa1XuLjvV+3jUUiHnYWl0BeFOANrP5ex7xOzkCVwYjkb7JH
T/0Mz78RDpnCu7ke/46Sn8SCpYq/kOInyEuE2KlEY6wsLteFjuQqI4NDTSnG71MrMOs904eXKK+s
RY3KQdfrHrQGkKniRn7N8/UAQGLDMCJjMGzlEhdcvMpSNeOo51Qt7hev+EWQr6duZE23goclFDbV
J2YbRKlNKVFcqHxG9o8JO+JbWsculUCky/+u4esXzWzO+lwqOZqM8qC35w7VS3OnKJ/kmAivtHM9
yn9IggPRvnz+4rEF/q+BONeP1PT9D3MwBuawEA5kBpEmU+IQRo01687/eBNdoJMWaAKTxN8Cow2D
k3q4qFCbu0lZi4qa5sthknfQUzUjYAmsRoPk7EwDG7Z+a4NbBoZxsnBH3C9zYVxU1ZWcppjHxuvT
G8QiPEOU0vK9RBAdjHpxnuGDrvLzTMPf3hhOWnGGwnCR2LTz+UOv872RTuIZ4PLvF725GnOguTWs
MdpVL6pUJAusP12EuWydFKU9K9PhnzQPtuhbjKHkAuDMxEg+BM2rjngIDo8phz36mhJ+N6a22FXE
L+tS29Qc9XG86L/MzU0TcGjoGlgUxa5fRYAzEKHHicWsREm0F/TTUxqyelG7x5pcs4N/J9Qgva7/
3TsspoV2HVRvIzo3k5Hio6+hP8fz8TyXG0tWMTkoLvMqBlbKbp4N1EGhoQQe/mYQSdWHdTrB8ERl
Y5cGhAEtQEKAAZ+WTbacBwEkQcueODas0uQVw6bQPRBzbv2OgcRnkdekxXrRQAJzcPGwb5dXpQnv
C5KFnRhskk9STPVkDMU0sJBXkvKaKABaS3yjhlrncChuOIKT4DSXsJF+X4FPTzsYGryLStJxZZi/
rK8O4s9AMW9qnAlIVZsfPoyLbrJGg82OyTCoMdOZP1ZpQfAxqjggsS1dCxQ70iCtRdm08w/Igj16
k8bjs9fMyDtkxFNiPjEyScnX6Zp8TEil1i6ku/ona95R7vidH8Y7L1/mX++Z6tOw7IJgE72kLkpH
P7YqgrblJl4n5qB+zfA/tlPnt3oTUuGiCUda+eaoFHYOtVg12zaKYS/7YQ3UIa/CmqB9/ado0QG9
3r1LJl1FdmoicaWgfGN0N0q5W0aGse6z0JpE4yNVLFNwbaIsEALbo0ZbHxgo6+ot6+avOKna1UpM
VKdOX3ufZ6R9xfBloPLzGkIF30iq9ERz+WK5OS7FzX757ueyM6JCsNt+oEh+3cxaBTCIa7qbeGrK
H8UQ7IVa1sUgyllUMOeLR+Kplk5KvlMqI0vYf9Sle16MTEZ2gObdYJ6JKqZY5ZI9aVG6pwuun6sA
ZoX6ixuHzCX8GJMDRfn73oPVNBGfX9WlvvNEeB7KlndFISGrFiR0NQ8o4vYp7OfLzSIGdgwdQZMs
Fad2HmyGmisz1iGqRtP9XboVG/E1Aq4FoFK2gZhql7BfybPNXcY1kYrjoeEghX61iqvNGBMnSuFK
ex8I9Y8CZ/JR2srnLNphBOADqOlzqCSKKp+V3JVMbXJoexQLwHmuf64PyEHQwPt2s8gE6e0RIsu4
PhttDC6FJKpaVpIQUT1ow3Doe83laHeYRs0KiPUQT0ueKByRLWa+DZS8QAorEdmUzy4soLGeHSDE
HepdKFzo+o5RvM7rec6vJOEbWhs0rpvraeZpSpfufYxeBfZAXGszpXLkK9c8OKHVWbMQYxDpKRBv
C8xUSLbWTIhVzJJc5Wl4LNIMNNNFuHEL1B8TYSuawMueu+tqtPQzzH0tlYHagKAI80x1TfVX4a+5
SOsECDk70xed9/Y43fYGNAQuGBPEQZW94DyopJs0o03fJ65ta7jX6sO7F1oMDn8FTxc5KjcjuqSX
ycWNuCYsyGCYMZqqqaOLgDmTma3DUo2i9Rv5Af+bzCJbHOtvX7G5g2ixGxoOeqIxuzRp/FSqsEZ9
/cMvy0AUtAvzexpTtbGzbyJWos8bj38kI9EA5I6TdBPhIdKgdmIhWjGxkctWkitweh9vPWNPr7zb
UVCnhhK8QIfcLIH9Owcn1O4j1OSMj+kO9Ngyioo49/63AyrYdOdcCidDDZwWKFBCiW0hqmyODNzo
mg9P30gbr+xa+4Q4w95AJlb+6SHG5EAYsz5hJU5ebyqYwSfltzmCrTNOuN8Lgbu1y0GeNKaFau5E
L3LX984Hkv3itr+RXNYIPRCgSHtvXqZ7RuhhcCXhXTRZ9/aUXuv66SR8FJ0G90nCZiJI3b9yXKOC
X/GBVz0ZLQ/51nAGQk5AmQ9k2tevak7+KXgegxWx/VdzyTywd3fm7gCXNU2y2rIYWKXn2YEdjtjM
rF/88dOhK+TCkcYoy9I1ka3KsKTnRTrrKlpdQVSpVXQbxZEMS7pLoOfMyqPr3zXJuXXKZ5wBG/1X
jHXCXtZmJtsYY4XpbEFtPKVarjElgu2p7PxQQkOzetmL1rHemhROzoLOh5fOEKpS3Isif3jbWOb3
4P9SHxqCU4XdLY6abu/a6aYWE1haXeZ+E/OyLcJ1gStyZu1QGTG6qkuwcWhrn1Ixo1KGpRwO10w/
hSjHVTvjY14PYz5JlLFvld97WeEV3pVds0N5+io4Euz3jcnNDayc6OAin4E/cA/i2tvPvqbon+QX
ZPFyNrZuQ0amS3bIL+dTO1MghuGm10PeqyzWF0sV1BQII1Dfm06uJLioqlG4h04pANTYyiAkYeew
uaiHMhTulgmBQhRIkAtOLR2i9iQNVaXfX71evsaic0E43OXLVz3pHN19ED5RtzKsA9g5m+E47/Hk
LwVsCfwebD3O80lfhsiikOIRZcMUQOF26nanTnhffAknOEtXSG/CROlx3vyNbWjwHZf/ydUNWhvr
5djwHzyujta1pxibcmKr27bfkkuLfAm71J5DE8lz7LshP4PvCNs3Uow36j/y3YwNHXQN4bVQI/ar
UVQxem68DkdA0aVqfTI4zsIBMyDVj5PFY0hNYNWT8dh0Cb/tds80fIeofPhnSOZd4sFnAyeMZAha
2GJObxT1x/uu7OSFWZh/LJBR9v2QEae8W9MFS4QMBUEQpYhl/pY4SEcn/LauI6UWMa01Vnsrx2vh
dOBEmr9xPdThxI291RKlgShsWfbbMk66PqUeOQWz7jyQs1Ccq8/reUE3t1tTNNOkXU2hmGgpZ5U4
7Y/G8kCMyGvoP+lXQVQ6sAUcR5tFq/r1vut1mGmnqxwAlINTSQConCpBh2onJqNQPTBMgilry+ip
rgGL9LWphoRzQ794k1n0w1K2HLSmkRSd8/77siFe3DuUyWjWrmKjMmvGIY7xCX5RBptMLvVL+Ic2
1Cx+AH9Pf6ARVnZFApayE0kGzVL72ZZrJaJXYwJvt5lCUGHu7mrsOklAy1hPKKKdlI37NAMmw9et
LpxACrGUO8aa1tKQX7obrBV9cOqGTu21RlXje4lqqjDsv8jWXGSjqbTn4tP+D4ei3Q+ilB2m3QGZ
2TJ0dkM8lRPZYguQGSa2f/qHVuBTb3iMKHAVVkcXeFS/zJxWNCkN4+JFlcV5eFZ/fLegvO75YYOj
IDVXdwpuVcuR5DR4PPc6xF1ooAjNW9+76mm16mclklDo4mq7YMnHZuVWgYFcBAwVH2Y/n7KbvKoR
NqOurR+l16/pOAAv/DzOi9nd5gz0LW42O+XAVNTI3AIQwu/Q6hDCPDEM2MHYvPYi76VQmIqwRJjy
2tq8qHoa3S8exRQ8oJd8JbNDFrLp7EdoJf1F+uht2r8Mc9iR27yvytsStvnU0Gwe53iQ0zy6xQDv
LsEw5LbMy+PoUiRywf7LaqZBl4vsFRywdOKPtmJS/SQyRz6DAb1TmCjowvEcBNEp0n7aKYDns2dz
0/StW+p/aOVf89Pv1Cu/bKmMU27ZGMe1uDU7W9L+B1uZh2Kgbil7bXro4lO7CcBl1voD1u1PC5Mw
hHp1G6mc+rUmFvzRH8xdpQRfhPlai2coEq1BElgabeXnG5QlqdNOBi5z16S1efky7iGbhrRnIk54
IK3VE9CVkPblRjya0vJmYjGLgUClF2SN5xl5utLDwxKdikz/YVvs/hpqr9v2gYCbgNygwHVxsSAL
7lnfaua+u6mWcdaf0f4BJJBI8hEKExcvOY3hNWtYtYBu13/4a/2Hqx8QniOcwRfPoXAXCqiNvo2J
i2Z6JzDOd+EqzaWhlkrkO9CRTBvlWtYXqjgsrZiKcZwBdK2i95bdP5E/Y7TbK0vXIrzS/ofbHGuX
sBZZ8lTaS20sGhhtuYRr3T3RJVzURlEdmnNnTvqpDXo7yVbk3I0TKt3XKqUf2/znsHdwTR1jG4Dd
EEwXcTOve1QYc/I7nKo6ujky2xQKOO0+xGJEJWlhel9oi6fBEQ5bEMFPYXalNN8fVZzYmNYt3PtH
w9ENxMnbeE5L+zfSaY0VGgyoPOfSqs1u2XgRcev+nWns0uopYlphbiCvys3xg+F5j9ZGcMBynmgb
LXpOxB+I+JRt0dMx8zpwN95f3BcPXo3k2GmHHw8tsAU3cnb0mslSbqdiWM6X8Zpe6y38vuSpRbWc
Q9JZLZfOCzoTEgXGu+p5zmzRBwxQWiNPZEsHuMXkNmWHmmUuzSW/RESwDMT1WURpBvAymkkJCf+m
vlYbnMNVDx+MlVW84wUm2AGhxraJHeI56J58Qmjfe3lcSN4t7Yb4sU5C+Tt9q2VdLPjNhEEyTjOz
uOkgvXKXQWEZ8gkaDCRJhNmivez6Zx/picUPfG23YS160+NqapzJ5MrRj3rZ4Cu5um8s4VjMv1/V
hKx7Gp16tXo9ZyFWcbZjU8uLzIcYGyYf8Gr2da1wOX87Blkzdn+DSUEgEj6kl33J5S/vT6XJGmkQ
WzETLWIdSOkI09F+WnKol47jM3wBu6syLXAe9fBfhODva87T0tKfNEBRRISA+oj7+pC5sLQaNYvs
C/7UkcfQ58sJyrio8ddIiUeSDe4ShhAXDMU4P4ijc5TF/Wwr4zTCxTQAb5Nk+MhhW13rExkyWj93
hmOn00tQP6S0LYxjuN3eGOJAQQ13ghwdC/E9U+UzB8T4haXuD7w18F9WwFFu3IajW6A9EoFMlxpp
gyMUTBI5Wn1GIwfBAHYAUtyMImNJ8A/cvRTZqUNHjxqzhdsJPv5eW4yal22HPHGcUbm/4asOeMyR
5jcg52sNTPBT48P6kIPUEqPWzPbm9PDJ+bA7MbK+9AN6w7APylNcka28GK/QqV+M2bikxrQ/EA+b
FUqD7TcHaDJAGhe0yLsSk1sbCVfsxO16t/GiUa4oxiiDxhIOzLbV+G0wgwQFl2hHwsvnxd/CYYbk
JGjdpalz7mNH/uG5OcTXmmruImWvWrHaFNTxmQspjklqg2DK6fthh8sXAPb8WYVEHlf82MYeb7Kw
AT0KIVumknWeBeuhXcCPxK/RwE2ajfYuErJRpb0+rfCYm7xfuNhpWvO4GKbQu/Atzt3rgreDrTNI
tSyI15Xb+jCJUJoCxI5EIgg3nnYcKVC/pdWsgdrSzPMRy25jH3cuQwPtdi9YRwq25LPwnziDy7oi
oaCW/+VYfjS/zZgmm+B6WPSDb/3+HL5QDyzeGCpSU0FVfyd26JgP+KsGoRbeSz02kQbHg+jB6n85
/VDlohJM3kn/GPEuN/ZRLVXe2quQZS1Q3kfY8AjqB2cc0CuZ0T7qfdffDs5YGTaWmqkInoiXUyyS
wynuXaaDDueLR0CXBMht1RoolJVF2zXq1FAqSq6lkSaryfssUiidLkmBzBGl4cJHGSJUZartfRw9
1dqwQtBnykqQ9gBN8E1Vzk3W+PacuOUxiDE9PaaFejMEx40QcJgV3JPpZVY+UkZ3RsRvTTppS8IH
PdXXozZAvhcR1YN4Vc01FWxWW7mhM7Ji//qNXAjsOAscCXBee+pe1i7mTFAowfGmnQdBOwGkf2YM
vmwpJJyb9QiWMCEXQDOOg5KcPIEwqXHm7+risEpdEmGV+jKeRL3ssUfMaiR7a2oFlFnlGP0FUClz
NJ82V7MRovkK2pMuuucv+GSHzlcYF18ZoIuvOlDeFoNWWdMXI3ZUc/BTnTbVpK00SuxKhYUD6IGA
aI7uWDMozWX4Hudm19ZrsBYDoMSxLrcJSxoZWe6xnZBpn56gQCJ/xCK1bHEbA2qV2brgsiGVBHrr
5ZZ89qVdAOa2eLJTtfnbd/IJyqhcvHbow6UyDlmBqz0YDnumYk8ZxP6vPX/Zf8EutTGMYomHcXdn
jipIY4sRR0iTZWkNoz783+1IK3gitaRp0aSmwMOrgTqJ4ggckuwy90R1/Hl4jzzgSjUnTQzkysxg
c+oP7EXNAS2gakprp5jd2FZNeZCOwjuFTgt06Ks002iWGU5MhSev/XWOHtLUTbSq1ufirOKrtxpL
/Y1sMhoymYSe+7ni6mZ1x/zdSriT+kQj8JMOjal1TgdwZCamVs70gUWPFjqKIxCNV8b92jBkVXrG
XH4X1OI6RAZLWEWFYRraVwIs9lcK5q7hY66iEYL0fTSMU1w3EAzl7fAAGfyDNAqd5xuwEh5ZP7Uw
wnH1JTGDwxJQCqkyZUGryeg4HcagCZXBUXkyp3Nb2x+mEADNj5TRtNw9qD/5IYmmLoEsBi6EuoxH
epgEIJE4mLHRiPZ3ZNPtYYHG5ERAYYB8VTs9T1SfCAhNuaMIi1g58uWXzBw+/5z6ceTxX3KGAADB
ngwbhACIHeG9wXHthfhSbTvA6+mGUMcVVUcLBjHnX0XwkFAstwACgQq5TP/a4kUmRDdgTVjJfGO3
6IUv4uYYAhFCj/N2/UlqEltRmJPSo94LvRzCwjVTAhLNGhIqLNwAmgYC5VztYuOZlEl9YZPY/ePn
70Br0I22g/gg1Rz11zDzjq7CP+/HmDyxOamYuC0iU6+4aGa/u/QZGzbG569iCqspZpzx3R4vkolu
ithF/xNnJ9z0Axq0u5D9elWQ7+sqV01aHt4/RPPiUO3qol2PandgfcXVl2n55Nir2M3f0RELSYd2
NKl31Aoon313ZtMIhx09kYkj7baZevRmQXqKQrfEYWGFxgV4hyfcK/MF9HdeSXVtzKfyn05rt26o
v7jd1eLGV/F6xPmro35v0/lI3MBAYFC9Rp4MXKkTv4bT7Hkama37n62tBiSNI7t3a0WukuDv//z+
iUEdc3SSTpL8iohGmlNrD//Qk9OTpNr0hQsNzrpn4x+gi/azmFN52Z3VdZ/R6NHnHv/EqkI9ZRnP
2W763dwG+apdgGmkwrwShPSYIFT3KKE1p8UBsTRLWmqk78bzJrxKSBQls/y+lj7mTz+5cnzaffHs
XoauXZp8H/qJkaR03ECVbIxXZl8+DnCskp9yzTaZuyqq62s+oGxTTt6F8Z9x6LWkOT3BfhZHeVLs
X1yagbEZEBWIojpTtYt5yAchgtnawWuqFCB4zY2BPwsZgwEOVPk9aZiaqNaRlBeRaXw8sFpDER+f
s32hELD3+/SYq7xyci0wTJYTKWBAV3AJt4tcVjvOLCB3DdtNmhm/cduD6kPxggBNv7lcpkiYuL1b
n1rQq5ZRVtNY7IQcCCxOkgEtbFwFzycDqWi2v8cDx1wjRD0Duhaky29BK56kRqS1xwpR3xGKNCt7
MhYf9eWhJc7UUkYmRoMA3wq/gMkWEDhDts5yt5bmptaYCELMt7H/SekifdZzhnXZO9YgDZUDWFAY
O/0CODTrg6r66j0cy+PbaovmnIrQzUL/MDVTvghnoMs9eIecu+URosx+mpNtRWPZ1uRX8LU/z6Lg
KIx0odKeJn6KFxuI14BFEokmlBL5xSVV2i7awVkwb/oB0dWBxlQMAXT9qLo3/C4+K+vx3krmKnM7
AOObwFZm86SKhPECBLD2S0/fbFsRyWAmH2UQaH/l2wyrArhgaWXL4uHv39uMcq0lm6tv64jUzg/i
LLtHylu5KtnQCCz58LMvLGavPW6xICPPxTBUEsjbshox37IV+RTIkltA7KXwsNyFpU0vabhnCPct
RWj2SF2mICmOT2cGOlhMUqTZi97HGJpSzukeFC8fep9PTJcWyK9XrvXnJTCjVtgkBivOLUnTdf+E
WV7wEutvPEa5xishcK8LuktbUf57H1ntKgn2EwxTSWR+0x1sod73sdO6kmPZ7mcBigYusmYEm+4W
vfGGODMZyQkcAIVVG7hDfDpPhcio9Q15RZAQu1feie+LnJZ5DGzqEqSiYFctpQcNUeXmjxz+2O1B
OaGkO/h3BQ609Ku4Q1L+/EwVNcAHyF+EqtPIlZqBcnRy7N0PUeeobUaovmf5r2qiu7RCw/ITxPxg
1K3XtVr81BA8oxLwBXT6nfLXqN2PVIrSSZa2sjHtL/FR7oOFzG1tcm9lPZfCVLv15p5PqmBSjcPe
SdttXbgBAS4UqEJr5hze+DsMRWNRZVc0PrXQ+eO3sIB57YTF0D7KHERFuNlIzSBK48TpXZErMc7z
7+BO1pMoiHxt82xszyHKi/wnc0pCCzn7/rv5IafL/rUj23Pm2xDTzqOuiWP2RB7EtSPwxsMBjJS5
wn0VfK9B5pMzzCwEtNaU4SaAqVtYayZRZE9T5m0IcUp0HoMOv+m4dqoJN4nI6la5S4x039gpHvcP
ewrND5uzQzbx0jfT0Ws3GIB7TCDbxsqLclkSJBQvOZoTVGRcimO9XSWcR3nz2mn10Z/LKtfxdH3W
DNgNA4nJc3Y+2cUps6Zqk9DjiXezG1AXP7NvI6OIprdTwy7WvycrHuOspI13N3zWtYUJZ+N/BvlN
hMEdPz1aXLRLvnq0rdWGTTuxWK0hqtooM+I0y1vobaOqR9AyaB8lIcHcxbUVV37KhiD6GKq/9enn
SmfjvHXho3bLrtoXVVvfF3SWeUlVcraIMmBt2/shcY2bM6s18VKnfNcVLcpHN5MNYgFSpr+x25WV
XXM1L/x3YEvuRXNdt4DagiG+Z775oELHALiDV3rOCzKXHOL6c9IqO8Wng0fmY6xSL4v1UdGVEENb
9Vk1t5/OR3fVLZ92HpGK9eqKJUU29cJJi8XNUkzqj2Wy/aEvuJYc7ouh4O8W6Lgg7OK54mUrkuTP
UGb9ypZ9nzTpTWLb5HjW4z1w3SQI65K71lE1qYkxF+nQnYHgWps9BTX3+B3go3PpQGzeC6m57NFk
ySqmArQJXDHS3sPd7sGW6wMhjW64C5aeyFXdXxr5zkMFHlRNJusg7/xfmuGNePc8q2M2GnED/qkT
FDlY0HwN1Z/lEwkLoq4C67nvSWA9oWpCEaazBbUG3pE1A5/AcqSBXG6q8qAqad1oxx1rplaWAQ1v
f6N22W/AGLVaGhEWkxokJIwEDDSEgQiJ2JDQMeMNcEFxIvGzGdzB7VO68v/oSSqI/qO7kYJCFVIC
Bbd5OM6HPtp9HCerlvyhT4xKhNuWHDLh0IK0NoGSLgo1AfAA1CyaBgF5kDShVr22o6VZYeokrM1s
ILGNti3/pPSTh/Br/bziSUlG9a09agdp2OIztvUMHkxHrlqRFs0MKKFVuQuvikMDn0N6FnZiVu9O
XS2xImcrGLQpOINhqNV66DlaB2XRDApG5E4wnZkZv+CKfw6NJl2kTkbg6yBvnY/GzshtjjBNqlDn
u0XfcVlfnnEFinbjhsJyQ8wJOsLZ2w+O58TBOtPfFRNcap/jwAR3ickGTNSeYcqHziS8p+uhTK0o
ZrHiJK3yStN4ux1wJnJuYQLZCO50eWiccSecx95XMU4bs7WdaVOq6oKc1Ha9MUr8TS3YqMY0UCBu
Dkcu9ARmeAiiYUwJoWO4F55exS+LdpiMvqFIUa3bcKqhceechX5ydVgiaQjJFPGpIFIQpEv7yOL6
m/FOmDZcu7+PrKvQPnlY+mcpd39Z77l6nxsfTLBwPGLv8OvSe6SxnMgSsQ4AUdZXb24b9umxp3B6
17nDYcGOoXegsRLEJC8+rvqn2yfn0olS/GeiW/73l5UoRQhAXezoqIE56cfsqaYw4Xl8bdHbRkHD
WOPz6+XdNowdN8qoV4s3aQVNn4hDVUf6RKiunWA/ryD+EotoiQdwA6zSnFhc9pP2FzyAyAMdQCo2
xCbNzsW5L3Sg4pSJirWTJzN+r4aPr3dwx4YfpWYtolrC8aAiYmmu58DvmvyyleMu09jvXNYyUV2m
Zd3GofIXm9gIZjBowJ1te6otslKifME1xCs6Z+xFo5II3n3K5G1xADCGt0dIhKU6Tqupv+EyPcyi
JDOk6VwS4f8M2ElRknHAfokLXzPm8LmQbs09GjBQ1uiAlmQTX8TFhibyWZ6Xew6ji8lfSlTOm9zh
JTNfoVVuwG1WBSIK6yyOrmyyD0EL6hl0/g2Qb88aWC5+GA5opyaS7oNzh+Av3axSGH4rWdzINIFM
sGg1i+puZ+YFBXL+JthhkCYZSNnvPI++k4xce1rhIGqBpvAzzaI9BILJyXFgBF+D5PsJmnsbX43g
9A2UEB+UObHa5eB1o+ihz1QmAeGspwPWPHZ+q0bz0uFQ1dwiaRhZ4BHJgOnPPvGWjk4T40+u2ISS
U2KfBgfhir0h3q0RAB2DRU1iF/a9PxOwAkWTyIDC8E4hBinhzGJB4YFYNbytpVmeGub557E5ki6H
EgIiK5qeRQ9I07mHuWi7Av85aGYlAWhkwGAm/vJYHdI/H2surLuNlfD6s4X+RjsQIiNGSxDim/1Q
RjRIQ1uEu4OfJbuRjKPRC/gr/0RfKOsGeohY1V2mbMhtgS1CNuAUzP12a3xGwqosVf54bYSRNrRj
M3ZmYVMd8zc3T3yCk3Tc9PKJDkY3Xp4+7jAo7Z5hJMWjXpQXyCW9oec4eiq5s/GW4o7ovQ+LfN5Y
aWPxGVvOgC7bJq+mMWebO/TLTHfK94FZEFbBlzV/x67s3DjwQm0604Klp90QwkGrr9uRrG/o+VwV
yq2y7M7iPxf8lbw/7f2cw9ioMoohrWkJogeZ1g5I3OQIKqO/qL5gM1h2pwCS4JiG+GPEkNmXN0Fc
Vbi6oRpttvEjaNIWdi5uigWZaYJUsHVePmnDnkusHH8b9BWv8T9K1W5ZPHLbVyNQzwz/H6MNKW6A
dMSjAMHC9ieEj+VYIUZXX21YC1RY+gVRpa82psLzCEpfK8Q3W/e3xLhPq68gJArzh4sYHcnec4Be
8nn+Smkz3s397LeTtw+sG3lqt8uZkUSJdRkdoPod65eDj54hGGV6xqBsCqJ/eFKnUjOKVnJbdZ8y
F2D77EAKrWQRdGN1/ysLgjQwCs2UJLkhrLJjmcfs3QSxnGycGCctIYO9qhkHuCvJ2WvoiNSfC6Xh
Ed8i/xmzFb0tKxEkVn34BGoZdUXqBzmQyNWLsjV9j/7526qxC0PjoVg+P1mjdBIm0tJa7Nnuqs7F
YKw8YHKjA5hpcWl6xNieg0U+9UQVLwgygoAaxjdzYJLlJEuoL05NNpY5YvD6EagTWBnYkTYLFcA1
X658Ui7Jy+KmBY6/gJJWEz72WC+M1lPwpFhn3FvZBJYEd6KShwpyVml17/ngRUZTra9ahfmFpvvi
VxSHyEygjtb+P4WKP88GogZHB93iyM/x6fpxbUFmoueeox0CBPlmriuP2Y5Nwxagtrk2AGFOv2nn
nVL9IrWz6YPKm6TLwJ54NSukX7SVjnj7jFSM6+akjk5Fw6NTbCQr7l4glLuzt7YUYXjBUuvRzX66
M5o0l+cBh3er6ENEu6xqKKkFW0Qu0zihaxOCCde5UsvTwrre7NhWwratafNOBQNdLeyNj6XebO4k
DzPhBwqzKu0mOwMcCzaR7EY0zC+R1dKv+eLyocM4+mvxFOiyq3IFx4vNRy/JOssoQLgAOAPZDqWt
9gYRxfuHHEFw6j0jqBq2Jyb7MJSCSONh2wOcYG6CDr/0bxK/JHfO7odPLvftECgkWTnqLSgy1dej
RG78qzKevOftPWdM0/RKsCrcPZeWyMJ1TlndhHDBLy96migSq66SB0FafEXJ+Eu6NIDlkR3/z8Z3
wkEgMLaO43D39zd2yELKpSMS+RWc/b55OfS4XT/GrYZFmYqnJdxYZvtVrQXOnApAXkQmGBq9uo7k
m96pF9XZbrxBn3gDQbiDWnJ9jDcWLJdz2Dz8lNjD0RI3ENyp/4RRE/JD8idKkP3PiNKGaCs9RQtk
idudQmS1NLs9fsr7SrpjNVeO+L6QiqoWhUJg6Ud/Fh1s8T7uWrZY1oJ3KfHvgluYtCtt1608srgB
EbG14Wk6KUtfvde4FndWMzzBH+1awE6gHyJTEqd7gcE8pgqbotegI1+1c6AM/8qPcQfuUmqRvPgn
F8ZTmk3Cnu/mDzU4EgQnTT3XBhI8zvkNtXvjnduRx+B/2TolK6PDSa4E8yVqjRxgL0C7kd0905JR
05eVIPa+OIs1FFge5q7FGWK9Sw6Kr1hItuJiF5xNOpOoZzzaBgxxiBQcZ/VHcMfyMH9h1DcmANaj
lt9nXU59avFVxqK21d3AJp9216ZKfmvyW1rcSW1lSD9i8UPEd2cTkc8lg5zxHnmoJHBIuxONp3rF
wdSo/jbtucn5t8GzqpsMOnevuOFKMmSOaUa0d21dKJajy3/lWiah1Fzm9oHQB0lR4J+M8hCxtWv9
Z7XTviEID22FOIjpyu9tW4JZL4fzXwPP0YLHoqoCDodQcw2WjcL5D98d01u2Tc4K3/0AEL3V5THb
Rly1nz+IHQ/owCTM+1fNx0ZxAURGSI4FpkK0UkNbN24D3eydVm0/QIs9OxpTndDO+m0ZZA4EUG6w
fATTwR78wHPDQmCmjMNJUGF5NnP3P0XHk17iC0neK9EUEiALUYO7h10WNTppkR2WzezULL8wdVef
LK5iOeV0mWz4pFm3zHKf1zM74qXPfxYTv6Kf7CnqxTSmVkIuBVKuwynGGuvyBc0dMUByl0VNOuGE
QGDYZ2E8/DGu1zfsXsxyBJ5/BpE962xrAmcC0Tg1Q38qx4CZ1wCGcpzyWIMpWMg7y6pmMCxynEOE
onTDNKY4zcQP1tzUkUHxATSfqNqIJZdhYgoD5tvvJ3fhV2QFmHbfNKR9Q0xR4FssxVTB2dGlGgc8
jnLljnUXA7MtZ0ZSXdJFTdZC3yGgmLyLg89V3ABDA1BTc4ckEcqoV7CXiHlCP0HNjiVhkzw4oMJZ
g8exBGsILc1xuRzIGRN67xo2EMVwqwcZanBurCZ2hVihvkpaPqSonRCpUxYaWnBB2q2E0RMUw+cw
mYJh46jpCqrK+2/DW1y+uS/B1bougiVTbzG0vAC4zpdi/TkoL/QaRteYhNOl64WpKT7dNTXQX8lY
NxLlEGw9wm1h85YoSfKOvxbxk1q3WeAKXW74XYQWUvlfxeFRGilA5E3MAaP0hJ/aKYwk6gYzfe6g
PbXjkscR0484nQAfvpepwVgmMe5TQ5AQlDcHeaY9vKpROfDlYP+T8+9ImfT4S3wxYlBLaBJ0iDZH
h/WhlKJsLcLzT0FVy2uqBEXhCCn/LX9dQ8On3HtImIRVgVaOCyRc0nHbLwoCExpd3Fin/GUf+YYl
2r7BiS3jwNZiU/0kasvUv//ao6FY31IwWPBgD7/+YguIuidkOITEjkkINXhWreNJbNzT9twUH4tS
lpOcZaAsbI76oTtrllund1X3bzjmkGJfRLhrMEkoHQQ+cbS4MfElQVrgjTyj73eoRu8ifz5AhkO0
Sp3F1lSkjISAJQ3qlgmYggiJC5qKyXGKF0rqiJQEN86Ibpgq+tme/4G5iW8YQybgPIYffTefdKEb
N/dvjGHcp/uL7+nBMkmLFVVUIXtPi9oHoh8cFaTXjkG5lUaswFD9VzeDL4F9nh6R8Vm2GRTh7UdE
KHtFuSon5GkSa6ZYpbZHDwI848STefAyL0xkVTtVndV463o3iwPOrb6X/uDIwttx6bMvNoAU2Wjo
ZcKBqg5cn3xW63rYE8F2x8BXbCnJovFA+eyfJLG1Q2w4jMms+W4APQ0iZXhNgqVD/uWGsKsFn+5l
MTKpTDc7GboHTbez7Py1/ICBxR+RSNsEkP/EPca3AGnDTBZRcS2frR84qmgSYbx0PlIHJnbvSn4p
YPlF8B0GNaYHxwuyGWjePKeQ9oTM+eu92WOQ5HdB2cYZhV0Zqlj5xdbdz8AJclxUYiCQjISR0+e6
DZ0vGykrXRu4aERMfrQy/rrkjE0eMdD+Nv62we7aEe9fVFHSJp7mHpDVbxPk5qSjLgl4O1HSIfOQ
ruTI075Rk26rps0i057fjHbV3Atwj5TQhys1HrNjlOjCyhBcjWv9MbEAlnHwvt1AX2oxxf4sZJJm
Cy6seIGfEEvz3hKKCa35u/Mw9ful4Qf4JiZtm3a/l8FEa7+1x7Y4BL+imOzdwzDG7CM77/8auHtf
g8BIkYRajoazKKKcvJuFaEACeGBXtAGqjGBeKAGflnIoHav8FBI99gvllz3KyH5q/QyfmYXBiq5D
OtBrhJEL/sMU9Ct+kiJlvb+/SG0l+KWJ2cZWJbUqkNl5QeYqDjxXV2olxJ4Qqi7eYgeSVItWYsrx
Nhg7rWjO+UD5rFjNYafzgclwN7Crq0ZhQLOKKaEeWSVDeDHm8e3ebq//2C6IcmaoYzS0U9QZA54q
3WemuZ7kAVLJzBCUe5p3lUrIIYSQiyPtOT3gZh/hx20ia7hUzUoeJQK3DQ6MuSqDt3IDaGwEq957
N3RtxOyBJuK8j43urY+lHniY4KQ5531Bnd82qkS0qAN5Bz+CmkiJae21v1QpE85yN7ELi3JFp1zl
cuaaCYTPgRSuKiPJ5Nzju9KTMmKzf+rvY8Z5OREVps09aF0mLqicA58CV/VM0fKA3g1siEY0/P+r
d+0gQfEVh0W1J0+xayQge2otesLdSbqryrHTRc/uN+TD57G+dxJ0YW0KXJ2yjVL9eCKviweB735p
gWwEDHQZWorN3yWhBXtFjLiQpPIyZUBu8J4wys2Mu0thn4auZqkHerB7KB1Uhq7uQuGvXENq4Mt/
BxedxmSwsHU7aI7lBoGrnohRdE7RwKSjwZx9LvjPX7dQyR7AN3FW5uJgQLHORUeVsvvFvIJ8LW9A
rlTRn3olSS+YdBuDwqlKBZKDvvw5DcDHNBFZMLnWdQTl0575ekZEv6umYHmWJ/QHNtW1VVYlglhf
aYyaR6WZ+B8k8eLE4kc2Zo0sb1YGwcr/nA1dNaAKqRJ/7vJHm6cPNLeL/lHO1ohB8+jT0jVSuEC1
00kXqjcPcIIxxI5+6cczRLXxsWxeCxP2dTcBV5ZOrZa0HTYbjrN392DJhXbvBNRtfjg1/APyo2A2
0FVKTTXG+q7dpv/JgYrFKdnJfETHAHjyr/qxAdj4GrPpG+8BVT8P17ccsHThyZURKtAYVCL9DwYG
aRMCmoDkOJykWHk6FA38S6h0bkt5PQ1zN3QE0uX3lOJWrCCsT1MsMjfUhfq2v2xK8pmV4OBciS2B
vt9WrluA4gfcZicndgmZ6nmzDO2phCRqOyNhBOJZ2RYz6JAl+nEP3mr1VLa+09nTcrBWLvNmKEUi
Q4P6dGglBhxrAZjPMy5fi1HB1cwnSxqWhn9MhUfEpqdCu61CRAy7sXKGCHu11EVVQhsAVA+SVp/s
4RXs/RNWIU6Ok9u9mTPpxDspHZr4pfJ5JHOTOSr2PuQ3+f6ltGoSud2XSXhmRDz2xGo6zRXn9arK
1R/gxm9QsCa2QddT6iGcbkxc0BEsBL3oyW//xCWYn16cBcjAeux7NIz2yg7b5ZpRrm8wrr39BiH7
VdH0zd9s8GAlO82KtTSnhdWJm25zGg8wudNtHWUFG2nTkWKxI4vvHmrtHZ+ifcSVfiZN+enjtJmB
qAeka0uzCOuTCOwxKNs8mfs7ZGzoEtaoAsxb9djTVyGSduGfQ6S5xcbN7+mUIgESW5Fxx0HjPrZ1
Zf9sthII87wrjVlYLId0nqr9rujh3DnbCyXF/PErJt2nn8TPbhnxxz96PHI+WWcCPgNmTEA9T4E4
9U1j1PFtHMTqZHebbZP7crEHAWSe+1z052GNuaTKwH5vsHcMd0S1pQo4SHGGm/RqNyVkbViSi/lz
bMRGh6lgbKpZ/hlsxbv1C821BGQhUmszhciorVJXTVSTL0hmIp0vK8NjRKcUgiz6mC64WVZ2nffP
VVg3EHObbcU+dMkpH330V1VJMJKs5Ac9JQMHGMtugOffELqsAXyo1G4wapSsFFyU0Y+0H2ou63ZP
zjQMHukxHZFli1GKC7HEmxMSNUVSe3zm48A8Ueu0efyLENabNj3xYPvSFj/36XkWg7xQE7A7KVtw
zF3TG0e1tv1Ws4aO8jz4aNUTBHE0bYUVjxxhMqlNB/CQ5jersf4k6VfSL364+OF8+NZoFjU7I5T2
jUbMiA9GtVUr2aX0eZkwIYMEKs8NBtFWAH6RdI8+Dn/wmwIyNzRxtIKklCJbj6Ok5zNPqS+jpvVm
jRLGmJjGsefI66dzFlgstXCBTYyfF1BT5P6sgyPIpzbd4ZqMvwAFQRdfCIHzXzbY4B3CSHYXMycv
4m9KTJ4kcQCqyfBlXZNPs/1ju9kYSKyazBTC5WTd847IrAZU189MUWpTS4cLHnRwUXHGwn3sT16G
8JXKmaev3an9sASC65u96tRWU7Qaeh6lHjqZjtis5JEKSwElGMHb6ZCzgjJhQVN+hQmGkJVbat4l
mRKDy4DqDmOE8sBBwqORm1QbRcoFal08NRXKFIH8uFD0+B4KClbmKyPDFaSZd7QcXRnrvGkSKYw9
AarGAzfWdUpjVudETVJfQmuHCVkqvlZd4inNRntwB8pYhwWUdCkGOqqkfY+9TiSvIAU1PKTTXwlV
EtqKs/ygMlCZAaLOtUEnZ5xM6cBIKXWdKXlzOdp0pOaRslan4Q1b+/5d9OXEnMtZsYquCCQmy3h1
GiBi63kCiOlnOxABJMVGyYN1Fz4yNBfqFj0FUTq8TUlEBRZtrv9ep2HYg8fHTEKPvKujWDyCHE3c
/RmRlqGJjiPrYpDoZI3FyTd49N+v2MAjENPmJZ5vmAsLjoJhnVnW+kfAMI4ykzCckrzfA0MIJ7IH
LnN2PoXx8TQa1csoNhdD4iEHBGPLD4lclMqaY47ENcic+FfUHUj4YVrrC0bmVydoO4sWh+yeOFww
yaoTCB/uXqo17x5TVTZFhbZM8ebm62PmDOfP5Ac3GzMbCwt1RfZQrk4uD+JozXdTvAQa7faW+AgO
7rYK+tHDLC19+wiC6oNmVN+b4DAHpVH30oDIusfkH/xMxDpmk1QmKf50AkehwfW/G6YVtg70Hvxi
Mrz/3Typek6H4lnxZw8pr2mn5WVuq/81ijPB3XQMitUHhB8f8BhICXgRRupuqVVM05gT06iPzBgu
8Cm6gE1youilSMdHoNNXkQnfS5k4pgfpfMuAKqhc11v2e4TErAKBKm8fakDsNnpP6JubMjyTfmKr
gK8selVaa8QGsXnHoepEf2ZFzcAa1sMh6WosxmKMc5CsCRHyFqeQLCwuNGrJyil7jPKOG6N76XPY
SkjX2JzgmOKD1BEOfEBNKMyBKU6ebCsrCX+wOXLdKHsZcE8+/UnFML8uLWcJVUzadQnEnaLwxgiA
8IoFQ2cbwbTJDhnob0tWrnMEafM8etuZe6/kWJJ83qZN6TygMij0JiH1L5D3xUlmgDRP2nJFVQDi
BNcEu9LUQR9KA9Wp64hIv3oFybwKyCamwStlbVWT5c/cv0WU3CJidFbjuUaU73pUn66kL7O/G9Fj
gD4mFjt7ivLERWwTgvLnW0I5qNUfDLrXlo4UT+Cd7u+8f4EN0HVZ0EWtMAf1KBbR3OhqHVAn7w5M
c32Dv4RDLRW+6ECB3AsAb++2XDBiOeJY57YvPVix8Z26QqULJr9xKRj+ftZR56ycuxrboAcJA3j3
xRTfS25OsUmBgi7pPEQGxVB5gp8yOKNzZH/QyXK6qt0OrU+wzIE33WmmdnySM0vyXeOONi+jhMLz
PqTySDML/VsPaaBVcLN5TcU5qJj3VtDYnh7uzB1wQJgwlu19DhMujQECYkCuag57kiGw+aY6eSUu
WySK2rstyCW4o4gibyw7yVbYrZf628QzlHLapNLs1s6CChi0LuwKYmP1IJP0soTfCquP4lc274RK
Diy4N8ryYlzIUah1vM5IaA0tQoBvQ59n2dcLnsc3Zp0MhMVhkJFv4A1Pavv+ObpXKfYhsPhwBESM
4Fk7KrmoOmCfN/Lf7M0nrJhOLIQBpfobKngU7x9sBOI0inCtVhzkwCaakL6Sh9Q+fV+Uz/Q1o1SG
V+SavQhHI7nK0X83371uir+2Pu+u7pSkdsJxaL9qcAqbdO+e/X23a6vbTjRAftXLq1bxloP4mb0U
P5hA3LIr5IR1qHrNfF9ZypS/JyKzgdGyjieQ48fgV8+yfLQYAto0SEm8wCVx88NkztQTqwSRslPG
lSkZ69Ofm5vWt+z0A5JjM5tKiDWwV6LY8KFpNsobEBMXIL7MvezFJn1CRcELoBddDWebeRJPO0qR
/6sulNT5Lv883QNE6N2cuupA/szkEykHgkb8OX65mFJBCTTh5zl3YQqvI641djGpELey4piVS0Qf
Nhz/iaX5gUo7nL+xkXNxLSSRmuwveIaA/FZyyPy5oS4zaBhUA5Ydih2yNFVI80onmcor/Wq2J4VD
A0GXIEDVnMzXQXHgJ6gTRG3W98AffLdwrMHY5LQTXfng7h9EDeNkDUJbq59Z3o7hBFIkhSjvHqsQ
X97I0DBsRdnUREV+GWzdudA8ER7J+gRGpxZKGxJ8YB4283cUg0ulhcOT9sHh3tXd1QG7QK1Wt+GA
poBHeeYTN5r+1yYYwoYWqL4Ur/JGX+tCCow+00vabdtklWw0vNIAQ1id5h6KR6mz0Gyo4+bpDyMD
7WwiRmNzCpqohVq4W3/gI9cQk5Q9lyQ2GJklhv06Od87TxN7eSHQ307dkE1sfXZCatHxW7v/uIvA
S3QdSfcoc9TWH2DyHYOnkB40ZWqxc77plUUKlkEy8Mk63P3Po6YONGc/91wlzd5GlGpJG9lMzbZO
tEXw8ASgoTFi3TKOfdLXljxAspcqKKzv0So9Z0R6pa9JoDFUV4Ylnb3sgRQAFmI4SMuREzgPYv06
HSfMSwztiJCc2G+odfmG6ee7mdI5SnBRipnt2fDRLKnZ3b5WQnSBH2+puCEysdpoo4ZisD5/tQ8D
RVPOdvpKHRVu3ALA2o2jxxyIXOlfUAXmf1bOSuvBK1xLGlaSKh2bn9BZ+mQfBOsTzGO87n6KgQMA
4doLn+8b9iVTI9qwwZKZXnzNhOIXXyttr1CtaA+Xu0OxnWVnf6O+oe0TOfaZ54+qQgBeGCUdELLH
DSZ4hikCxLB0m+xmH6rjuC/WARCxMi7hFDHNoTQr5dYIMAL4iklFBFu9omPYv9F0jMbJ9a0//XJQ
CoiowJplBwEKgEK1jhvO4EMb/+XqxacUKf6M34o6onzYjCwS+yqNRXP+jNXtFGcRbir+PkBmWLTw
kcdk6SYabAco8a+iG+LEbECrsK+XrcCMuFIciEC4WU3e8aXVcyA5J0max0iqp2ZlVDgihInEUl1x
kptIbvy7dX265eb1UNZ3Ms/rN/+d+JYq8v+qqk7uvyXtMGN63of997IGJp4anJe2vXheui8g8HxD
qr4w2TIYoHF+UNMtQxEGx/EHylUw63tsiVJfv81oMwwSW9zStCs3Z1BQlfegxF5mzC0pRz/Mt2EV
rEGzou63pbIlT8m0R/XUUKxMqa3iRDY7MnZmm34gpro7a1VR5sYKF6bAKjEJIXgq1ewSYaIX0YLw
tkA+ecMZcbVXHTacYkxV7zwVMwfgPAyZ893AdUZnsgIDS7uR0wxIbmrP81fgmugjJwQSsQXCBbBB
NbloEces0qHlPIbKICnDmX8SxgADdxhDrbmD0IOmv5GKCBVC4Q4AfFcD6HhyW8IDsKVb/7oMY/B9
PBRQFym8TKnQsdCxjW2menRAClS9U55l7FuGS+u4Rztkb39oZCYAk/OPdZRi2zQcg0sutX1ME0vw
KKeG5tNKvGaoXviIHGicD31kendg/btfx/tPsRuXYn6e19EHFikBrn1lfKlmEWPq2h1E+1/W3Za0
xNNg5jDh/1DJjy+ZjTdjtBvXQYUN2+E+f8l38wqPYD6yMyzMNS7MqfjtPfI9lE0nBHAc4wFzKD13
3LhCdmihqA6BGNj8S9C0MCv2nV+EpVWc/0cbdE7b3CmfBgwqtwW54if2CYVfOej+uqXOIpw1hfdT
qSaYaeFomxlkMhGEMgkwyMLB8TvXh5dNSNlUKPK2w71Z58YFqaflpRg6JA3b5w6keMWR/RelrY1J
8T9j2Ya+lKFY7GKhbTdvRkYRC+ldjqARnx+dOXwlE0z1vEJNkHIATUDpds4ofewxvaTKvf29kk4u
Kgxuhw1YgHEctZj7uPMf4BSTqHmvVYenyJ7rLoaeDREMylFQFZ3ZqcMJNedLuuF/W4P31ZukLZLz
A11CMceVkn79kScBS+NALgCA56r7q/ODrEIyt2g+PItavha1bUjkY1SZToFCkriqKcqIQ2Xo+ghZ
KiuBcShclaTQtPE8giIwjjtXai5HH4kDlajPZdtrOLw+2u/cGvpGte+LGe2CdmENsq8fcWopKyWl
quO28oslTRS187B8JvawWpYr1HL99QCwIFXnXjudOSZckCNT+AkYH3iA4TAgKLn1LqOQsfjgA0+R
E1G0zxAXDP71OM3wstnKQD3Zqtk3NYg7XwEYHeyZOBW7xWBZTAEKhhWTxIaYVBN2jumx4n7GSjYt
TkNinfCLSIy3O2TUo1yn7zAtkYD0unTDXclRUYiWKWANpMZHpWG1WBv1b+iI/kJeU9iEGH/vF3od
ZCKnGp/supvGX6DL7WdCKom22NUS+ylqq65/DCFhRZdvQBMujUXtg1DNzoLx9jDlQrFOUiju62A1
tWWE+Ex0LMCZEn84TWfsY+Po/HdmfONWLvy5cRFAVDl+E8DRPShYDUIKPSO/pxCTugqgyqeMh9DR
QDnlEKrZxOAJbD6my2VdaFl3A1VoxMvRzK0lI5doVaZ0C+55mFjEiNfYMr0qVM5mhT7zZTeDLzEf
X5B3cyj6xnDYm0eewinvOMW42Zc4LhmtVZRgNfvLcqBB3lEREcwkMnlKCWSetx12+nm/3fRrePyp
4He/7AhMSoBCL7mu0zuYWlq16j0h8MwfWx3o7wYJWm32B/wQ/o7sn0gD6dvnVAfxPQDRdBWDIjzJ
NzMVca4rKgdrM1lXesjaZ5C5lE/RWkokq3Hkr4JnslE6FiBx29/3ubGZmolqYob3JLDOgTowK00u
nQ4TBUi2fmJKnvmvDeTsd0TiSf61PDHNQkZpnJVnGzhQNz9cJFABPntKUJkkGsR7f/gxk0XC4JIe
kOCgClfxBtAn/36kKsWxF7FVbEfF1fQ3wv67F+uN7i1GXGqSvyM8vrStQxlAXUGPm4ZHV8KuoP01
4W6QMUHsNM9oVsIa38BGjyapgYz1DR60t2E599AOxabGxRlOy9cDeFOQSG/KNOBIzUpQvfZ2f7nj
hrDYggMZLVFj9pYzdRnfVPXkKa+BUiAB77baVocy4ZScWyQ+sN5PX9nwBDkMNwN0PAGA8Fv7FtHK
peF+BEjdtO5YQdSlLZb4cu+yO5ssPiDKt82CP7x9L7t3H8jNbycIDtxseVuDiecJVF+yP8VCwOv1
MGrQICjAf4MqACcHTIawHAAJlcSvFlw7VrXW/rY1UvdgBBZvSTNKGzmPi1HcdDuVlouat9K9O5+i
FtQfX2UZ1z1Io7p+On6jby14ITRkxQRA31HF9hxt5euVYNUI5S9mg8xwp8Gl+JsxJSkhaC6sgjFf
kCLgvNAxrj5G9sNvbp6bar2GCCrXhL3VyX290/gc9LLYTTltiLjMbkEGTKvDlqKdvBpwMGzo47m8
9RulirWy/ID/xXsiHlidhGP95TGw2hy80QqNFw4Q7eLne2r0XStubASIHAuWKN4eDBB+CehC0sEQ
t+LV/TZQT9qj944SpsB063IDPxKweZ9B2mj/Avwh2YNck9isYbHOFRpECv+TOuvqNUTkUW/cI2jX
0rRQjDYg5+a7DbJfOeXY5p1QwE++B8Ms2I+Dm26pPz3C8Aii1CpVqVFMG4WnVl7ETembXuwV8VfG
RN5lGdh6+SgkKs+qj++VwZO+R7Dc1vgbGobuMl/AsO6uSJPNcQNS+EwPdGtHQSiwDIjH+TLu5NZa
ZsWeY9JK9bYYh1hOmvJqEzafx2WAIyHI1ZdsirCBVmrVsPigDjpmGhZWfFIZcjl38CBHF6zumk3N
3aVdCTF9zr03v9VN9R6daoeT6je0Wa9mPKc7t2C6fzJ2bBptJco0NqnOSddsSez8lK72doWiKHWx
5csVgoUOLqp+Fz87vlJGQoUDBrf0mviYvQimykY590G9t7H1GXJwHxOqroMBMnzIZUFjVL8JkLNI
XlP/n9MTv3hkeUjL63RBu+4MV82XmxfssnJgKoyEzi7XZDTPPqjiTEjqBrDtH6F5trjdpfRBNgQp
iWKQ7A5U446Xne4PaoUJtziS6rQvW2XUNADmOkoDqbacNKmIxkqje0NsZrHQnduVrsDms5+0mIxK
iC9K+T2vt/9hrKVEESRsCKhayqAJdiQ5abu5B4XTCNCLKogAafk0upTjJ5l76vGcScARIG7KWNlL
EB0kCW5I+tTYZF5H5nlZsdQAqNJcNNGqzUUmsdlZHeDa+NNmzSZry+a/kw3loG5FJSxxGZNLLeME
L6moU4vYwVn5PqtnRVj/R6KCugvRNalaqrYomLc4zetbAbku4MbHSFKz1AM1hBWb6HKkPjFWUKwv
PGifGJ9SKjX7xnQu+vhDEYUIshGr2Ob9hJHqOROUOo0JyJUT98gp4OleRBKMGDNRyF/nFCfVW/YH
IR3Oy58bPqADkDF7toaR0rRFkqk9iJSfmRJf5U0uG4lKLRyqRSZWDNRqnpb3w09oPusnk3xkaAv7
qC694AGkLQZE8nu2mzrKPUHta928rRL2ddyiUhblReF53BiJSjW6wOcUAED89reIQUDB5txqmhPq
6NSrst0V+zFzu3T+FOE1h5wqiIViTwANW3ty/vRTAzHz+cWtXzty8po1uVNhmshrFM2vhqOogx3U
/Z4YNLtcTHm+XtA0RomXion5thG4TzrYZQkXMzIMKZKXgE1Mg6TKtAwXPHUplhHmnXVDO/wmBHqT
R6XxJ3Q5nqoauL0ejcqHhBhhm3zH1FyoVIfsse93R3E2tPAYIwM2twViLxfhz1LTVehSJvYXFiLk
kjVej0hcAW2gFW28OzMsxb3K1/X7Cy++YWo0zByLkjsZzp4aEjZ3Cj0lNJ6+fZEZfT2HqMrEx7yc
aGVU2jqBWG5HHiAKUC6m7G7pt5uhFNp4y/JOFnsv8BvtXQZTNnGYeCEScqIuQngHGro4fD+zI38j
VKj1KkAFYYwKGAh1YsndpGh2Rb2AtNdLGVWAcFuk1tXNCEI12OrFlGXxP5baMn2TYVXarNbGfZeM
UC6EBtVDQccPGnt5CofibPt8PVqytTXoNwLJR5w3mnT+BZlSeM05euyNmM6fRAXenIWVy+PuMpN1
1SMPpzadUqixEHr60uYCW5RokHtLMCJN0YKrdhfkPq/hXUMnB6skTHdmSLDHX5oikZ7yd/WjMbsZ
A3TdyEoJgk/mBEOaZAtIrmNseWX0Ej62Uf0iVZMsbTsIEO21C+IebypEikW64orNN4vUHtD/6Elk
X8rQQg89aMuJ7SKSnaeWNQ77mOBdaQK3gntGh07W9qsR6XqlmM4Z+L03BiFSiXyu1QqbZsHtsInH
eCNLOnPPkb1obn57wLTA1FyrrwUxppHdz9+bOBtWxgdBiN5DvOVaPOPXx+xWf9D8SUzD0CAIA3CX
6ryj0VpKuPCUPlgbxwq1WGHULyu/i5cEWH8LxnbiSfGHki99tHwRyDCzYLXPurlXu8JG5VMk2zzK
yP830zpRzzbI3AyUYYSy0RCeCoytu8Q6/68fy6iUkxXRiIreIxvmaxbY9oScbV98ynRqqDYUOOTZ
Ywp0Rm/0uuIf0J57tV5khGFUjlNDiufpxD9ImVC7pLgueEVwvOxUreffjwOUe6Gm8Sf3b5fDnJRn
FiLAqmMbh7oJiPzt/IUiBCAsbUJM+YiBRhUCWDSpYV02ryjTAP6QoM6gyDlu46zIG8r929nE4rrd
YZn8EWLz+D5tNt+R3L9lX3Y5L37ZTj2lONa/YsMBpIAz+8lRJUFEywzDrkoj9f/3+2Eo8xDikgdH
EVFVlvbsMp8BuHFSVJF+FTkZHM54vLlZJWuzKZn7KAGj7G1WGaxd8HYqPEWgtbdhrrkircU6G7lI
V0OyelIh9i3Lpd7a4bqwXesZV4wQOfGV5SO7T/N+V6R5c+zQY2z6ny82ryeKS8443gWI6n6Or8vj
AiHL9vJHlMM1aNUZGa42+k+LVPFQUiKpEGi0wRwsUar2qdnOCQUmklRX6oW0P1PdpQe1EECyJgb8
ozk2dJsbL+8vXySZemaEnbib0zGMU0Ri8y55AKNJmPZ+PYF6PLr1J030KYvDrtElTCwYM0pD1xEa
t8vzllZtqOzpMWamcQ9HsNB2Hs9P80bVEPpol0j7/PH/BO2C78Vt1+0FRo1y+MMGs6dHxvivNhf/
dOD8Y9fb3xJIwhRKsMX38SqJja/iHRcsOE6IMnnNFRJPy4VTRXZ7NTCzFrw15dQJNS+CgMiOpk2r
tQZ3PkpmhnnP/KloUaWF7FXeVHAySwnSN1/RwiRmd7/pqLaHSPPCvdRkb4GiVPOatbGuXLDuoB9r
DSq6Cw6AZru1mnoUg7KDRE/Vk6spax8yGMD1fQCfTpHtopj6XmVASy3dnKkT01CeDqMXR6YDB6Xe
PXunJRUyYeFgcj6wq5VeIokw10TX18Cs0iD/xL+NUjWWvqDhjW/8bNFS2gmSVsYCnWxiEFQ4x+AX
MOcsnEHWTPixmyGMcWXXWWDZIrS9AZeI/3k7x+Lb/CjUhWBoj/NH0uI5SNdVUmhoA81JTfac0L96
7lAWPPdaeIr1+0+F8IgZF9mc65n5atNpw6AjPqgwv0QjoYBUOOkHmWV2TtI2l7EtuO40QsHANHso
PGtZhESQd3yKAM9uiBT33twX31rxvCkKGy980h1EaZM/kYXSxA+d42zvUYZQ8u2ln67J/EXb8+p+
zVs85w+v0SzVAszlLrbqWB05yzuAM8hhH6Ej4/uNJwYXQ7CJQ/JEtlSZOATPXWAfVbM6OaSz4Hbx
OgUgWbINy82RhsNKmJmjxdJlzjb7vNJqADIUT9Znls0f44Q9McwVOJo/nFjrVFowrY19SDMtU5xq
myFUL6ceDwMvP6WKmsq8L2po8fCH2CmTQRa3U+5ffarldModRBzvfOLVBQqUxeNteyFoKNVXncqg
SIeQl0UBmDlLtrYQtoezBo3sxcWw28w08KzSHhLfH0VSPOmgmhukOiznwcnihEbWP6FiHtyA1kWa
BF2JNcDYumDNr1fwR8NivaMN0UNJdYUFA5M8HAGahc7NWHGcsq9qks0rRjOoeBjAUc1cCsER+96c
1GNPXGKPq/tE6By+teb6+EuTque7KM+2foZB5N08mnI0zCXMxoCizd8dRAvqvBjDYsf+GEKVpnrc
w07pfFMQMw7ewqvXFEPnuNmE/gIE+uop3IIaX+hUsO9vE98sCFuaIZuy1O5aW0UV7FBXBeZb33z0
EQYGgWjMcdTdJmOsvxwlgkLsvPVpBBlZVMnYwnfTSHJtaDlpBycKuhfAeSti1L+hAP5P7bj1Bz4M
/rdMoSq4UmuEwgNZu8TZ9m6L777O2mfPYqcJ4fBRdOHzzmBfG+5SysPjQO/Ce+BXFV/Nzar4rzDH
I1LxY9ZtETK04vUYQbWqtZuHfKXBcPPk15KGxDGdscbwmGxMpxIkkjBWDtWYeZ/7VwDtPGJ52TGx
y8ZVkhpC3yrg/V/mGt4rbFl69vVfYRzIEC06MkjCcNnQ12yLttY7l+XLu1ObBN5+EUQwl+75Tk/M
0lzp+ylndnYct6PTUf3i+ty/O2VvbM4jphhTJUX4LPmlST97WllFnm/oi4NXGaoQYYhU5FJm+GnV
oF/Cbzii84E6+JO8/X0pazY697UPJT+vIJTSVmLUc/1AG6B3TpwrrEGm1JXTusKioefuMtI2hCdE
0L1b0xghmgo5DQ5yhHFo74L4oGeRa3Sb+5nJWNf4jrOyNUFDSJnzy2Bj+h9AaHTzmQZTI0M8WXlW
lHF2jqcHhWR6X6Qpvb2mu0S+MfmyTOkqxzRa8Adm6OlVM1ajm8IXDLliWQHcIAmYsrM+s6hRqP0e
Py/tQ9s0/KL7g6MQpng27L/kYtj9n9YR0jzZ/A9k189LDexTQzIHVGCPcFtPVafXBreEVnkJsmXr
0PJpuYiFY9vxbqDuRQoohXly3z3cTAGotn8cb1iyXrxSLiNcDDnkAEgobn9DGmo0MUo1tMQgzhe3
7yC+7TLHCXq6DhwZJLp5ooOGUFOHbXpcwfjpLATwdAKZSqovZ6vvvIG6Y62BLo/zfiG2QZHCvZvi
vFzs+AKkt1AZ6CTP//v66Q6q++N0tjyORWga4VVKp89wLw6EwGuI4WZ7LcZOWVgPU2idUoUrIa5X
TGuRveqAhDDX83Z6ZjI7yfNDoIuic8CLddbFXBN+kk4yiMNn+qIWkRnjvWIWr9eN04rUCS7mzh39
NJxJjPMNUHgwYis77qkKE2+4EEKcJiises7Z9p4zc9dr6JxId3G+fOOjAfon8LdCz7GwjN0GC9AH
j8BePt9ee+8u6W6FScspC4ct+fzvv8T0FP21ZfAVBDyulsrWx+dhaolEivrriRBEZBuEtcXJReP+
efjo9bNV2JPcYq65PyHCCrYQMjqDzlwvlNdw1b49BvpEhLC2FA3lTh+9w+o7qoENUTGHSqyrV+2h
ha3epOSxufmuGTC1ZTz/HLnWWl5vAE86nodSHEJkW6dZYsem+FePFd1OxLxzQzvmQqlVFLPj9LFU
LrWSkupyE3mcTR2VV2Goj/ViZmIjiauZB7uSW0h4ar6W513sGDUbkyVCw2h1fSamJ5ZtcJoyLz+6
7s0FisebjHqKtTw8TpohvIsbisCvK3korkvcTfglTxNtSEEVtQzI1D9nXaQVmZIdxaM3Glg1F018
uihe7C3AF6gZhBh4gsTF+gbTttuAvotMD69ZTmScb2T9Nwt1293NRISayX/ZA5sLh3zKXT9or3eJ
R83bI9LhDkM5bPHJZAwH+y2bqQASmdG4QUPA2RlvrvF42XPsM1nkeTkT1pDkMaDNNgLpe2rwBBxl
xlfFX5T61vM4IkzowKers4heph0DgkZ8056V0pG/SlshOELRUJsILLWa+NWT/1KDwyMYhspUVOkq
4jioFfJx2kWKFj6R4UC1oouFTydQNfPxo82cbvAABr/cYDcwof8Tqk1E93aepU1yYZOIdU/V4jRh
WIe2SyWXgbkqUh1gjE8JrfWVlS1xPrjnk0zRMXM38uCIkOGYQCsGwMh7sSff6vfrvxGMXuvbllV1
sZyscW6IcvP629R8f+Br8TzmFWa1FMxP3OfO3c+4j+/PLseOIu5DGLfSciuj51MaLXzMyl7MakZL
bEuHPyscbZmLW9ZEGuTjOBtLXx3lbhid0hdVS3/YzQyXXVNFy5KMJMYfjcUzmUO5eC7c+GS9ot+P
UEJRrjv12cQQIJSVHL6HkeLM8r7wXEpHHy3srQ6grURf0xJComcMQbY4+gcNuPbvdoofSTTLDdm1
qS2cy25hMlZ/0Okoqh8Cssm8p6w2mGWkf0cD2b9Rq7RS2jGkiDhQcMEPcOaC/ZDe+0oiXn4VEqG6
BsBAcShHZy+Ybnkk3NhYJL5fRdgaWNX60pP9sSq5OdV3eZwZK2wlp2oXj7p4C5dZYn8LVQmBZKwQ
pAbUGttgr01+iRbeb22NAmcFKX+zvttP8KMfRpqi+L8t7V96OQjRHNdXg/+bNWY54Qs1TQoQApXi
OunGrt76zirTvd/vXDW3sEWZ0OnemopQ8C1YGrRS8tcDkm4nCXXZTKUsqXlbtDuJuy5j8xaqUp7Z
gP5ckLhIuveQI1Cxzo3Xu4vHc3EBce9QYhSo2z4nwX7IyjTrULTXtqkbbDsplGCa4rTR8s3v/gVN
7T4Ykz9zwzBwGzmby2k8m47+R41bAAgihMwRIJ7zeQDD9Og8H4sjiEsdYOveu1WNona4JtxLyuAv
WeQqeuBRlk0L4jveRe+BOp0ztUGNbY7+yZkWTeC6W15wlTkJ8HOYDWZvl4d82XjdXBsspFTSRic2
e+WLsMBfr+KqvLfROrnj5vFEWx5fOLZGMzJy9igYoQM5ybtmPCaWO9on8lhIoVtud7axgj6t2jOI
7j3o+54IpwNvdm6ZdEJ0uSIVWSJZh55gFY3wtVbbMTrNwsIJ4Bby6HnO/epJxSJBtauWXgZTbPTH
2VF+IxFsALiC+NR7OHwI5If64YVxBEDgV+csfSCv/pZ+sVboTZ3/kSCI/EnKIe7XCrS9e2ennFzS
NAQFh1PrRJrMI7NWxCIrAL57gOvJQiujv0JOW+XoA8uUHbuZ8uoWlTIH3Xh5hUsi1s/dOb2c1HG4
ABSzIGYVNH5JqesNn5CBS6+U/3IAq7OqE5oHQIagqx1/kqYs0irDAwpUYs36YmG5KmgAFSzthusa
uXMzpCjIwIAYb+qjXufE4iUeRU8cS7q3BlUis9jgYuWDQ2ie5oO7aL6GQFTnz9TTHm64vbKOaVYK
eIMI6m2zsLyYOAJqdf8RFT6Kvtn4bdeTtuyR16hIugL/fMwVz/OoHsT+p0i6c4vfHp3dHM81I6/o
ptcCWfms9ziWBdjNSmkXI9CgnJiuzwYPsvhIdQ3eiGk+XwIZD7tpT86ARR6UQMlCSINDBGkKc5JB
W96CJCAqPLGWc5HRNa/gpKeuOE4zxswI2DeMYFhi4+EKUGzL0fK5R4m5yrqtMKu7Ows3Q+a4QddS
CNdk9jLrx3/eGnyEmijD7RNgToDi5mCyvsneejdaufYjSnpBkvF9QgDzeqQUFczBRHtQ8nTVj0wP
wqLpuWMwZV5cUwsqRWp3cqU3tOYLYItUph1xI5enyhMAIA6F6tk2HitfT9pr8Dr0ZfK1UdQC1QOO
LyjxgAthUcCEFCwjPVMsz96RSLe+2GQYNdCJJ6OQ8NPa/5wMGa4KN9O26bECjAqIcs8l8+vSu2x1
V04+QubmcfbbeCOLgpPM73C8YCIzjUBlp4qQ0fNQJXgr5xgLgoG9nnauj6FZfSTGTHsPJdvKIgsD
nGZbOhD7PeNG7zIKjTLetqvGtfo76H+M74YwNteq2Qjc8Eus5DnRluH+gqDeKUTI2kpmG6Byw6Ye
oloX+VBWgWam9Zyrl/A0w3f61cPVhPxlp8kZi+XBQQkNAWPW+hqfg87WqBBStY/qBZGOFHPULUPm
xbuTSH5ce8Fl76mguKUxs/He1UzQq1JVntvlAk1/M0R1ynfyyyV5/Ip2PBk1gAJt40PcbgujES4W
sKkEKbMDjLalV8O1c5Ukh+CYrVaDagA73wJP9GdtQoXeHTNa1i39D/w4riQMgL/H1Fnl9sWddF89
JWB4zaIcXVWGJqzT53KQDHldb/3gN0pBbW5aiH/Bjeuvvc9/D4VjGG7luiu4p2QDacINM7gozlo6
P78rtyhXbhewuAzT2UWeb4p8TqPY4cBsyzDiaSKxKFlZezqatsGhOsquSwbwOw4dW3ORTsY5yvGd
o52mI/agfjeY+LCqkTRVncEg50pJJg0vXhpLIqa3dQW0AxjVum8ZY2ukkyu6F7FZYV17brrB4+rC
Jm9h2gADli4zAlkvTN92D5tWT+msuxSeEdBdIrSaAukHBWjow36c8MAYAPheCNq1/GXaJaMMAV+T
1OB53XeQ7rHl4nP4FJtIp49PbA7bi9/07ZQ5tqHPX2Om3sk14smukLyKffcy/CBguGlFDbV/3/iY
Tv2AIElSmmmkrU6etRhXhd9psEkbUUMypcq9uc/Mz2Lycwf+bSIsD9sLaTpLfPKQxI6p1uJQFb+N
y27UT+0T1M7tPfIqGorcm1zmpE7+jIhqrcp1RulcSGnSwDcQwmVGvtP8Unq1F98NYF8oM3+gs3dh
zKyvvFazqUTEjRCOg6c9gpBhjaZBvJCx3Kogq9NkZ0snZyiHe8aYAc4SZjnRPFTGa9KCJr/170O3
r+MoaplZuC/z/cYwJJB0OtIiQRyaLYPq3+tfJIGY/YXBS5AXp4OCc6L4W7aWf06KMVbuHrBlz4i6
tf++A06/LIkxs1dHKFgt8yNyicvwErc0xhXI6ocyVgEML2lEg5wqzX5PIl76oRtUCHhwjTKzHgHs
hbhvqogu9ffmsmJ9tvwc3FfFfi/jsI6AIv1nz/vYyKCccrUcmKV58QYLWwYiX8RYNg+53D+DuQ+8
3E45HHXxF7QTYwFwrSdsnX8n1arAMIsGEHnQ6FsWDfwRNBb+CklCP+R+ztTHcw0fhtuuBGvOSaSH
LuhVXlbaQTGlsrcGUX18kmdr5ZpbTVI1BE/FGloHIK98mGQx50X1frqP7O6lWYMSEfxpswxXKAhC
GMF9FZTjxnJqa2pIFesOhQUCSOgNLrgtAvYVX/HTpVjDIwXoCOPeZ3w7iMlSSV7mrLFECO4E88AQ
Pc8kBhgLRIZdIZ/Nn6ISpv5Ae3hWmS8I/TVk9QEBphOd58H5hYAwS96I+/P/u/cY3YFkFuBjV8Mp
eqRXNO8UXLf68rRd108k94DQnB1Ird7j4NElY9ILN/U2Cj/mubwR0vYhcxlNpH5xrEfG/Ai8b5M/
mg7AD7OCjVPE0bUIUjWFzznsu0edGt77JIvaHjOLqRc7flz0jk8qisOcFush0CjePzTiBLdShNyC
CPsL0aurZy190eHkXyafUHUc4+GmaPG+tAKAT815P+YXQ64OJZY7fFTqO5U+szPAlYRxtarbmgbX
nuY/O+mu+fK62acDQ/E7lH7fCqy+fQSXroOhz/h5JeZdcJYwKWnWQhBIyPU5y/gaRBIfaOBUUEw9
fxeLbcZXymYzHbGPpAElvtnL5txjchzqPe1iBLTfbmHgj/q70ll8iQqwCcfKvlCVcmkmIMMpxV8k
SUvggyY8uLqwxFSvsuja/tk79AmcPWgZL8XWtW+aKWcq3vu1BDARYWc6tIUG8PuIgwU0K6eNc40a
xryWDjqkg6kvnPgPLnXqRAsoChgXILAYjwAqIhHf2duScvTNNmN+gRWvXy//aUQ+eq7IfPIgScKG
zVyGzKDyiljPzAnIo8AykGV70+Egj/MBvVAVp/b6pEIIOkrvciEtHdqfhfnJwgD7KK4UZAHkyEe7
4A9TJ83dN4m8uy+g+9o0Lwr78bmyvEU2yjqBUldFsFo1mHHQid0cs11QbG0e6j8jfOwKf2U9zBmG
Jj2MVclRG3Ghu7k6jCoK+AfZ62/fPnZ5lhkcvR4Aa6F/3Lz4AjbqRmafEJ0Hf/Wvd8z+lBTLS/C+
MuVSwocr01PYNkipUxeJZv41aXPFPlmZ5nemv2kxkbwqxDULFiaeVroD+33eZ3cVsW12NzXYpRXl
UoCe7Zk7xCFZFoJzCuVQEGwf5lcDpGoGdOp0tYw+aAkHDvW+W639VU708MpMlm0ypGY2dxqOKUU0
9mGehGZXb+XFC6xptuk/1obhCA+BYyPKDGS29I+7ja/DZJJFBGrsnu7A29F51+SlxnB/H26JZ7En
oEVQop11LJ37wMLPDEZCRL1125AUtwsx2oKoKtQpkAjRGzeVoboAESveAjQn+4/fKn+AnynKzNr4
uYXxNi7BJO6nBJhujzI+7M0qFuTcr/nD1wo5mKU+p2OHhcN8L65Id2OujRfehAWC9tNO0QR6t46p
oNY3fHCeLsSQhdO9upOu4cQK0myirfXP89Kokp9pMlP9YZ0uEHvvxqwu3yzo7vlA0UgWItDIGJg+
5OKDv5GAv/ej7H6yT61eYbi3B+TXr+UERBibttgkZVL4LTtsrmtN6i4XEfSsTX2SwG/hnP5fxx9P
l28a8Eoqfp2orzjoEJPxOPnk7xH/NFwLhS1RnZdA9hIQIlZ7+cmoA/jeh6Z7G9IPiJBPcN7IuX5h
G54MwWUzm0vSPdV/EYrRNK15DSUezNJE+33By4NZ9MukcnKm56pCa6pKyjAPF9YQtxor55yh3NJM
dULvX8wE6Z424v2oYbWfAeDzyIt5hwZx8vARwY1uf9ePHD835V6S2JIKGKKiWwulIsUHbWoEkiYP
VQXC5iJlV9jtzfMqfIWdov4cIW4VihiyuUr56MF6tFrE/iFYinP20AvvHfwxuIFbb7xTlkjGbEOm
9wYT8pgswFB0AaJ3X1nuvMkcYPTMMKGhtabkpL9E+lhaGe+7wiLv7AsxsTgIPwI9Z7fXQfTvyugO
l0xLDFaLg14yYGmPQl3Icq/yO8UGqs6fnTusiNlB6Y9tdpdCrSVjFE8EaggmFLnyqwRlMm43lYjt
K+HneBB8hNQKUNr2//T6FKe9y7J2wyiav8b98t35FZCTBW4qjqOE1LPNcjnv0xxVhE3AB6tAuV3d
jfaZEoLVLHz6+te54D/U6E5TRJoOmec8icAJxW/pOm9tzmN63GmjheU2yfmlGNOR3ApKYmRzvl+E
/GaK7at8UKvKwcC3vD9alRd0YRpVHRAHKTiz4cFNv0plYsMwzc+jIaTLVS+qZ3wqqKd0lqPmEAK2
iCwvJUA3CkjQWciOV43vyXcrfIy9Ezm8BcjpvyreUjMU4zaRtpdFuENuvMT2sE2hK3lzfOQepchP
oyirDFavcprIgHAnm745KugTD5ckWT0jDJCDNct6B6PFl3zEk8e8McmOx+ReqFOnSfwI3XJgGHDa
CKZYZTuNgcTLYzDSGCQMA9uv0ONOejnnLMnh0Ky0EC0bsUrYtKgHBoFl1Jh6m6WAKGI4RDVugaRd
aX5QHgcC9vZPTXHh0QYMiRhKyFnC4qfupfgGCDqL3b0mMg39ctcB/iroo+Hulw5aGWMwojgIM/wu
Djds7nRKcT+82+NN0hjpg7zeYe8MclC+HEpr/ubxMK/+8vIDkzKgfI5LT9zsa14o+PGIa8xLJLK0
iKJyM2VaXIpABAN7m3C9Tp4wgqE3gUZ/9HXrcH7YsnMv3InvC2bYl18XMuWEBfj+djEe00Il6cgu
J4bjBN6E+ScwuULlfhHAR/rDKZwWqF3xbnJp9dm9dhWMbSs0fjnfAj/S9SeCA4pxqPqXPqFt0T7c
ADXVehFscSdCpVQJEtvEqj9ZLhw9iEeKqbfapRNSZZaraBZC8Aq8ryRgbfcgJGnnIBxMZ0CcUKFS
sOpfjTmE9jUAs5LHZ7EvSVNlse35Ia9JJ80Zq1LBWhnEbIQGs1GOOIufC6AL6xwseelyZYqSdAGI
o96DoCAQ253uPqkHzB1hm/iynegOBAZJ/x9+TWJ2XEXdlbIoH5Isu6wjDlSHZnKZL/jnuFCGEc92
Cz5O6MrJLz0Nl/o/yl1GBrfRfAYQbKCpBpLcSl7oroCam2MPPpA0MYBeRaEY5aHvYPGV9nsEzOG8
biaASFqmhplesOI72cdypxr84g1pZMyKD4fgV1pg2N3KBnfbuCMmsgo9bazV9fwQZerDkMqwSSQs
2/qYIP0jxm2a7MWod50WfNywWyjn8FeAaGwcGEBGD4e+nz1ucHUaoBVgvyhYy08hXUMlBKrxxrI2
771N/r6qjYwmcGV7Jz9V5aEor8AX9KbMXoeGaUL0j/3Gz0OXzLD2OKTJT1Wdhccp7GZMRXl7WkB9
Q4nKgnoHxvZ6p2v5knEBst/TGvw2Qxl4jXUhfoJyceTjCbnlzWavYLgXWIIb3gtwgY+5bGmn/kEB
8S7gzKUc/oN5mgjCzCqocQgcnhVRM0CSpDL42iwKO2FLwpnM29mvHpl2JYlW7e6O0jswR9vqCDYv
TsAvTPc8nj4NlZK3vDPSQDBZbrvgHkG2Hlb9RnOSlcC0duFIeqQmYe7MA8j9EWtS5ievTm/od/A7
5jHqgGeM2+Ie2L571x4TmUw4GrJPdd+ytW3agd3HYk4rzk3g38HYn6UIXLH/P82TrtFZ/4LWZUle
LdOqKLKTCS4brQjoRhGdXV6hs+c51sXjBVhSTTDC3WvDDzUDlTifBVZibiGn+qtBCcLxmoFE/zC5
qctJ0IWiDQrZr7CqilrmHYioUxPfAA92114Jzp+G/uD7rUHiRP5fjXu8MRNVRqwaUJzFw8XI4h8S
ANSrMnpBqfStiwPIcUJ09GKjcvV+3Ax45P1gfXR4LtNw7o+7zdTIrixFll6bQcNIyIStkZn6ulZ0
aFoqU5qyApuz8Tcd04Jv0bGPe/TzcGBGgo5/XUfNVcNaIBZRj+mFIE1fkdsgCvXpRsBVyfwFtrh8
AK72bOjKJgR4/RRZc7kIyThmLsrH2yCaFPBZsKqLAgLFexPe+rGJ5KuLefxLTbhPMMmDCoYwQFRQ
7G5ZPEOJ6s+CHZemXlB1JmkesEd/8dmmK4qq0gZV84cTofPgGprd2YqsBf9bQGt5PZ/05/h6n1fB
PYl3GNWVV+mBtktvMnh05g9DgaBBlzhLZAJ6Kj1FDLBT8RcApsC7vnDslKYG3SXVvAifk8ECeQJ0
XwHTIMAC+w88rufiUabV3CTLG+tJ95kQOjJ9fbwiTdvCISG56vJP7Elke+1uw54uuixJuk1diKXE
vAbK41QlWwOJzp8LkH4d9Y00C8Zs0j6x3+WMqmwXo6zrlwd5KC9vfGZHBMwaQEvRUH5WnpuOTFd/
0d7p/HN8AZCf0UaKzb7ZSnx7rYu+Si2VJfF583bFv/wz7W30qS+v2GIyRtiRLrlY08fU2N/QJ7RB
AODSpcZ0XKrPBqNVBQOgSPJFw++eQz91nhiMEQL/P+7gODiNyKu6Y9rsvAvgb7glLzoGQ2zSddL+
kLPplDw+D+Ywqinj9PkBqY3mGdMEsbLDJvtqByHuNfa6/FihRTc7AqgnUxqLcW0KGER2tBijJWPz
vca4sBoTdivERMoue6AZvqXg3lU2DEoNHaT0PjP4VZnMqOXPItoRAZxYbfv5ouLbZROtcvUhIk04
GhOVefxQ7PfB3hWyRay8k5OUI7OjpFc/WgQEfn/XbuRDFjjxq1WM9pxN2Vy5PiWyV6Zt7Pre6jcV
fOa7KuADt0wL13AvFmxz6/bGsAjaZkf/IuH6SaUkQT1r1cJVLRmbRKXG2KUCrjUbUayLsi6PlZJK
M18V6Ht9JRbATap95ToxtOA5P2VYChN687wrm4WAfzI8wQrhi3NSN0y0m6mAnQ/2oZKeDsgfw9G8
Q3yNbhkHhpjrEIE0AmBzBzJDLh9Vm5++AkI/B8fuzLv4K/FnD2nOo8vSXUtR+PqFy6aizjLeocb9
s+oCmXevVuqsPb3a2ul7sFdWHJKQIOIDXAgtb4ZezvuIMr07/AsbMT/u9d3AXoOuwP97OeBcf4+2
Ck7hOmgDzdUPlzsik2cwixze51KlXv5vm/25RXbJ+HN+zo9AeSVmVABfrL7GQ1BqrV5wWVjTeWyJ
I7amvLk+QArotYvm3j/AhnmMzW2NDeaXll00OG5vnuR5TBG4ftYi4uCUu5oR7u/Wgm93i2JuDmM3
Jm9gDkWqvK8YJI3xrZUeIAEamuyHl2pmtc7rKPU59EqhhCdxVJJtbbtbUYy0Fe6SRzsHXz520ADn
qaZ1h6WeGeaei8/yLlcScNw9MuvBsXbYRHrAO2ACvUm50TpUwolzrkShyZMtCHTyBy15ACplpSxG
F+6QMRRLsPtDkK1WE+K6KRlagsJxpi4bTwh5AO3qVEW6RtS8sGFo94jfZzNiiNJETzOgNa90t882
QUTpcAXZP/Q44aKscaeambUlCXLKniD6hh/lKFFFxtql+YhwnSrRZptiqctAZKMuGP0RxAu6XG68
ZpFzdVPQWGkD0iKB2VsvGAEG6oK+G1rAL47tUcKQfWtYb8c9Palf77wph6zYX4qgxvt9vpW5zEqx
1qOmLivdpjQB5HQdGtNtPyzDuHTTkf7khYSqHxih6TedgdxLAZC4qscT1W/6Jhn2kjKp/5FnRfqh
IGCgyfMrWUBZv6KYNX3jR0qpy7ULiNOYNbDQgSSYBVYY8hOmV6OqHPbpXr17aIFQHE0nsyF78RmM
LnJ6X+l7Xg8nfDH0Gx8Zl5LvUocZHQcdRRpWgX4Q+TB76d5VucLLx309SndefWvcnUki1Z7fDBFb
r2qmEV7aJrJNysquisUgV7siKnr/wHtL4vdEX047rcOCgLhLah6+kMCFWzwl36CNZ2AWeAFt5gAY
xLb1zYb+o8pQUBdOP3h8qDWNVOMzHRP+EHDs0LZUJaApkYQrkOqpk2h3A58en8rCWDJVrje27QQX
hlAMUkinxOIKLSWPqIoVxooSTJt6+r1GS6T44TCWhfQ+LT7o1VLHioaqXYjETHgMhTFNWF+dVrF+
4p0qzSazaouiWIQ3nApvhrjrGyvNN4+grN45SSSmYvwTtmz/FHtwV9gOIhvlgE1TTxu/wKtV3wvf
ze5+mnRa4Du97fy1gY3x0RaeGtCyytw4dOytfDFgfN3Ad/fSusMPYTDWw8gvXVZb76YGdoHEQxbY
XRsmKU6+z0e41H1rkXg7eb+4vey4RiPj7Mg5YfNEY6mUiVgfy/kvsc5GsXcvVA5SCYmi4PkjXFOJ
4Yr86RqBLHt5BjZXHIFvGW02S/KHhxraXcynGIAVxQhvqWigq+x0fau53Ig+I4zirdZubGdh44BK
K9OysyRk+ErZ4anTkjewZRsJZIQzIBZc58xd3EGMPEMFJRGrJCUV0WalIpLRrUOnkCSGNEGne/Oo
yKif+zYQ8Rl+ws0Oj8NkbTJmZ341G5EDC9T+HeVPdgfFhU8AugDdB+Vn/wk8cFKvJC9xInAIh832
SC76djdl1HSi5BNoWdii/c1BTp1ZsGWpzIWknGLbbsEMwxDixfjg9qR589ds5rRuP6pshQu/qbg/
Lp0D/45qDAAJtwSVNN5K+CMee/E3YgKAnDfgMZ0R4iRlUotHj0V7RLcNsGOHJIPIrpiz+S+6t5Cr
Fv4vbCrKoK/R4b+DgBffkp4EgFfVVkhpxV1MxfBDPBP0cuGfxJ0ddMcxzx/f/CEizpufy1Uv9lI3
Z7Bs1kTXRHuPOJwx5s1cz4y1xhZ8tibKf87MY3WOresN8Z+nr4uOTGO0hQcRU8vkEGBJ4xFPOtvm
jZ7n4PCTqUiJrJezn4zby/RGi8S27T+KIhKfBH7yXWlSE9aobupbx496fwPpYZhRNJ/QIimgjy4/
j+KocMwFQwbrDA+ClrmTo0eqKHVHDVQhNgYlebrxmMy0Wkl9OsdfIhAjvkpJOanNolbCP42Q2xhM
YO9a71nbLzoRWa/D2EOXv4wb4NGmzwaLPUvB8Fb7VOlM8l6nxWCxA5JAVXeHSee6BzzDqLQ0T1+X
6QFTtaAuhf8p2pI/iqGMJEEZrdz9ZQWkunKe1AnfVeuGQ56ew7sUV7jnsc1KZ6sKbCu7gwsinx8d
WHZhLn7EBFw/Pa4OVm2hD/wBwJebmbPqAyWCqmm5Rt4U7OaGsYzJasCyw+6t3KzL/liH8ANoiAH3
YdjRqeCbEvhJQ+OoX2zU5BE6UF56t9wyKd5V/tquXJutF4PZ1wMYPhMvoN77CTInkF4JJ+JG+M3w
w66J3JBpjrLQ5oPE1JJKUPDH5qSi6TFfZcKA8lT3kYVS1msi0+CrRihNPd32A6Vu/2tPR4Jv6tcR
TYBVM1GlguMpH7zpfncseo99MinkUn4OaK953FTDjD4LMwefuY4vZMwQMl3QcBQzUhBg6kX0n0oZ
nJ1rkAD3iYjcPw1MuRj8nDXud0+TkLuGhsjNGEv0h3f43mMrzuLTXIw6gTWYI2N6NOl8q7yDOBvW
QyUswYwulhKP62756xYzvIjoI5O6IjyCG2F34oAmKNCkacFQmOFEWgPEdCX/9trsgjU6Ayhwrfzw
ztYQvHN+EHC+bUFqGpN33nNSNXmFhv3BgQLlkYlV6w/H/CiGvennUfqu+/JAbXpRYYx3OQljtpJs
evJFwpfKI1cTk2CYRAXY/h8aqhQGJ9b/rWPgYOFVicJWa2ZdRR8scQoIm6uFqDbNGMG4zUxwlcOA
oMy5CsXMH3b/mTUsPwSWaMP/nG6NtbD6ZbNrBw5vcc7X9+yOXQragrBm6CqLsShGsuvzkyjtNyLu
y2PPwnrarQ6/ZG9TJ3hONK13CdsgmU0869XayZdyBlpTjAzCvPw41WlkEt8av1q6S6lKFUmTXA6j
6eTx5Pzw06UudyiM9Vhel4GvYzu6JNujmY8+0EfPQgKoGwMXMhJd3fehiHtgrCMVZZscTQIZt5iw
ciTdimzv7q1GOreM41tUKw1H8GwtglVnv8Vjt8c3d/Bndci7SPkEt0L0ES71FZ//yPyCpjZk21Qd
tHNB7IZfQ9dPU4IkNgFzE5xezkmQyaNdPEmfi5VhlmHda3TuC/rUBO1qXPxcDzcxR2zmPuJNPtVj
sGQFbAbfY2jcBf2tn7S5g7Dle/9q8IL8B+bypeJSCIqiC8uz027uKLJixNwrOnzUHaV/GWk0StO6
QGDRWXLdIHQp8AV6PdYFyIT5OtYIqwKQIL1e92bfpMX7K1myAIbVGEo7smBM/SV5xASOkW7e0SrJ
NvN5hIZ/j/dni5NQMsAGrXgLjnONf1RfXd35TRLYORS33SgzKrAddKuf0WLf2zeplKHBvOxRo4L+
ZIqXtmV0uzUt4hmyFKiMzSM+eQEVVea/YmGA0575sUGYo1C8niYY6zE1t4+SWo7/oeEjALevtcuA
fp5/nCA0UiTR8MD8TsNHwraSsxg2MmMbVMLluSxUHW2uD6pRoxB5FAONPvO27SmvPiQl2OpXBSSg
3QVXojxEfZIHCZYHd9G5Dvbd1vagdtST1UxDNFW6ZE+PKksuon2CxShgd4P95Gjjq1XYRhtz+GAd
G3fpQVGPaQIuXOMjrzQG1I3FEZn8HpzRAHfMN1mvbbujKgThysrXgMkbzAy0AevXgiZYPZbIz0B4
Yg4r1yZnx6ai7B0v1b66iCKWz7dr8q+E5aEe7srZBXS720v50UrH6rkc7S9St7xnmqN0QNIfFrvJ
3vNqFaeOiq+aBLexAFA+HZvthf+NhSmLGDHdHbLVVFexGntgwbaQ3UypB18k5erCJMl/RmqiYpgo
2ySe0otzECz6t72O05U08goW1s1ylaUwCep192twZ+EvBT2m6DApAxmtQTzc+o2hxpn4zELLFheR
xEfcY4afzufaoHbQkG9cTAWauD6+frSOExIOUEMA/7/xlOwxnC3B3IXut1LgIUFsroSFz2fEJyhF
84Ugyhtwxwvi2zXzeQ1FmjbgqUe062rYrN6j5m17r9HRnuCevK9h/3AnHP91aGVgh98ro6CSPbxb
LsqiboRMilVbRuPretjOQ+xBhNEeA17Wt03N+/4ORYxOC2mNZmeTwlIQ3F1LkbZQwwDYqgLLMhsb
SyS+odZj53IVtAevgoYVy7jxBvs1MCSm5N1FTAMGjsExMckZwnVKBT8HxPqJeLcf9dbguqGigMDK
WZFckoAC3AMxreyvx0A1+sDh1Wfdq3t7f9GGHHAFdhHB/Zq9uJbHc2Z8WRPdZBHz0UzzX/fxY26x
a5omQuPJIh1pPCaO8RhGQ/xfcOITBcP5/gX6Lp0jkbUgQU0hJ3jmy/oIrYEs1BCpk0Qe6mNzK53I
7zGDb8XOptyO08581sgmL+mXASRpNUwmYoG5q20JU8be2n5E7qk/tKtuKcMlCgNHQfdvA3qwFJ/z
Fu8sa4v/BSSKtkmNinoicskAf3fPUxttMlInvGCmSCRhJQra76ln80+bzV9IZCFOb3CEeu1ggwyJ
PuQ/VqEEBYS950BQkCwYUmPLdP/aMoREmlWd/UpntyYHw2pOSqg3/OGYCSqum8Q/M4qqmDwNi36r
rYBdIqEDgNGKL75EQ0Pllkr1JplFrTRJoZDQme/26tKSrqkV6qesFOz+OP7bEe6Q2j+J4UMOEpUE
CYmFco01y7MZxrmSwXev2z80LuXB8IGIWErza1+uPakFFf6+CFh8HbKBiuRDUf0BjG+pNZe/4rva
4zTt6ktvOrdawmzaT0eMmJCDsgFNTvGpXxG5z6HZqYKe4g8D4BVMc4x+e8X4p+g3NHsQKjUbjRKW
I29qeXqWZSeW5gTQmyxKLzf11QkO+4aocxVYNJM+1mtSxxIYU062/AnBSMZ70j+Sd2LrxVjjKPhV
Ywz0oPxeKPDqo+Gim+fDBKbwQ0asQN+5JYtXctcm5Ixoe+ZiQoBRsYMyeMHwIbfCtgu05SjyDpth
Fxu8836kGBykdLYn8YYNdauJFxcKXaJAaLlChqSRNch/nkz3H7EmTgaS9fGHNFIXjDvh7YVWk5p6
h8LvGLZBswhPpUNK1GFJneF0O7REyNV07HtcFUoSuRCuFU78U7PE318jIkrzuzIA9fC98Rlrq5F4
LnBf316dllvBDYoHwg6RLEOyPNKYtQPLYbRVLVt2CvLXJJJKs++9FXjwN8kLYP3YuMs3XzYcy/Ao
fbXx32VXipqLmM3bDX8MFvLBpD68OMT4li+YM8JFf8iO2kUKQOctJ1jv3ScHzB6Zbuy0W6jgkvZc
4KDJdLWjIVDGRXk/HlSybE7ZNDr32s1B772mgq+//Mkyv5d2SV9XJiuBxkez4+vM1JDCSV3ovBYT
dLhKManqub4B1fmdDHxYbFGXn4RF0/GUgWk1TOk9vWaoWKz9v+59tTHQ5psHoH7CIjcod7CpmDzH
Mrx/Zz4P/ZfuY834WJOMcMQx8yJ1FjFk7/4jppMBeE3HPXRXY6fT8Ghttt+4J7+1v+jp4C1k9vrt
c2cV+PyFyozQVtK8LFfxd4SqiNSOtOlT8rk7URHhBsK0yayKUfjeyOLKIhpnE2VWIBwdhYqCuCVo
9QAy32Y87M6Df+EpbQYDwZli7rMU4q8DsJJ1DNjTms5vZ9o5wG6kpAmxfDKVaQiEv24YwA2+DFR0
XqsEVNmZK7lh8IBzFboMA2DQFX69m3pTkIp1rd5s/dH6GL8DBLAkQytdQTQ3mJIZP11ecg+pTErk
tx7hHaIZjL5JJmLMPtZ/qlEYYxfd1kLUas4ORF3b3RZkLTcfsYKZHs8CwWj9r4yMMyhkBk6jBnR0
mKty/NWHRAcj1EKaDdKtvlGGzhPmO67f/yHUC/ofw+6NVZOoJxnB/sVqoHAT9Iu+WoT/jxNcbowP
HZlfHgHaB+m0lWgOO7A3FcVzL6zVZzLD9s0S1GiyNDV3vwzAczeYx6v7StL5gjbfw1KVTGFS7q2t
ormohDmAOc9twMhKIEnWgCDRk84gM3/Q96vjPSQk11ki7VlTKV/t6o3GHabBu3PhhJ/IXEp6Adll
PL+ydRTF4u3uJ73pIArQ9aM9YLgK6APcw94k7RPRiZPuIKFHf3Z+8prjKJhgbp2sJGbMjK7xak7z
R12LD/a4rc3aIBvnTEWbNnu0BE0tybBRKgxj6x8+eOJLz0lqwnSQslTxpuHvczWpp/Sb0q+mRVAr
fsmHcgl3LPhot6HD52amF6ytl61Gj0NV5NqNbAoTivpfHcRV/yq5tLcBdcStnVfQ+Nfirv3RsoMS
Xw7m6oBxvelqF6cQTLQpnn3dbivPFeyfOszDCSdzrSoo704dMGDmfh/X2a2+TS+lKUdYyyImBsED
LYjrQeBFmC1+B+CVi56cgl1torCRBo7xXI24AhrzH7uBx2DmfowSfcWLN/qz/9p8iegEnSuw/uuc
zCF5fqRuYKekBVpQpScaizGN3u3c97OSO5w+u+tMT6Zqr4TktRN+y6lyFQYyd3Pe4C8g4LHqxE48
xEQYLXhn26SudyKr3i6Ii5AyCJZu5WByqXy3EmbNVfcn/EZ0gWAs8ZiIx0nAUOyZmNqgIqhw7CSt
GVkRXGYeYYzfA4B7THqGEopm01Qb9K8p7tUxz/cjvhcoaYCu7Fwv6KJOAY5QA8yU/G4E8Ndk/1OL
H+zroN9TPB3564hEIQsmWtDsT8ABF+JgY548Xi2/kSh1Fy2okA1amKw9VuyuL/mqX+ssliRS95TC
KV/VPOdGr9CqER070Rq52u/rHR0zTIUJrvd3av/jzMNtB0t4UOg12j2cwOqd4OjmW1S9YgL1b+TK
XcvNIBS+AX7UweTBGT8ApyIOvfaoNNpYt9Hhw02ZGBjomBgGKwSb2LqCIuBxBPtalD7lfgOjIINr
Kcl5cw1385J+irzt5UpHgJjVM+LxduJYTlj2UevU/wGFjvndkjd1krBqQFQqd/7gNtabI/IoDbE5
sdzdsluSlGxvt90LHXEOLOE4aMXeSYQMlYCbG4jSAxh/TKsq/HTag07mvayJkZsXMxXwLYzcwqFm
5sz2W/VnLrEXyNO+m2+uG1rNPD5saC08ynYfymhatI8gRxM8aFCuN/jNV6hP+hTPw2HY6uuwuzdG
QqNf5t1GpmLUJZGv3u1XkLUuzqupkbj3dGGNYZ4sh4VLNMeIaYTNoSJ9HnYLW+XQuGYxKXV0VXUy
bc7MOT6zryHHjIbBKBc4caSgsXAxcLIYWX729j+vpOBzVvVgYzCc7rq5FM0CjTo++qk9O3yIEN/a
9iJUtvRphW/kzJYER5osqNqYWJ3IfTEsRs0tuIcTh5v0wsAhu0sgnGACNihOPiZsZucbbzea3D+g
CRG6maQB6P439vIAno5Rt80dIDywRjjZEJ8Fbyx9meMN5yckFjOnNk+36ZIujA5eP1K2zLCjKUdz
iL0R4OyHzjPXgrur+4t4lEBAWujJZSXwbls+rwmYSZdEchET2VtaB3vms2yoym9GLlhaJzcv/kJ5
dEFlw2l2b9jz1iEW7rkP5idbD+nROBHoQNpZRcvmEkSY2H9Q+3KU9vIPYOL34ZElPaQiB1OO2Xql
eLZ9IubAhdty7tkS7vYX3G1Zl0XHG0Sl6/tozm4Zjenunv+/x4yro5SJIz4zXKMRoEAsy0K+C465
Q6Ni2nHcu9YloW0ekPHchGYsFzc3LBvUyE5M16jksRyxzoPuRhKEXto1JuxlrbYiLGvjAO8hkLNx
lvvSD+DdYdMFqT5MLP6UdB70FWz75q/XueaIGgMygZmNV7KMUWqXCl5wmcbbs2DvP+tXzOHStDh3
B/cy26v05aDKaVEHavifAZBdlfi8DH+fsu7ygzJPXUGXNwp7V9HZCulaQluc2vRP+P752g9lAV7w
O4jzNAsINmhuV8U3o49s+6Z1hxXRJHZLOLOcn1BJBdd2XZ4OGQDZ+XyceXZSXFKc8j/ccMsGtS3n
sW9hTeaWtg5n3Ax3wd1VmGSwYXWSyMjgc6zkk4LTf1zAA4FwMVFEKlWUKYEQJDqRo60gd/5LGhkH
t7S8GgQnP5qlAGLvnhkZZ6Ig/7BUNgMy2EXNigBSEvd4B+voyOrc8I+xc77gEtdpCKWAEAD0CATY
LQKYBVav1xfWxVh0TVqlMPIMnI0aQaTR9ObUl26fJ9qzlfcX1XwaUqliGmnPtue5gapueBES9rly
VmsbOsiFuRwVLIN+9fXkMxRFvFzn1fml7BdV0EDNSKL/IMj8EJCu5aPprv/D8PTSetmWLN+dJ8QA
eIiKYOm2YlLNiTUgu7x5rZThc6IFIAaAT7MxJa+ALE4oRHoHCeFMxMvUgmnEEIb9soG/mumuRbbx
GLrd+5yUPIuvp0oJrCYt6AetUDulfW+azzAypAPxOb+0gnAlaMl7p75jg+kq4d0fAXSgRTCnbkfC
RQiYfzBjihV5pGGGcDW3JwN2bFvZKQnARD8DR9xOvhkv4aG+AjJ43/Z94dOZ5WbTFhx05VNRvxM+
0TmvXPKtj3VkLTYoJdi+UJ+eHKhuSigcH3wDRPqu9rsD8ovvKw4Wt0m5XTQNkgWcefjDXu+++YfD
vRio/2RsEZVWStIikku7RXrLpLBIgLyuv7wEikLVel65MovHVfNMHE9K+0EcKlY1xpFBwjX2PBxM
uZ2XTP7JKxupMVkfYIX494dNkeTd/E/lZFuhUk/2sRiIU0gBSa1LbCoEdzK+CIEsTWde+j6biXIc
GqsS70bBB3I+7pY80eQz/o1SvK94bx+g1ocarVUICgI5b3NJ8H5KlzJtnC1Mrk+SsBDunZD/23xP
qC7uht/icVMsgPCy8qWLOrEXfwOvwIEbQY8X4pp8Kfd1QkG9ckD5g3vNlIEPuQbjY9dM5eyZr6iQ
HrsXGKSl4sGCIXFRu8jCDHqxn0RZ7FuSEDcOCyxfun+Y+bSHabd7rza8uAdSBQCXkKPnwegGhPg3
Ys33VTpQECuQMkuaq2AwiazKULey2SN1T/vfMDMipNE5JBtxKUwC4nWzP95fb7r2VHMDZbzxriHP
56Sq2dtbvV3u5BEFgpBw+ErfO8YQ3jXpdnOcJghk8p30ArYDPS9LA+Mnoy+N2DvASkhdND/KYCQt
5mdhe4/4Z7eCaRle1m+YGZpxB7v5MkcvIffOaqhpRrjMZP+PcKDhJpzTz0tb7Chy50NrG681sO92
x/SgWs8c26JZoL1KDHg+Bf+1ud79LuIpAWVZ7gC9J44ktw1o/JkHmywQ7idObrJoTVFFVC/KRAo+
9w+F2vdeyqDhacJsaAxYO1iBuT2EQwsxaa4Tcf8IB0r6fCpGZbASY+JXcpcItQhPsgdt/QWeNiBB
9XC0LXDTrDqPiLGWwJ3KfnIJJ7tkhN0Y4PsIv/l3HBTDS56EwRXANaV2BSNkw8QDg+YhQ7ffMUVD
dcaWoXodrmeM4jFGfa8PyoWIyWgIEz2iPSEvwSFfBKmtTlxeWCnj6kam4f4AVce6iPaXrUFdTDwf
Bxupx49WG4AFumLmf1DUJdCqZXqZsMpVfkiapvbGgr7yYyMZ3oA1ONvK5exYlkIhXbilWiGbmMMu
lA1aKXpo42AIdWEfFOX9hO7Q5WPdE6T81WtAhoPdiO7TjUzkkmX6dwngmIMCzrVW679pfePgXGaV
qw8uF2FUfbVRe1JlWt5pih0kPumwcregIX0CFMDo/AUnHV/NjuIzKDn0XMlWDsdlr11RZ5WmirgW
0FlMyTE/GqxWlcBdoVBskNkZPb7iMDwXkal7++IA5xZivYIgwqa9rQQHkLwQXoeU9sRz9lAwrRAz
4xtsBEUrChVs/UhrMUVXLbgl/G9XNSU+AolRlFf1LZNRzM+3USHYb2Sw/F29Ryk2oF5p2d/7k5tM
xtikcVhlG8Vq6FiUjUU+HhjvRRQS6zioCo+/hSvqLi2DI7iCe8TmX5BQpJriD5yff3fhc7F/LBcu
RDcDESZXnZHbVcDL/6MasPzCqsxujjLNb6Dk88jl28cbWUIs83+gkZOxiSDR3+VZVohGlWQOC6Ih
rh9SBbjrbA7m6uMnF7VPyALv3zGfvMQwHNHbkQrPGrhxg9SnM8icczYLK8crvflgwC0LtyVzkGGp
YXu2Tr69TmzH8DPdlkBdIEFtjblFch0BDdGTpQsOfTR4sTTFSNyJ6Qq3O3w+gJSj1TJUYOjca1uh
Ll1TKdF6cqiMmjiE3A5rXNYZrXPLji6cxI2EHrm3LzX4F1qSxsQZsOWt8vCzMCk8MNEo5pairwOt
bM/0DZW+mcrNeeXY+v9npJuBzipt76fOP2KDAiqg+yyWIRqZQrjWPKHmCHKo0pHC/zcqNm49UOzs
sQfbxzWNaDzbsJJ8By4ldNWZsKk2ogPWG81T8eDokU2HIMTCx45iFwiN+yJtYLqP797TmglqtBJO
boeFccB391qkojfXXjXCj3UYcDsa3jOdpvFSUNWnePwrxjvIW8VnwakWuLH5tY+vmjrLt8tbAFHR
IvxjNtDROYl+TE5uzrx1tAwf6KlmDOPjbx1s09/wtM0AGZIFgoyJCWvbwrC0HbsW5yvdO8Bodfxa
RDzT2cWSmqvYm1v5XFLuql3AoRV8BBHcktAgEoGeGJgq/SLaiFARLOFxwaAFsNJpcx++7DvlguJg
yCrJxy8KCXaQTrV5EylOnedXeer0BPSH4zK//AStbYMmRtfLXWLfI3TGjojz+jVjORDfwBCcv5bK
PvD+OJ9I6VgJ1Ou/EHvaYpJzoCN3PsqAoUQ0jKwmDm18geW/9s2CNOhtPesJtJr6jGjxibAfoA3P
9sWD5iGquH48PJAzZF/CiEjewnHBpYkp4nGro2oWML6H6gX8g4Ld+ouSw7LeZPQelpvb1Gq4q7cI
e6iLMqtlBlDWUKb7NOX4AuAqm8H5De1DangsnLZ9R6jCIa8gtwkaK1vTStRMO/sfLYNmOlNxYIh/
jmCVjgJVlzmW/YXhVQj5QS9qUwd5SHH9P6hEKRdEs06GokkSjIHgmY9MYLNnxiDe1sZ3RXOH0oby
Uv1V05yNZEpwqMS6rS46zy212rlFTIHFYh50oFwB5WnoVZ92NV+Zbp/LPmXJGO7vKpIMd8iuySEB
3NuVfNI/pHqD1oCZaONtVFWv+1wU1fEgyZOF4uG0MFnXDVN6vm6wkZCZ4wDidYkJorsbcmSFeX6Q
j3BclbgzjVBbALnzCeK/mSIZt3ObNjXDD0jSnrHD1kRh6CjwiWQMyh5Jd+UmwJoQqLMun8hIGTis
9OolvQ5e8lZJ6iyNXXfAmMCk/Td1H4drMTLUymQUJrcSB+TXPPiNk9MfXgqrHFmX3dtiyMiNdaQq
WZzq87QUZn+Ko6/oxv9JSCjwCGM2etptfhP9lWnt1R3hCK3UKZSM0BLQrZN3WjuimJkrufFDbFVn
2zlUPZ/lvz8vQdwcQ/bjXPD/R+BG6NxhISvxoL7haWNDgEHkv1avaXCDBgj57LTXSVkz/0UnVl2R
HsVt/i6L7yr9/sy7EbxGI8XgmpCo2f1XLW+hGhhoKJlrESltnszyXPbVud45cQ5p8UOXnGSehYPu
5fsfCWo62XSf95zuPS9x/IeWd7ZDr/Wqw/cdmYTAu2D7YWmuD3aLTMkcARNH5GRUcb0xe6TN1YDX
iY/sKfutF52Sq/B7yF7EkTwbXRt+w3lHM4lZFNZL5x51Hkzgx019dIucAcQujw9pzz9qNYpEtGQW
o2ms8v50CZ1/nvInYgjVzE484cO/KMvqIqueV5rqT+b2BHej8BhL0JcIlE+EK6I8yBt70pWmfCtw
CwOsR9A27GJOvOpG25y78lh2t26cBp6k2tw4a+yyW0+hwBIuFZEE1lM+h1aNQGVoqJk5L4+fOrdi
8b2uNy811DE6yo5s48aDqMJrTr15sY5UTQiEyAVC+dE2C4O48ef+Pw9dGZgV7y8YqHxqgtscoAQY
gCko2uXMj2X4jOQyWj2kwU5vWd6TcPswmW8pNl8mhv9HHuPqkSKUtB1T+Yn0MRdHtJ7eyl9mk6gn
zBzoBGKJjvw7zMtfSzphTQHnu9zdYb0RNEIWGA33rHqJnK52E9gDGCx2ULecV7plslDUfZE0EKGF
rxDcgQiwoH0tFlMVjgubyiOOdalK8mVpZGYOUAR2Jm+daBhMYuug/GdKPXCaqBGGLoC0y1lxSt4g
TmNQhPQ0En8ma4UgD9JND9x0tnOx/x4tAZ95Xn3mlQMMAeWp4U6ScEQGvClkPhEpNMhci1ANAw+s
t2RQAH3QnvskE09IODeeX+PWNrPlo7NlIZVDf4hbexGKLoEubTY4Ja2RQDzRkJ+a/ZV22FCw3EuT
i6KoFYYCwA4WiulfdCGmELNiBQvyX07YxRhwFDt2NjHkggUPzfFKihsuXtUVA929boQHN+sr/pRK
2CiZ2LFuA25fKhFq6YRcK7EwbkmIX2APMoEc/CACrrsMM13qdZkITfdkVhy/iT5eSTmszlFYdw1+
dfIiqTLaocca40HeRZVZH5B5pm5HKzT0a8NMc4xrP4Rg+jpXcdJrfKvYbq6Z0zVY8OiFKLCkbS+C
kIUfRZMMWNngpP88HYdYm7NNSNIpQ5DGIbbTATZWZCG85Qnxi7RcKh1Da/aJJO6fzPdtbEPBJplC
wQ5ZAc+1zwYdXCuwOxkmQJy6gyyr+R740rUjVFa4avQZhSI6kYRJtFUeorPkgPqQsjpjC07iEa4g
rjGuJ+GGF+ML+pVVB3dfudBX95IpVMMhIWnRMY5YnSbDkhk097lCB/ykmF83Dmyf1Duz+1coKpA0
BYClWI+hFoLAN5fQFNhc0fDlG3WiCGV7kKXqmxJxuj/0RgJJzFFcg2rP4Man0iXcRpdnoXOBf9XP
9UDylfQelF8gGHcYGWtaJI1LzLaYkphuzckafbP/7H3dfRYBUgH4jR5Gen4TjSPf3q8jNrdbjf7K
ucxgJhvf6G/GUYyJ1eWWWW2DHo+kcchIOWhF/SrckYt+D/u1OLgQ7Ej8XDD3CJQF475XLtjJDNog
7tIoK6nm7RP3uTcmvpoDEAQ80vFJ7cnUg+1X+1zfEu3UEagzgLug/oPi/6DUDZ3SdYT4MJYixbQQ
IBA1430diHLKK+WhKS2zNJZzCMdgxEz2JozIH6R7FgVyjcz9kEZzIVx3Svzu6mzJKOVPWu7FaEM2
L9DYXr6nTNkCWmUNbxFua2CbJ3A7Ck1mtRgWLaagpasmjJyvdeuIWeQ/ZRQZC9+BViWvQf/1qG2b
127KmyTOC89bdKWaLyE9RKn/6dffVSM41zC3xodsDbylaIfmVt9lf51SDMKZJ7oyN+w1JfDzsXV7
NiAaqiaupSTY0D5hg5Qok3QMTobYoE4gXpwx4CuagW2XwvcPfhR5LNeTdyBpoxCIJbvJuTfGxqWy
JFle7XZgN+q3sfVgSiSUQ9Sz+/QsdDej37R/5AuED0xfk0qBIJ2jlQXp0P9WCo1VgrE0a7uihVVn
6NU9AUs8ci4wdD6xkxif5fA0I6LCPN9wCApcKylN2OxtJzTq80PGlkcdx+v1MCWbKIU0K+QNFBRE
mxgycmeSH4EdJvMQfoFJoEEFRED90+wUBEbGf3VkxJU0djGhaj7rZXtjE/pXWCwCxqesv2VS6Z4d
4zhXUzA24KNTsFOXhWBA1+/zQ+UhOHSNOuOYb6bS7ixAA8vQ8kt6IQXP4ONVfADar2bMQKz5sGzK
2kY1O+DG7syaowscUXpGDLHjvuLWgzpufc7gMIhk9Dn6haRQR4F/SWpmDKWGNFCz2xWfLGCFWSiU
HO4hqbu7AJlEre8F8/Ub4k4MlNLe4iW/mHQzn2yHDMPsh9K+PRg0hDZ7FzoqfwAFU9+UxdOnDA6p
T+0edoa4q/8Oi2+vhGNYcgYbR3IwiHv08rU1D6XRB+ZhJv0sVxxM5fPjFXuSZOvGUp0AuOvYfsdu
K9JVFAxha2JfCCRlLAu30spF8HXAsnYm4bX325LkMfm89e2R892nGrxg7J8qGdykK1XHAsH2I2qF
8dcgp0KgIkuTiyrr7k5Hlc58HzA95xOJx8NhXR/0xqdbIGKvg9k0od52SaHxTzC2A1uXP0B/BtWP
czdn5nZO8WPdmpWnHAqmwmlrwSKhtYM8Jqw6jsjwyGxhIDMeRag347UMTxUja8Wr2zqsN99hRVmy
5CF+ObG3XHt1gblYH5rCxBN+D7UaGUW91nBDRY4zHqV161TMotxyNGkVkP210L4AAE+9MlqZ+yC6
czU3HR4QHlgHzuwtbZeiWbF2e/LrUm/dOLyQZiBcDeT9iSQrv3jG811jzAMXjGSZvHJb/59nRuSA
ytHciwV5254tvn8krxeF6GVd22tUWBNQxtT5pUTSN8Apy8uPmrEaoM2s1kmrJkTJja0p2TmGRNWU
3Y107cn3Sb5GlIGLzT6HgZ4YmH7yPD0+agi0jub541O1iZgqPytq2qW7bNaxCOFF5Fr5l0kbygny
r1AaqZllnBmE1Otv0cFwR9x04ewrEyFctX0XGamPDEaeo19Je1/MC+SOwKhY4s21kfaaalKeljLa
coYtl+5PGFSfGiJXzzfFcXzT1Ghrth/mcP5cBrSsoNSgWEp+0364wO+ouYqkcr3VXvvUezxt16Z5
ANgapUqfhT7fhqbgkOcRHU0v4GE3ASgsPjWA3w7fOIegys2+cqhlMaDZY7elvLMfqmSTw+Pjf9ms
3xC0DKKB2K0K0z9Dls3cH230HSW4F44L5L1SKR6kBUZjUh5/84wsIRGegca2e8HFr8tLYK5C5RM/
cfnpT2ZYzyRfePdAv0TZ0yZ8OppnlQfmH8acra8Q8NAPWeNMgNOgE90p1XV9rH6BjzxEXNpaDdFI
xMBh+ZNkxBririxiygtaqnU8ybA+w/KQw1NXSH+CNYiGZmPNyDS0nah1ivwJ7d+ksGGyZnfqrTDr
hWiC9mleqkQfWXdHvClA8WYghSYke4+dUSoe8wbB41MK/VnVCn8o/ket1LcPBu6Sadnz2yIEKquO
UpyJ365DuCBykQ8CvsY0mGHkCE3ChxXfZqnFzbXXj7cBnMPGFuNccx/oS0nhGMW+0+k0qd46lS+Z
jxSCvPUwNSygKP5CyWI7x4+yCK1H3+UUcycwwmJ6CagpwgVa0B8U0qxBeu353JtAS0sW8amq86ow
jw6bW363i1lVBKxMk7ge686+TIgn1o38SKNV4IgXeDFz9XOajq3Zo5ieYcwFv4simyhZnWyivrqX
kuyEp7qUuMwftCCCvokgLpdT2DpJvpu2RGrul30pwPiUAzLxJEONUT+Q9O+fW25uyoPIJVLsyL9M
pDH0GtwYuSzagPwPfGWAArHxxCnxm0sInT17xnfLanPb5wDlwee+pOSkaydhdPUlYAiKl7dpI0Hp
pVWqJXHI1BGvent00AF/IfynGvws3HmToCOvydxCNFtBKUSQNP/j1RqL+vJDThwjuhCN+yyrpo7n
bR4OnrGNeu9y19SzTc5IyAk+R6GV5Nx/E62PqClZiBLK8xyazXwMbr0n6oqWMrJzodI6En325QYY
NWNQgMa7DNnDAkZKy/RiVfRrECJFHaM8CUBqG72M3C+hDLao1HACHjLxFVdZyHFFNvWHx7h0XuSh
sWyG77imq9fTdSccQQhn+eFfD9TIdMw4mvcgeNjljD+wq8b0/7+i3knT/Pczozuu3dlZz1J3tLlJ
a/3iHV/o0aOcMB7A3Mo93NNy4yiiqQi4nZlzPx3dsPfAUwTOkQXrxo6dUJBdKwyJZPqI1sLt3SQO
w4RPb1SX1WjFWshGNpO2+kJEpyVD9HmhRrCB4k3+WxAhq6K0ODtjv4xVOPPmjAFAb8KGsxna1n45
Fxjj08D5KzI/hs6lXXnt/filJX186veViqYTCvcEamjConum4D5bCRHSMjkJQIzvOVCRa02AjuUA
/9qdsi2ztk5MpZLer8v8A8oFyEyGT+4OVysJi+Ki/1stQD9ubhFqjSfA4O84J2wK1GZgU9/eVvwg
zH/BlL719qHHeF1WaCmhg7Pgs/EjrndemORVL/RlZu4Y8RuU0e4Zf8LNFek6Yp29X7kuCboYh+b4
WScr5NwFpFVh+bdgIfXVHHXinUSSzzY6Fnlo+SxNWvWbpWBQXua/mi8SxiqmDpMzS6Id9GianK8H
U5NSDVLDb+Jv22FM9PK0ckMUN1kirU3kzMawYi0KUEsr7o/DDvmJagKOwFFJMjx6LPIsSRJ1g87P
LXbnVy2bTuB3p02xv3FN3oR9I5kpggBnM9csjXvgDvMrEd7ku0khLYfR4lZAhgncZNj4qORRTe7C
kewb0dFR9NKgWCQvh9IrH9Xufj3Uf8oN99f7F/r4J1S0E5lPEsCO5h+3NyoXPpBneXex3hyzUKQp
Ghfq5tFwUrpch98AC5tHd+Ydl3JsUZJkk4jp89tUnicK2nQVZTqaqRk9uEMedOw/IZMGxTOtmBGg
s/Po1yEYIoIdahT05FBDmLakKP2nIaRI0/TYejrIj1a0nVD3YshMsTLGRqdDANZm1UP3gh1lpReC
QoM24KnP5dfoyN9lrgitX4ubljmjAlcocLS7EONMAvrup5/hb9VFa0l/cYHku6AxEYwdXOuTwGyT
avRevdehOLBdQvdOmFaU7QdqjOB5opHxB8mdnEt5y/CPH0SwqRspBt+jQ/5+0NzHaHd0rMHnL2AV
zbIezl4dUYscnnE630OF93iPV13fGFMov1U41ZKJLpvUHJbj082fMla3NGMaa3PyHlxA44YaNwte
6ErcWrTSqGsJFSORUSAHEUZmDpPiQUqF4LBYL6vTm96x0tYmGLAqFOhC50vDqu92RYD0s7WpDPm3
IKGSzAKF1ZHRjWz5TY5zxJgzaMxzF+QrRr7zSRECktO5P+G5n6WuwBpOGqsOgBN93xTJ59Oo7BvD
byVi5PIJyvztue6iYLzBod81rVs0ckctlNuQLHiQYeMglk7Mjp8T7Uv8dulFRO2js2vwzntYgKd1
4IrkH68HscA+hmsT+LnCU/A7TTH11IWTF9GF2l95QHgGxA8nncSNT3+LIJv4ts72sAyrQ4ujZWcl
IhhrAMYDfK4yvqzOiOVddXdsvnOCiNf7bjBemgRdFYiwKI/skmJyrDnYUK4rRT/IMtEv750MGi5/
qmkIzufCgu+U9kU8FgX3ysXN47CsWsco6wWQhAtmSykaQtDe8kMUDIYkjSOzubvmq8wGblVU98o6
pGJylQb8XHY9PnXcUupyiTOeUENHknMGp2TGbUJUKiN3dTfoaCd+a7fy97M6Rk/gCKPa0CFPRRdX
kkAZ0iGZPH0h56ReLii5xtJ42y1RzuWwjX99TIiT6qLeTN/3qDPgSyoKfpK6NGcwptSS9bzLI9Jb
SwH0vlqdvQUN6GHCddfRgQeFWpDUqwft/uyTF6J0rWx6Zjn/Gdt2PD0b2nOPX8az9JVirk0qEis5
yiCtzQzeNPwka0HET/wFxAfx2r773CjGdkAE7C5Hp8rAVxh7YFSGrkjl2qrtGdonJWw/3RmWO0Dr
lG07mAqeeIGVYAcAnOiPk1x1XEQ3xl1Wm9FrZ0+7x+8NB5AgqITjFCbCAPz9vdUGxEVS1PEY13Zm
c+vIuNiSBLu6HuZIlUujhm/XiS7+/pFvSx02gwbOGrGLs2IbxoDd78KUvz5SjoMe9tU8wFyCEQJR
qwxcKt3DFq0XXN8ZBw98AK8mO+fI/b7QBiJkzT/nfukTYmzd6dAl8aChRJP5reQpqf3jYeb17obW
Gy4nWwH6c30/kAN/prmUqvoPdVEUL9z7fILV8Ve2XQMHqaVfGrYyby24quvvTClSF/pyUBwJ4qLX
v5XDzCpxwT4aQnnT1DkqnwDUEshiOIYOtfY5sp2IrP3M6L/YbLwGgcW5rgKAXfZRZS+hHscfxJ9m
ST17EUF/1BFhWnGyMxGKg05Cwhd5q1R49majWKFGnmMibnekifZ9UFVsBmyxyHb/DM2KW0XOvJPi
nYwCtG1Ufx3XWVXvlPJV9yXslOPDe70KrqNMZM87+6Ua1U9ZSpYjoK+BKoUQclBNWguz8iykG6ag
ui7dLBO+ztSFcVIILOolrCVoGT+g0mW6Kfg2VtYFj7nG05E/4SoY4M9HTRwhbJJz0cievfVD2rRu
ExAtsnlG1KEc3pBG48XDPn/rKAJFPqvI7OOApcLCRbkVUyBdBGawXU/5VGVhuyMlbXuPx4PJoJM7
K7IEcxUVvKHIZkM0z4EAt8bYPbgqUFIDCMg8UrDst9jdjjvTmXv89pdUMD4LzNH8kmx4Euth/9H/
mIUcAt0K7AGzTRFdNjGneBCiduCqHuXcSNeNiiSvLoz1mxT6GtTlwkxNpjo9v+dgBUs5BItR62hw
kQ18JPaUrdnzoWMwuUKPS4datr2wpycFhwLC9cdgWuoDL+qlNPD9bZ4neFBDfhZix+5OqV18Qu66
lqv6Fa9U3i5831Ggv5FwP0ZF+Nyhe3kKGigCIFtYhSDIMXploqhxxLyZaLBtz0NVaG7H0MHHjvQF
Hlpt5XCwPtGxf8wg820ZyJjgLdlY6i7lUhKNkUer8pWIAd7MT2GSkRsqh+mu6Vbgw3/QrqcptNMW
OALrQ0dGeXQRAObS9230In+aLoQ7i6fvcSdMm9/PgIF/MS5t+vhOUEq8zpDT5M026O09yS5bjq96
E5MJTMooibVOmcrQBwm9ZHIc3Hm1xKhQQrslOwRxhKXI2oUJOSZ47y5gnWJazUvqYtB0+1UGm5LJ
I0KUQfuL3zDTpa7DcAY+KztVU1VhfOTnoqXhATxzM4LX5GGpxaOVwBieojXpYpCBkPPWXIUTPJbr
pBlBj96/iPPCiePoJKlZGXNFPwe1ahBQMZ/csGSFlaklTWSdrAev5IWBaREgCPqW+6SlCnTh5ZD/
ayg9ivtLPiJzjmVXNrJnCx1YGoO/tVNXfX8AsPwO2Rwlp8QxDJlYFubRapFg4jMeIDV5oBp8xq4w
Bn77XRpbEOC4gARq/RItyd9dSgdtuE46xBFdaV48nWapEknl6a2qMhCc5xnstZWBZB0z7CkIY0xO
plY8l7PdlwpOtH77xJ/deGdL1KPnuGWqkZs+HFTq3jju7tZQoL2CN1CIYawtJahH+pD/YhSxhMxU
uxPZSAnaBEIzQuw3wKjRzraHmJElvxcGqo26Ku3sA869CSXONyzWF4xHRYO6NA3eTdsLOwz/szKo
Rh/6oygtA/aszePMTMjn2NjKnqgcDKZX/IFrPpkSTojgM+Ez3PKoHCm58vQbsrhnpBta2j8g4czU
HlmKHXPT0CV7GL5P/cLHevPXZLNxb72AALtDd0hTyBz/kwAJpL28pBTaqm8bY6JAYst7/7B/VJeu
KmuBE9/qnNCVBlPV86lj53NqefmdG0JQ8GOrddrRX6Io4hYqAQWJbsh4dRuJmWO9pC3cDhXwcxk+
BUlNaQRRAi0kx9adgHI5u6w/ClkJdDePw+NC620LlDrssV1vQhzETnUf0VjjdTDIao2WMCLLT6tI
TKqMX7VlYly37s63bJKBjnx0FocJiBI9oRUzsHd3GrqnmI4xY/jXuyL36Tvpc/0qVLYhRLhtnbkM
3nzxIP2Jggfbg8SE+yqnZkKvp44+G/0uJUZFD1pmm4SIU+yAVk40IT+Ii27TQzysV18ObWVkOHaF
oL+aGxV/Y1mAVHYbTN0QWMfaXWRgw3cBLojJMJyHkW0PGkSrVbHPb6LPuRR3GWh1kgW8IEJJjmBu
FaB9BWx5cgLt8rEoknIJSvuDIjLvJwOWFZyPq+EXt4MECmUsFk0NzbOvWBrKDGkW/NwJxbwToiii
mtb9L0QNj9NfWJ5TcyrA3PLm3k0MrWhCfYsxpFRXit+0njCIxOSYS54jjPwquyiKmH8HXDR/QbkY
9BNEMfl57fhtAPtB+PV3W90VlKBsiboXwa67CWIAfKcNEitJkFqx17QBk+8PlW3i4tbrqXlKjKAI
exRLVgrF1g/kmI1oKcs1ZwKjlTpmcT4d+hwpQV5jrLdekqjQ8/hXbYz5PJe/uKrmYWXrkyFG/v/3
yfjBXW05QNTVcf+uHzXIdeqXVc8GefrPELmwSj/PC0atRZWHqweRvJRzUl1JHInHtgTAyMAd4X5j
/9e95cEfBknBLwUgA9H0mQ+ut5/7kiAkA6MnGzdsHB/+mTHnL/OE/jNOFe9e4hto6zwsyw/p6GuQ
s053DG5XqeIzso3UA24RExHnui56+Tiw/18V1XnBDF91e+9+ah6WEC90svR8YJHv9jQmx0g/0/gP
GYNS4ssBmlolpiOHldhyFNgFnszkQ5Mk7RKgs/0UoywNffO+bCJKBNBcFxYXwbuWpVaZaNCAsN7l
um54dB+iaKa3++XRBi/NmoZ6IBJBhGNN++17zN79fWWuBDq5XSCrIime7w5NSAiLyDHhOcGx8roF
muf0Y0Bqah23wzce2Fq2nKhGCxalcXyWDi/hD9hHIw6d9BJx9xjXiYMnR0X0EYLQ8EQiJmN7fA1P
zSrjAqqdMjVgos5dWS2GLYVK4rZ/+EwwCiqhz9Y4QqYqQUmZUL4AwK3mOX/NrYO3oyqNHKdbq3me
FWYar/MaebZIRXWFHDfOw2UonxBI5FRBi3H+C7enKtPMRIR7jFMIQZn6apG/MNbjiD5u0J2cfSgc
FY4XzrH568e11IsCH0IND7t13yPaJxsuBCuxX0vHcWhN3qbtEVpbm9OYhuskQhsiQ0j0WyJU/DXx
n0+qsfbyxIiUE6v3rKvD5OzM3OJwgYx6pj9aqt2OiRDW4NRtvJOHFvCcELgQ+9JRh8raiBSUNkVg
azhNONL76o2+v1L5oIr2UxUv8L97TKi9SsR+6ZTwwTDClca7CpfZp8PyvCcb4HjLn35TSeK4gdLb
wj6lwAbif+3HjG3hTrnCkVwiR4pKLlGQrjyl0GPQDeRxkyL7LVFo6WuCdpgueZokNNpeNE22gzte
VmYk+Oenld4tP09Ci1fjJYS4490q/b/4qloahATWjV+c+utvmNvwjE1dIvOaGsJy4htxh6pMkd5T
RvtgrYaky/sga1lszurMCIV7OSCC4YSxDq05ikqA73vf3g2sGfN9rSiblRnKDkKGePiu5E6m0fsR
Vq4EpAm6eYR8+O8ltPL+DrlykGC8djzAx/N1fQqiFYaqEP/ksrQQZjixI5nTlqwK3pi7gsRSx2e6
kbyUsInWKuoyD4cGRVrUGL74ZPqFcHZi8fXO22fJzNA/lVriEBM8yNtoPEd2J9bUZb2h8KPb5jLB
EhKbudnwhjmBIt6S2zI99sH+R6EbWHFqIdkDW/dwpKIPQH/UhVAtcKMXfr9IOTo7NsN/BtgK509S
3qboaPygdBZlkrEtY6aWF28A8fvHW6GhOdXyb03RbmTbaM2UrscvdHi6ymhOb90NuDNoVynQh6WT
8dzVQR45VVnDUuIKNE9sehTmVAOn4IpWuUFs5ASTSd9ob8m+tzSstGmTDrSBcTDX+OAlvaDpc41U
4QxYRdfXMkLen18kdjVcPYg5hheWtcmNc5SwqjtFxwmLfhKKCmiqvPUE51P9wZTZ/5UhocLrKMHN
34MBGfYsSo6o+50WatCWnlXVhssRAP/Gn8xrCTkBDAXDHWcX+PBb9GIv8v5LFcM4V+oDIxsEsHQp
BlPUGws3aDlOEqE7CqVOUBchSHGPAQGZsf0jbKY8huL1NcO0m8BVjVAMe4T65WB43c2d7/Ez2Aj1
cgwJ2OqVRZXAqFNkpLxcyyJCBrYA5Hf1kx327CoLiavX8hOMJPZtx98uaDyGS4IeBsgg4VPGDpDa
1+naWr8NDGwBfjl8kAnNsGSLcS2WC3+MYeH90tVvTrcKSETMgZK6K8gV2TziiWHKhlcrBUq+bJAO
apzhPKCgcid2rHUwQS1gTjXObWqzxV8aKSJSI/a8/xxacLb4x9y7twH32WFumGxR8tyQVUn339Tn
6xKwA7cGjQYulN54wxkmaXoCPROxYxjVIwOuI85ASuBg96ocMglYEg8Bhxe3pUY23QnyXvRmsLr7
oqMVCDW7/ij6sNzEXRI1N0gJ36rBpqh7PtmygdRG1DrBvgyAt/pH5fetYb/cty0fJx/lYEsdLaMZ
YZbUmu0xzwmJiXRB+TcNhxQ9F9svhMrHQQ8V/0jFN9z5kRk/9Zx11C7ZrbY4Frv6k4w3TXCjqOkK
trv6BpJH2p/uxEs6RpL7XjuHK13osoDnF/ZLlavtz5Cr1ajNL9OkX2bQgWQBpNIhLPptPkNbD34l
2zpNxv6Lo2t9svI/l4DtpX+bPY26bziyBpLGi1OqASw4Nlyw+OVMSudCgdEjAuQjec0NIVTrVNNH
22Lq1dKgh7gJmYDPiOoXaxZEYJEfGLItqBkqqWd6BEWHVTaspz/nYG1RB2cjbGNIM/usL4yk6nhs
g6JjZCaVZvd9Ht7JJ6v5xXEvEvAz46d/7voSWV2+Yr2SoNsQgssn9gtzQTo84qLrTggJQEPwWIvC
ieFgXrdkiyaFr7yb3kI/DtZX379In6mq3vqZxuwxStCuMFzbNmJb9UErL/F7Yb7UXUn8R+pfT2cj
JE6a5NhrWNnRSQBBUrpQqoImhszcXZ6hJuVwUy2BbB5fQhXvsY3jD7gKgDGKArKKa6HNbdvaXUGd
h6AXsPhjAMmbtusedyHeZ52SJO7clVocvQbCxswjScqWgNaq2jkUEYVqZ/WbUtKXUZTk70pcEIHg
WBGIWllMuWK1/uYIl1btuMryuMhUy6C2W5rP4tzleyaMe0zibdvU6luyynJtodoF4V666IjUww+Y
f2XJQj1SpedWYUEmR2Eyz+7VnRwY/7IyxuufNOYYTZ/BXA5s+zfgka6pBcCTF8rD5jhYtuDyILwC
XFw7J8x9/zjNP/Ro9JW0l0iDW6LUa711cOZUSo9orOZnbeuPTgj+WA+tb+mekbX+aD2VwPH5fWEN
20elq29nhZ0tnA8G+fk11lrsb65BEUtjfsEwCwx+wiPDbZmHjd6oyCdJel8G7l4bT2KbzeTRexOR
6edww6SBk5gvCpdg6RhK7EQ58Sb+TIu2BCJ/GqMv744Z0HhII8ujdH5d5MknzkQjqmWfvQ4Bli4b
5U0JrfKT2Fr1s54Tk4/0ucQOrBPzA/+no59NSQZB9GXj9CSi88ZHmcWW0oCXyhdKpVrNrX5N3fMI
xk6D/A936t7tiI4MvbfhP3TbWA4MRcDJ6FloVUTSZ/jFoX2Gcf4oP1L3ffalxOoSWwQiTxE87LLg
TSLdabFr2Zh586AE2mmYkkHArrBRmFrpHbBmRjWdezPb0SQ7QC2vCLWZEgEj4Wg/gmiAZHISd0s6
vaLH2ivFs6+c5knNqeN6z1icAhWJ3axgp4HdmTSUbUQoq01w2g5T+I73ps75xBz4UakeKEnNK/Xu
PXzGC3bUr5SbM8y5zPxf/7x2IaUQy49NTc7qefdjWnUd0Pz0wkBMyMnsgMcIOzVQ2ZEVTq2YUktX
QsvudmSeXPXGBhLgnY9CKvmGlpKinN8XHuGXskfcD7aprbYiMW9/ff8+fA5/vY2q9LJ/pit7MRkP
/JONgyiKjE8gOxFkz88vqf+PTHqd+76vdCNp6kcPgqdEs47DND0m2KGhkikSpGtrL37DRNFNiSi4
Czadi2bkJ/no+DiKSDal1VsVkYzRAuoJbHuO2hXRE7Nxkv4HoKePZ+oG9foQhEwQrOVWiAShpGfP
sbcazw1BNUs4MGHDRpV0fQOHnymEOX2ZvcpcUP8nRmAb2yomwEjoM3ukmsZVGaytz2Je98tgykZE
V6Z8zB7Fy632ycnqpJWEjYUHkEHQX2bEN6dbyc4HWCPaqnUAiZBvr0tiiLjBLV6HhiU55vuDJkg1
vOt5uLo2Gf8zuSsTtnZqj1j7pH5gV+YDvx17kBYLD/6XH9hl7rTrZuUGEFk/LrHRZw1x1U+zy0WT
x/1XED6pJT12RAoIsUjTvSN/6JZZmudVZhLeetn6fwSeV3Kp2PboRp5ezWpss2hEZKG4DYgaYY0F
n6qrwryRt0naVJc2p6Rby5TMTskC1LzLu2fWVdChugaHxwQIH+z5+Qg1vJUGI+26UmOpNc++J37g
H9+BdtlBSVccb+ZebxWpnswJAzlC+5FcQphDatcX2T5uBhd1hzjSyPdQhDX8UaTSBo4v1eDDhFZ2
+6kkTGDhDVroPrRRCh8vau67Iw2YBaLXQTjtuqHcHmiO6wfDSaNPAT0WUtToqmXJ7nlLHYsvjZtu
VGV9hBJA/vsM5lGu3SlI1+6UC2dtHaA3HLc8GI63+KHHmGGIguMP1m2j+qPFotHhgK/4hED0nAFj
2TWl7VTd+nxofHSyr+AI+QH2xHcr9pTW6gCXJirMPEAoRfE1K74KKN8qD/V7Y8N7w7tNvB7Kp0qa
BO+RTNPy3CR8TCnxKHaYxxikkJPtqKZx4xNmyGjOiYAsWZgffiyTC1h1m3AQW7s/kbKx3D+4tEAr
nX0rllAdrEXwA2/Zj1n4P1XCYjQ7RjrqCpukiG/NVPg8+tGnpb9ZT6Iv6yu1i8I2tpwGgL/cLuUg
QVe8mjdj+/YEoGpdXZGshTKZ5RrKO/U11HCoy1ka3vf/p5SnlZezPMhfrW70ABJ3PFdj9CA8VWkL
SdCpdKCkaIDlMrGd4bdEXdCUbVBc6CFnK82myBBLvOW/pxLUhBLl1tIvarCv0KnhR4fcbLiARruM
O7KGMJzOOxgzBBLmvHU1O/j/HehIq/+LZqFxnxoTrngA6/mZzVNegXyu9tsYo8rWi4P+BdJCeAi/
N1K3FX4otRLvWCMvDZi/cVcUIwKmvb+TVVTE0zWprrPUdU60aG0EU2/U++wq+kbE6DD7BzoMheNI
kNfTx38t3Bfst+vtOUoaTwRLgJcJa5HSHg5v+inr8huelvlahRf0/vw95MrYKsrfccqS+xuFmEeA
uoMaqIhI3IkiiypOddQO06neLa2fM4FKtw+vIAAGMfnWx30R+EdXmN9rcMNfbcI9TQ4Jl8Ab7R3V
0HJkWgdWYpX7d4EPcprXVXGnqQh4cTdbf+Jrab4vnJbDoarqt/4oE2HUsJ3+krGNFnN9w61XAbG5
ZdnNjbVTaGsEouccH+WNSRK0cmYmv3qVhfsBveAGnlKBRS8Fi4jtjMab17G0vyAcn3xdNxRn4aNW
8oqICUqJoAAHEU9yFBhwdnp0N7Q8UqPsmqJKtCUbnElqv+4j517t5oQXM6FvAvclnyfkQZ1tAxT5
IkFeeL2vK8mISbDhc9pZrq7A6rRv4MLmZrLlxjghaD8hzsm+LgfAXtsb68PD/1a5hlAwYouwJipG
aeQaHQK1mJ3d/gRMpmtOVMpw1fw6sn0L8/fiWC9ZEpsU4LG2+mAG3rTWuCLNKQEhApTxCy9qOXTr
aeOpcF/jvUGxUW0tOErxoqbwzkbH+Mu36SoNMD2nKk0NeD983FOjeduINZE8r5T6XV7hV40I4t2h
KrykMsOK89SJTd1mBijJY+nN5f13w/ESrVZ1hnYYhE4f5lOimduf9Y/5fml9IzeDBQg4yeyLZQZ5
RfWRF9uX9aLf6DRtLLpQ+FI4Rk8RxXBFuNWMHFFwYMIVuMgVXyHfv4wSc3IqGgqzoQU421Sdd76q
iVEOYTGLxZdxxi7sAU2eeDcGT+NaCDX5+YXI63bPnFKQpS7SkHuzVTqCYc71dS4Qy7ms0yINtktt
GKQs01aBMrY3Q3IQYQlLIazV14F1lmHZvb1u5KOIcKNl6ozdSxg5SApShv3ZmWNZhMx2n6T4tREw
Do8Gss1HsTRYZwFub0I8FFYMWE2KMLC+z6DFI3Mc/aFBsuNVChrrNEb6KQH9uCkMdRWXvVRAgtCW
o+Vi5dbfxpjENxpVmP64Z1q8VlsT0/MPDJA6lNrWFwa8D8ft+NzchsfpzhI/Y+7plcmB0RrhL+z9
N0bauA9qElB5IENLpnuKq9eyL8lB3PZs7oHtUWg1GIKX6TD+WsoJ9CbSdHO5+pQppkfwX59TCQho
mJSrzCuieRzAH6p5f53OsA5G862cT8LXh5I3Btc6lPr/3z+5rRBRqhNzSw9eIv3OvMuXvbOtiyly
vdEbgplBzyp3t/ihPSVU7WKVYqP6qFQs+uT7Y0DmWVArgQqTE4LhjV/Ph0cNaYzoPXgoFrBzvD5a
Rf7hqAR+PSiNiqNiBUeHd0G6SKfqsmeBGWK625IXBfIpzrfieVdX3NzjpNOe2ZfpdIfb+Zfogt3j
I45Bqagjgg8lavP7Y2784w2G7QkI8qYziM1Nl694MhXnQfAaSAvAji9+Y8ntSQKCnAYIg3+WPdD6
2KaD5k3qEEPLxZatU97FFFIaqWbfjZvCiuYVOo/w6Wq+pqvBh1hMr5JXvdiskN9zG2iCd3Nsoudp
HIkMD12jYMPD/KThPjGBlhX7hxHFsJFP9gnHwaljDBi5Wf3oPQ4PVMt1SJz6gNIwkSa00TLW5YV4
3CFMIDejB9e89sMm64zvCBOec7T1zeBsU6tEn7tmOJrrBGMWACLOEFvmfQgfw6YMDedw47M8VFIF
pO817yeQY4GcPIqaejooIGowAMqTTU+RPd0wv30pA/aaz84eJ/XmED3ejdaL/2s3MQa43mYRBjKE
cGsUzPUzCyuJMnUsArBSLYgDONpiDDHm+pSHPE0pnN3UI+AeZ083iotLAM8fprJNxRIVDBk6NjXr
pSvgAlPZ40p//9UKL1FhQp8gvW3hI6j+VJhe2+fpU1G9cCKUPIT30kuc2ubKaw7FfNcZ2fDdgiyY
e/b913YShdML9rAreLUO9ARsZPl/CgH3OwGm+VODTb47wMGFEHgdloH2ty62F2tj7eG3/Wsmv4RU
OwVcCKxpNNOSad8tEuQfOVpHp4KlwlZlKmBz+k2eeA/OmqwqWiN76LSq1F1H9DKZfwpiskhyBy1M
GEQOyMkx1JHXMCkel5npouzJdJ8qn2/955ELYxo+6ZZtSxp2WjABtzDmv6Dg1dGP3lw5+Gmqk4+p
wArtoHfNcHq6t06o0ezVGx3d9W92b97B9H9EbIG+LHQCSA+Icb+jSJX0iA490dE76zHHO1Uxfac5
CGYYx/SxfNGTydzTkoQzD4E2nTZAN3YSkOkshLK+N6o8Ah9WGna5c/xAzU63b2xuFfp7RHQAY0OG
vtXGy9ys6IYvZY+2upeZC8bVDjRGQADr2vbWF19PVtrBeDl7lFNAl2rkytQBIfCJdHLO1oyw/QTr
ukYIUrAH22M9mhBlwG1KGjS08LNli7AZ+cE9ycsDuQ2c2pYSTInSXJyliPDg68ILKazLJ2laN0jN
D0j/J8NOsDZrtvHwhb6jAOpslj7NGIBkPpgTSB8EmWaT9KA2BhTSWp5YwsrHWNqtd0Qod/f2ZoOj
aPPQ9Vk12BD0CwpA3e+moubvRV9Z/flPXy3ppVCM+/nA9mDIEsjE68dmVbO9LsWUKX66JByO5zGR
RF2/Ilnzo14C+lEMKteYtZ81Hn6gUUu0axmY633bEvpcVGXYOlwf0IlfhjIAd4Anu5j3v+lXJwm7
q6EQOp0iT7SBpOooKLEg4ajujE+7sqLtu3Evff8kP9Nbv9OgkPM9WXKTHnVvEEEO2JW+HnKESMFS
K39fuqRcKNUKS9P0ocRPrvSFKWOZ+aVD498tLdq2fmlrNX6G5VD4FbfjP5qFMvPPPo+83LO46a4n
EbmgPKHAnHcZ4QtywiwCMGeHcmzUTtzsE0qoQeweSih4OpKYyGdrz3Xj+qWLbImvjDn0d6M1XOW6
fPJE+dLH1Ag3bj9gBk9b6bZf5644CIE8FsLI5nXOgRVI7CP0y2aE0wGvm4tdxoGlL4YqHDc64vRk
/q9/jqVxnxSVwVd+NeBupcOZcQBzgbOB4YUG+mOYno7XttjIkUnImed0f8O9i0FDq+KpxKwyGwKz
zLL3FYkr/1J6XHjfx8opaIaHBIB12b/Er5kroUPVe7L7PO93VDc16PdJySX+L+h83I5OMKTO1a9k
13gwLzRQnxCB+yHm5xPq95wdWNWgIgMQNW83gheIGY6reSY2zL+pJjAgZLpNHXa7yEVLKhuYgUhx
jEQMd+GRod2aKJ8CSi1dOWMOdMbXF1kF2jVm6L74Wmd8vTNcMmVarq/bzgzphznHmCmMqEVzTU/Z
85F+Z/Qofmb5BZnFNCgJv41dPQCAxwppsMa0eIPOjI7HSmWw7G11hTeAwmLME7AUkAw8FUTSiPZq
FG4jd7E97ZxjS6HsvgZg/i24ARnLql7HVcxfEQqXTwi1J0USoRYavAnKCpOkwgDMEhk7cBV4E9hX
b4Nly9IMcLbrf3M0fNb4+W4ZyIM4TLwZJsbJIl/k/mw3PeEFgU6rCPLrUD1MxAK2IOodsCg+33dt
NKhpdoIHzeT30qX2nCpWSk2mX3GQxx4EARgXwkgLGP6i302kbMY14J8AYlUAL5h3kxjo4hCMbI6O
3yNGhuohTniarmBhGaEA2aOD1T/luK+25RNzkWQX//PxIVaE8KjX9NnOrXNBF4qpncdIgMGhhmEQ
3q244z+2nZcQpyZMO1yRANbGKoYFQ8i5Sy7Flqv7hAj01di4sNdOBcGRVz4EVL7cWhrr1EfsDamc
g2/znrFY6O33M9i13mAij4KmjOfLyVZuc/WslLMFUaMjAW6q3MVMQCoWvdIpr7GUolhUJ7ePSC+H
TKQg0zXn/npq9OrwkYtH6AICycO1BUS9SeI8TIO8gqKCmp8/CMiL4JzmCZa4vJSMUgMxubI6+t6e
uIXZnc3McVzr+bfx6qlZJcv5oN2O6evpn3DK63sJfcjrNUex0TBsgnAdsiTcgS94Di87uzH5QpmE
Aul5LXSMR6xQzZWnYxZRIHWeo4E/jglqdUbtR5aLEbc7bCiue/QaXp+45z8jAB2tileLbvTR7Cd+
7mfVs+QaX0AHnMbDTA7MlzZkemfJqGPqMDmlaRboOhnvpnCZ8AVFeRkXskdwWC+gyoo9AXtYcdyU
5GPKKmsWF536UajAJorhJQRjAJoOnsCaxFsrquPvKfDJUvpAxvKJy7nBxX4FAs+qtkw9wklHuRFq
ODJpUZyrK+eecJKWa6zYEZjXwELmNdOi90UVMPLAUHPR1/6aAe8HJVowoJV9ylHv/VCThDa1gs9+
Ba7sgdh/shRRibM5N+b2LKwiy6eZ4Bc18igIVXbvXh7KukPBIgz/d61H77UmGHAYOIPu33WrKQxn
mwBjhQDv6KG9rehtkSvgASD2PuBeJLNYG2JTJ92upqSL1rdCSJ2u0EgZ9RNEvXt5gke/ztqomtRy
H2ev0kqz8j2R/dQljrvDicN0ERfDt9f7182oymgbSmByvq7Yi9asM3aIWOLUEuh2idBK3TBaTUp+
gaGCNqinFl2Dgt2NZDPKci17ESRVR3a4S725scMIJvLNreiuixiAFBr9iSyp87b8XF4vercFzXEo
jyOmb1Fr2uX7k+n6O2S2D8DTekxk4fDx72fJTtbyxt+P5jrkR+vabMTyLZVbsHKyIYEhmNecUB9D
ykeWcGlht87tNZBiNr8+D1PLZQqsKwp+4iUEoqcmsqkeNMkyOQJtxCHw/jq3N6OpVVFem8nWqMaE
TETbpFpK72TEJ/joWhVf+qzb+7leVrhurWA+8jE2aF50MwxzYW85FsL3ugNINjMNtGfskfn5ETr4
rPBGWdhSFZWpzqv8Dxs3GT76rYUgihUJPPOxxfpJa6aW0XYgq431drUhz1jqquXTpdH0Q0jZPLKr
A2Wsl1hBRR/CSucvIzPts8UtqFWPTpIYxNIvafYldtgsLIKD6p4ctAUDVmSJnakuz2pZ0GiAUOm0
0KX6Yu2J3ER5C8f3ifm7/n42a+ePlCsniNDQhRixVCNyGLzBEeqvs9IeXtS5uM88Q2eJaZN0zF7I
xo/U8IzUh4r42B0gPKcMzkILoyu0JYEHb92D/Phb2Mcjw3pnsaMvqybwJ297jqpGJ4gX6XuIJm7s
2T00xqzDFJFTy10CvNaR4rE7D+rZm/HWe0EEsNFjuwQZOeEt1hVOaY1I4rT451v3r4aaMqa+0E6k
Fr1+iGeW74iOiWxA227lZCtP0Few5V2K3CBc7t+jgcwHyhaXDer6tsZoYn+afaUUoSdi0aVir/Ou
5sHGKWllkT8He52uG1UlhR1NgrJm8O2RGFupjOxLHseCoen3opj8QRi6OY9iwe2piAPET3yz6nEu
9XaTWhyGZJyUhc8WcJOnCtHodMS9QMZg2A1eEoJkhYwaoWLwRrMz8yZ+cMaXV5ncd+k+wlVyBrGZ
/LvgCB9UKnNaaeKRDAn+VNUFLWPvQbyXF/lnEOjgrbJU1Y76ZwhEZdYqJMhIMh7h5q5ki4Y2nVM9
tRHS/2QL3MqErCq55cRemepS33JFZw6JWRGwMaMfTJbaObVY5Jiffv9ZsT0zmG+Wyy3MMxyqcgJa
fcZT74b5ULCXM689sOqydfjPI+EmZrS8+jVBwike59O2EUS/P5/+prUY13IpqwPyr5Hyl/VZSuHZ
gZNvs1g5ZUb0E7YgSDnt5bgjT+L32oqlx+QGz7gEtCMf/h4ZbVToEqF5wgbKvL0nmXnOxGAlDP22
tM1BBZ8m8LkvBS2QGQRqksw94PeMy+32H6J0fnRXXF4g/+2jOdozEOt60E0GArRPNd6nDKxEzPUL
J0fKRJvH6mg1qUszwiCpVCYs6mqGtnkgccAKKr5bTgzBVxn7P6bf0WY30vnlV3ZBGySnQ/Wc1lQA
h33TenIV+zPOGdOmQ7Ywr54pe83zBN8W4/FkkCPnRa3j0wQj0jqLjX8SE2tigQRxfzHxRWesG4iM
liLuilY2HGiIazsDQsDgI2mO96Ren4MiDlz+clXsVSAhuLOAUeEdaMGZxcuIl7S1+bCC9T2B1KOH
B7tThK06lDsRQ1xCc3nl++KAEuzifS1snrqJhligvW09/cJYu46elUzWcWpU4GYDXAvYHrFibNyL
by9HxJB0ntEEyvsaVVQAbzRKhVR/+1eHg90qYGuy5JwQLrMsnc7OTzMjzcgyqJRf9vRv3aztnB0X
XASeKmq4B83Wlbb50TD2161RhMTECTL39KJ6xYpMqCSQmSeEpmBWOp5Bi5QQ6CSF7uCBLd7de5Zw
CbmguulNISjUr2+B78ZLYhUBlLUFUufeSsEd9jPVR1s8phSB76xYKdN9RV7E+uTH8B0EVILWZEEk
UQKGBGcTDwkcbas2G1V4ANudloMq2zv11ieRe9AnPV8haYMQ+IJm9KUmq3eMcoFBC60EVKitDsfI
A5GYmgoGsEjAaausC0orsmADVhlQWGVeCiBFjx6KpFmwkgcng0qtj20jogNZhxFF3sq68gsPDtiy
pEOzsUzg7FAyxOLCwmtFhvwLLytnfzzyN/Lmg+H41KrwtTIA523ikYKYTih980cKVtP4NRnUqmEp
M67LDBNhg8gX0QSyD3cazYHmkKgMzJzVnE8J+1XM9lyFwO5OZUVmaVuhD6Kcf9ihXBU7OY3UhDLI
qW+rLOR+rXJugWTF7r8Ge1qu441k3fStnM/d6vAW1BzWw/WQuBgDlBZlU8ynM5CbFKg/tQ1yhtl6
pxUtysIAiuL6FPuMrKdS+ilJcEkgaKxSeBA3xzHRAj0zU702KQTph94xzns+cRaWVfgC3w5hI1aF
++OXndbQoMEe4TCQh2UfBVAUrU/ZpWpqtZm3B1iwFcwn0qGapt+O43ELKd8DNnkmLckFjsbApPWj
J0zliZffvyORrtkrNGvE7q5ElbqH4ygRvd7c58+XYLFDDDw5zXxsOeBK3VTPcgmNVwrEANKlZPCi
DXEqHK7e0szvCmVkrsKEDw1jHFb8+MMJgN+rNTXQ0wjnbgO4ZGZegph7L+d66YtIOIsWKceYbDQV
npFRMQl2nCzNhOB13IkjUTjweVghnXi9gWWi0R5xuoCRgJNOjgcFlF1cFpPCQK70CXmZXF/NhA79
kfzE+o8mAK3kLxoV8QmhIhYESj/j8YUtQG8pZkfM63QTbyhTBodINxlAhey05oOqsg7OQ5TERCjo
hvgxVHz1VdCJ/VokfB4RRRb3fEJh55KVp51Aozsq4xHeSXzPASTpCLDMruP9NH2PfaZC2xqphu7h
EcPWBEw6NxC55jpXs0lVMYpu4ZP1MWNBMWw0tV4ea0sRC3Via0bFtlx6TxsVi43qWDn3gIu5cdC+
Cp/uc7uIILABcBvXfYFegZZonn4me5i4cjo0qlMxNABGPjjZjI36ySXAEuHnsg3Dvu0Kd/ZAKlC7
Kk/m4xMYVxkgF3kx4y3QouRIwYEMyasLY2NsPeK9je1wepQK5/yXtBFpaORHj2fPKCoEbaXWys/L
XuvDKZgnCnwXwZIrlZ9XZuiv3W3FAzR3OrLDhh6wv8HC4RDNo5IIlpd33bCVI0taLVIHKFJ667iq
wqlOmNDmYJuEJZP1VaGc6EMMc5M6nwh+wuTnmRJBmUQq41xaeDBqkKEhNtCl0e6obT6BfmX5IBYi
8xERDKyqwPEo5hPJGzvLEQVm0L+4Bx2YPMO1TjhpwMmBMbBzUl8g1Fg7HVEMyV0952qMFWlrRABE
8r11fWluPuHfQAfEQQe0JQgIA8suJ9ZuRkp0Z1xkNy4UbUmwMCEltrMHdXh/ueHfvqAWxlBogTzF
yul+5dFrUjykYcQ+RVGANtpnHrDr6O4Ul85REOHzjIA4zNXpqXgrBLiM6wVprDpYILHeSj1JJmk1
2FRzD7y/sknMmQ5ZEoniqGw0GZbZxIEpavwEW0aRPQoLDcc/f9lfGpEjjQfymLttPgA2HPgQ0eFY
/eAOCh9XOBrtpj46JV4oP3DcfbjcCvQ3BYZUAMJVhGhe3Kr5UQd49Qdd3jI9mKuxUbZAbOsLxK7S
0DpB8V1bCYrIFogk8XgjH7byGBkQHMasUVEPlBkkriCGIVuLk8Mw4pVf0Tvd5zqtQlJhAuigE8KX
ovxLGDb0HhxI3gS1wXL4cgmM3Il1+Gp4y3qZb1zkDC7qMm+3f5fbGAs7XvWvmwduiZRMtqWBusTH
E1fZ7314Z9iqX8+CEDdBAVElE0sabF7NqArXzo37iYbreQiBbwVTqZ3qpme/K8DVou56Hdc0U+T+
bGoXB9lZjuevOADSYVgs64Py3P5ASp1cU6n7ZH4pPG0VatvPrwQEQcxbod4KC46sJQL4kR6HXTdw
IMXrfygn2LimRwk7GKIlww9OSCnUKdVF/xI/tkdymBLp+xE5ixGs0c7EEThll3kWDIml4m7wib1Y
set2wSCBR3xXIGrWlPFIamIYORkmR7uMJENyjJwuG1KGavC6iikXyIsBBhUnBPlCrfcqnZMZrN8Q
CWqpjXdHdsatKo0lzjW8UqC4chS+O+pOhP3Ex7Pxpy36d9ZxuckvQCvyOWZvQIEn1HpLd8sNSK67
BFvUPT23PmxxzRQT6gh3pOwqy8+Ss1dm13cHaqs0XAkprx3pRtXF1kN31f9v5cYzUqigKmduag80
9l1CxR3k4Au9Ro+qVQnUtW1xsq5j+H9yMCROHYJwrQDiNSOH7fptl1Y56IAyZxJt6gNlQgSYcxZH
5uJ0TYM6st3HyrB0/8SWS6NP1ivCWb3ImrV2yaHoHdVuqiYu05eFpMFc8/2bjsKyDtoeqpO3hILf
JWGkymaEn368J0oK3K/ATOo96gbHaDew6D6azz5kAtWw3qTMbjNb05BkYhUciXDNVNce8G1v0lz4
7N57O2MSzxpaxU5XZjsVm0zkCx9fqOLHRQzJar2qmiOSrrXN4kxGyDDPYrM8zvyPJPW16ssqE0Z1
zxqiecPwNQVvSfuXMV5usLkiT8b44jboQByq2tMFt3HDhoSbC1p48f1c79MuHjnhr9jkehd7FxAs
0XdjoEtnzKSt9craHyw4w9V80UtcqVDHXxTHLUHcxgauHJMMbjv3IV7W0Bsf3YcxzPhghwsDQNFZ
9hTEar4eUOXj3y/RPdWS17HBASO9chVD+a4pBGDPxhXqvar1IlzqZO8mDnLIDNttdFoY3JW8PDTx
5e8NguvMtRosTpXRT3SkGlSTz3OfUhMm4FNcQYnfwDkaEYDOCIwVvVDQXePN3C7v7jR/JvPCNNg4
BaSUC3VUACtWeKtcFVceu/nDg9J/EM1aLiSIeLGI7gpny+3pZ01iNL+YNAzgMXrs9pWn131TcnRB
N2pPjZhcnfuG2Q9anJRsotSgBOgbxBfeTRpEmtQi+2ViOfH0BvxhFnPS/WaH7YVFQyWmT3vnYK5o
+fi7txm8+bkmoOTd+WA5ZT1fvgFyQjC+Hli2C0fF2VN9llLBbeNpZCsvWGNyuyUrfh8Qf34Wxvmt
86Tpb5pFbp84VkjUZmet/g3GSPDT8kfpUG+MApho0LMuj59b7qP3PB5Rv5/wIM84axNRHTPJRPmr
yBt6D0qq4LFpFtYzzz2OC8v1cLTwistgcTEJwdVe6us86C+CnAqtgIAUztRekzVrVCF/KeytKP/Q
0apD946JK7x0z6WupYoJl5/DfKEmnrBmCTqNDEwnh9evd6/VXEuhZc8Vn9HCRnLg4buSoYOSiFKK
DGP4le6fZy9t8dlBI9A8lS7TnrVagBPTiFnCcfThZ12jale4hcoQpWdWxVmIc0MQw/HHfCkT6B81
l6Ze8rwDKF0rXCOrI8k4I5Eag3oY+SB/ugb85qA9VAEzQXwglV3aA3v620dgbvRtD+iIg6r2O8dV
jgejvzb7A5DOwS6yAZ1RWpZlEGQhaJT8GORZuZw60/5FEs9rQ8Wv6y1PbGpbLT8ZXGvwruw4u6FO
Iuzf/g42wVQw2LMAtOw8cb55UlgN3MoANcRpxweCk8I5um2xVZyNHfV7rz4i5zmofkni4FVVEyXU
qjKPFOuYFtgE1EewAnw0K5ubz3pIyrc/3vTqPNRi2qpukL1XO1D5T9gDuinrKqb6EZW+mj8LuNSb
nGAgf09OCqC3MEMtyKhzoLJZsTea/2Jleb6wikdYSWV4CEUZDRT1saP47RV1NY5U7sr6NWdsfzew
ftUj8feSFu2PuJblwmbyIweJvGSNpqOwZHPpSdvJs+B5oFLNewd9aa2a++QFI/DcsPWE5YbxR1ds
pgb66nmZZG34/iL0KWwENBJBVveUsBSRfm5XaguXvIzLWuhueu1xcQCLK7yPKgvqpp2X7wjnbVWK
74ohIwoeVN3Gw8sTYgAoxLnOYlmoFUlu/KA8BCVGT3Rwuuh7B+Li+fi+Mf0/5BWKOCADM0rPsQkZ
C9noOWm3o9I0BUL+wTsABA9hrbs4hjO21TWfEQ2y+gEc1hGcSn0CNRmjpklr6rKmzNjEeoz7deyP
QdS7ey/OEAZluipS1IDNcs6Ctwjz1S30urz1XTuge6ukFbcHwpSZMFsV0GG/iDnO5jvOJrh9MpTE
zEpjujPLyveAsN46GG0Y+MMxLsf/CLeLRcaRLf/SS0Sai+fGRlkhRedjTw1Acsjdv0D7wwavQ8rk
ih+UGYtMmiNWRQ/AMRc334q98opbwA4CClqHiOMnVa5fsFi/bsnX+AENlkZnKiwskTpL6ADiZ9YO
sSrkMxGlssNDAJJtyjzyEzGSfltZ3kG44x6Ye3B59uLaJ3kfBbUV+giDBbD1QfFXpbX38Nr4MbUF
0EejtS2n9YwGLUCs7PoaI3x3Ba0BygrKGJQ/Fm0RTLjB7H46Nuj2v9rL1pq6oOXQZ9v4LE0eszOF
ba9ZkBx7PJrUAqjPROziQQ3ECnbd/8hQ7GTSaC4ZDvfXGgwWMz+PaiGl9iCec+E9yoahdNe7+PQM
i/QLoXJ6H0uPqlyprja9QyL0bN7nzUvzvs4nqTlzPYgtOGdolw4E2vFrj6qTeg0S8aMLyyzuV/09
Fqb+YyM1B9HLoer2z7MS3tW+A5agYt/G+2/D8SpSFH/8Dqb3L2p8NlkDOOI4uaM2OpN7TRmt7CLG
eK8CZ8tGMNbNieva85kaKcS3bn4DU9PCfNfcQo7ooCWZcrQan9sua0zZ2PDkkTad/3IML20fPgyb
49q1mnjvg3AmoiLS/+OfDo6PfYGkjut3W9OHmwk2SkfZjT65gTsJ1a9xkO9F9f2vS2aqVgUTWqtf
vFyRNwY5XFkF0eeVz/MQUW0sXG48YAnbhGsaekWCTnvG2BN1adD5OoYBPDphJp3YXGHC+fLYHuzc
lcSqC0fPEx+7XEGu+S5klc9oPmadHr8s73h/tejA4aC7fMJuR+iHY3kkZLbTtmS1gJ/aWcJ9KTHw
fGIMPJgV9qOJROIIfDM75dbNpL0/aZ1M1IYU7W/BPx6ovfZWZnoWs5+o/9Sf3vOHcmLBE/XB6ZSl
P0qWuTwnFSBEuZ069RWYgc/e+n2k/R0tUR+b44YZ/fT8sgHmxpFHNlIZhUxcpNycjpw/+SAdA1sL
QpVTveGuF7ipJggsKuaT8m3YEaIkl+Qspr82F9022P2JEZtmK1inUjC9JWBGN4J4iFXVoaoNlIMD
fyQPUzaS5OH1tiMCxOu7hVED9H67wum4npTRjYzsCGzsnycOAk5UafaxsvAKpUq1uElbn2kjziv/
NUCCqqBW6r8Pjnb3E4Wen1SVynLTgPx8EiBUyu0P5jKRYFdrKcr0R3sjZch/t75IAoMu3kI5BYme
t9LNVZBy4Prsqi8Ow6k2V8N5ACPkaF2y4waCAS4ak2rXo+h5RLCILz4C8dwfgAWxNPlc7t3rHNhz
HteDs04ZALUqaFanb/5u9eZjN0l8fAIG2NHbfBV5gUlEoEpibuY5oEaN0vbH9heFudWI/dYEGGYC
jV+Se9LZ3aNXozFlRbYl6xc16uY7WiLiwh7FcT1JWdY8HjG1/D/bCPqpQrNxg6TzT/zqzxEl50XQ
dFx8IUZyfyAUIefjP5PVslMtb1c5IPV+ujw0MENlfvLHeDggzcB7P2cyPQiYZkDQqLqw2aOTzGX8
RW8HmtfX0kLf1TiREB/jrwoaJi26mi3TGV4/T3ifsYadh1tp3zr7ACXs282teW3881q4sNoZ5xpj
1CNkARlGnQf3l7fJp6BeGSKNLG1+8NgjLK9g1722iBCtxT9KVtrCxCzBbZCoESj+YCc3NBmwgQg1
lZQgfE0iHGOmEXBYOj7d2xzH/OO0lQdm8zgW9IPM5teln7HdUdD7sFnKHKzIdq2iPOAzbqWu+Zg/
hyh9dFP5sJjrVmFh0T1s9JIZJnl4xYlOHcLgqVuw2O8UajWupeKI1bDVkFXh0lCK6V4mvouzGJ6C
HianyrPfkOAgTXoGH0s1mx6CbIiThRpDyxj4Ksi4s4RNXxAJ/e+6QjTZvn78rmcvKvoOWN7uI7XF
euGGfZXUvT1K0cWJxhKuTc6fHSiKjf6xuYqH467aJIu5tQ+FMd/BFIxbxGBrJdHlYGs7jyMD92Sg
POr95VHN6Kw+ld3hIV+RVUqfuz1K/mxWWNRB/XdKhBTwgoYBYh2aUv6XldRa14LbeuewXQBZ1Ojz
UFPwSC74i20JHyADeRi21fKMLAVW5OK7mDl21l4UJvsK/Q1pftubgtvw+vIvdXZPot4YgqJ9m9wk
pJ4OyOAgXVOSDC+WMQihu310RUpKAXtp2VYDabg6znUnYw9Vt2MdAjWfPv2qjdSSsYxXR87s2C+w
W8tUKazN7rQEPj9tavBoXyFd3SYHef7RTbpYou4My+OdrVrjriIvAA2xJmqj1ZYK2J9r7soDmENz
NUM/YRAkDrEJ33RUavwldzrLedcquHiX9Fv/ZQxeEo9unKUNIkszRwyhw7bC/EjzKErLmZPJsTwC
stGinkW6aQ6G7PomxaJVdxbC1BLRrisiydBCbu+O3ksv1hQ7cp3MD/ZoStHUcbNPPm0Z1b9LQm++
hQgncHEEIXfA5UWUNH2hVERdbXAzPlGLi2bQLgflCYb7LxgarIbcQB1DT/8jFc/B/Snbesx0Tb6B
3HmBazhnos+eAlxLMq6Yh+wCNmC4mwlWmx+nwS5roqmUCO6QLT2zaW96aV47xhZoOPFvdOnll9Wx
9nLiP28OyJK0mX6CWroPn1K3yXZpNspyDriIXGsFBoo8EetzvkZFyUzPUwtCmzxVaMD3EdoWdUWW
Wj+QueNS7syUye2U51UvYBzY3OUWGjhUsJ3f5QxaLv4QCBRDpcteWyDucB9hFk/VStgdykUHxB0L
fhE+MSICOe2UmedqiUhKClixZR+LPy8HLRS7Qqg2onH+IZVMMz/xLHr2cX638TozROyh0+jBeHtW
ELFlkU8p/fZWPO2TAO1JMpxEqNxrj26aCffU26MbYCGvb9dmxQw3x01lsDpSoSEdP0sc3ApcZNUD
r1GBb/btDEihjShM+JXpdmTrrr3ANNb5Xp3tzkUpEQqv5UX5z9oAhN8SsxVf/3f22hwbznZRPYrb
lQAcS+gT1HbT5sl14suAsMvBkDdZjBn36kOTz5BNKIFD03fBN0jRivzCe5AiCoGZTrifDSQ1p6M7
LPnOzRxmppE3rVL5qUCAfHeWl+cvtGTnp8vMbJieGmjI3h8Ftd/d2hvQE7jW4hO7o+kU6IJ/UpBV
mcNlLmwNI4VLH0SjJ6CMnfiHnlSdHxOvIytJ73vozdg9RcT1gkvEJ8HHFik78z8Wgc9yX4MtPK79
im5ICFCRlhjS+TIKgobD1a4UQOFuAaBjQOrFDgx9nfpMTAjxlbHciPUynaSI4GJ/kpBbrP6tIRT6
gLzhl9C4+bDan50AFTHLB5/fUT/IGTni79sVoHnJr/yIFW0cipbhqPyzlFltgEWrMW0QlVT+TA5u
2REZMpz5N8K0j8pUPNP4mXw8vVww0WDNDXDf5xeJyrkGvbmdE2Z2308TLJi2JrI5GZcJBYdw3vh3
ZJdYqnxP/qhMTZFwObpiuhVKi1beNNKxTOfOuDsYA5Dj4KT+pHfzFRJ7ZWiujORucsd9p4lez3L8
/c0lITrKJjpWRnwXLoqSdKMF2sy741J6hIXyAva47LBOj1t1FgB5Q/wtA8lzu/9DGMzSAxKy8jXJ
aZ5RS6xLJaxB1Iia4sWyCaTf+ENRLmSaMgCUenkti5WWD0Q5mkZqeRqWv5AstRh+/8k0m/374N+m
xJgtjtbpo+1fRITuOcwxF8K7hdQltGDONhhmauaffmsbERn3oVT/sWvdP9+oS3xMyZLn3GCzub7j
+ymr/NILwELDQ3sGdHzG6jkLdMceu4poQ+Gp2hppPc9Ndx4zqGoJBMWFF8/UfABM2dxA5yYrIhRt
UwTFGLpOf3xUlTqivGS1/ngmleE9Mt+CvsXLobq5q3aD4O/bXq6/uRpRh386Ei1p5vOQ1LwLSXDr
DKSYCEEXUMQruLOZ7CaCLkgATFTzKXjuXH6h14WAFmte/1sBNBEwmoNOjNO3hVoj0vjEzBIB0rSn
LTbR7mNJcbP5LZjRNZC8OOH6JjaypJNmwI9+fOYblwYIPsc2n2VuUDyl3XHIVQ2eP+DJkdAstrjD
EfZwyOq0dSi4DSM3Aqg+ct7KjlS9zOOTM7wNiwvdEQYUvhYks2k/yZcdA/JVxr695H7PABVVmMDI
04G7iEIqh77INkEu9aKKJ5hlnGY3WmGeId/tA0ad/3ogaY4akSOUed2/0pph//CEWqkSox4PHcVl
umNKnsg4H8ZOBVWK3b9eEKVJF9bAfJ9MPk7lm7YSmzLOruY+RdrybJukZgYchCntXd4TXU4TTe4n
LqwMNlB4pG1JGTuubAHZlXVhdJ5Grqltwb/3MnPuXGz9ZXQalDr7SJVAVNlN3WhVgJ7U7U4mtzjv
27m7CoVJgkW5Rs0HmRXoITumF+4+SymZoFL7wc66wbQdQxj1j/N+5NBXE4sHAWoohjScA+xh9dFt
VrrA4VwbcL3+FHCvtIfZhl2+5jc2VrpM5zAkgmwi+24nSfa0xTbzj8oYyYKuYNw9Y6YhBVCsxItP
88k6B6Wed+h+p80iG/iz1QkM0DN10YO/oyVWPcW2Ek5Q4QuQm5kxJJ5t987LrflUcGpGStoJZdsw
FQOlvJlxLRM675EKYOFpzKS8fU/to4UR9BEs4Om8SkEfYK1sl6SJyijmxOfl4Qyh+/A2CRXAjA8W
jEpRb8LqT6jV3VqXptMeffgBbVRLZ7gvLMPeYpilk0UIVItaf6aT3vVSOE+mZH/Lu9Jcg7IyVXh5
tY5uSpeTkiErkiPG7sG/Lf6aQYKNtYjA7bu0syY9BLkcLtTFKaIUtX4gTM4Rjzkr/6pQ6zHO5ItZ
y4nW449q/H0TceXCYOHuOGgG1eTnMrNRKu9vbmv7QwONskCsHzwh5Js3N0AVwzFp2BetxmF3VBHx
QxBumIVC9BG21/+9StQqq8sfvIt5gzufTAMY0UENfexzGelvQitYwVUM8VUzHUj9AmyC+Usu2tm1
KTPpm7+rrw25Y2bzXv0AfEN0bU40bdhoHdTFJGU6lza0wHScDsHQHIrNJtYzpcYBnh/MBMd7aubL
eBKKQpAaJ4cJhJbAyR2y+mHN/i2tjiWPeD2vXnE9g/163Fe67b1OX67wxWTyNm9wDsXkGslPOFEg
K+dutUCFzKNEXrUcuZLaPHkA8sc+NJTG2KsZuaK/amFUCOsEMD2sgtvc3na8Fh64DX4NuqjgKRf3
Z1k6XYFu+m8cYPE2FpPP6dZbnbIqkRoypbSDvdKaMS6egIb6uHnP6cRqIYaYaWlnryK1ZakKwXjo
OeIXD6GsX6pAW/8xkK2QSSZke+30BRJupScS/l2bUN9cpZWGswPJk7BUIEAQ120gEYyRbiIAlelC
ApcfT+NyOUqc5R0J4F3jh83CXR5icHzdsu27M8R18q6QVV3JdwOFyTYudww9QYepBWxp+VVgykv9
IcVFKYLJhEdAvx7OuWKlkYFlszBxUpwafsxJq8F/2GU5cjxjfB0OkMMLb7lhICBDG5xmEqQtb8CL
Dky5mwHGHsko0hRaRKqSKpVdC98JzGuOyn/IesgblkZxwC5bpT8OqSqH2xWipXEzQiXU4wue6uTM
wmHVVY7Ufo1jLbwCzNOmHRfYwnpB4i1ei6ki1oKAwVFq6QwZIzqQjuqseb8k5TNpNRXp6JhDeBb9
Pt+ZEQb8Ghz4haKrDxTdPq+lADo9nnMCqqi0b0N40to82BUqPYReVSGNGH/NoeZvGXc4om7UMKPM
cminikAlbrKvT3Gr8lV7ANBjzhR2P7H8t9xfdKvwOXxT27H2IqUMcbs81Cko2ekRAXHwv0zZpfEA
cZUurJBYEvS40neu29OzHoB36Q++krYF9y/vWi+gdwE3NkkGknt7wa8vqMPGTr2UqhhrFJsY78W1
5U+xheJENCyuPSp7lsDstweJWfCKyFvkLBVXNMX/XAq7OIDQhXF9JUIa473uwW5DGUS8RnYR2EJm
neRyr2QaiGqkwQ5hSElVkREcyKmAcS69KOikXHejp7SHRchN++TRcCBLveOyp86ZHPUp70LZy/+A
yGnRhCKH0uTlctPNtBwGQ6oDp1UmOmWGD6mpWd+CtlTeHG8cuL2lApjKgEebXQ/NXHRDkqCFqBcJ
V9f/MsfZqRsCGbjLALdT0uv3HfUA+ITr1jEXRAWiN51yHQpIhtv2T5xng9ofK0D5Pgg34QrY483X
U0/DqrPYpSe7ihShotQp8Uo8On7QpB8nZKro+0QqW53bh+Y0RJISHbN/ZEKRB1vRcN0O4xGjKNeQ
iwTCwR366u5SjU6c/2I+ycOg/imi2QwpVR7KcVRFXzI8BWRT5ywYcMmNVb0Vbl4PPo9V7j9hKI6A
00DeU8AnSL49j1Er+q8F4vDab3RMhD5/0970bWzA3C9Gha8GtaNQdFjhACuIy1cJvrTarFt2yoqb
NnvXofIX++8nhhoSa7RYt9qaLYGobGa1sEUoQSrQb0TNLdkW5u0Wt2I8OAf4EtuXJjypAdF+fAzB
2hDOTDIDCyGsMcm2gyln0JfVwUmcrg/OjerWtD7R024tE4Fhf/t4HkQSCkOohDMEEqo5y7J4UtAH
U8ro+LtxtQ9FzjMWn5CAnuY6RhLrs9hv69ko9ClTvEA0Tth9JwOnCk6G86cCFQ5oco+cIIr759i0
gsW4XYCxEuJ3sUdgd0YFepcmkwS/2I1JuaQ96wuWi1+VBlg1DtpqaqFx0O0eOWu/S57QK8FO51gM
5fKYG7oTvh1se389aU0OZMPL8LOUHHkZJJhQsVi70F0/DtC+gTEPE/xZVqQHLT1nCAd0T4LaQfrg
nxAnHlFYTZz+kGMVJ9M5dAaKVO9SmKOTj3VhBM/GpsuyudUhvvEDjHIvU7I1v30ceD7Xzg4WchaQ
QqQcs2nSlYYQ6MlWjp+3wiE5lt1a7m40/irdnUHhh11aeQALTO55GGPsdyGE94yl6zqam8Lf9dY9
eBN451MDy9FX63mVRvJrPlASPR9dS+72mePA7c8OkW5R6CBYrp7vySk/w/9sZKwBVr6PU20Sps7c
18eBB6VKLzy3byLsiOvbuS3fohCNZ4J4g7ZeX3hSBV0x33NEkCMD4cZlCnDaWW1N/0c4/zFjvhro
59FociKFLW9ishh9TEeJrKuAy7naAQMFl70nrxiYljBYbCC6AnbCJXJyE0KxPpjFeFGW+ssJz4lS
aFqsHxjB8w5yr/DIzwxP4iysdjO/FzMmUs2T/dTiLuj2vVhHpH8QFrPE+2JDojn0IsA98WGwIvLX
DEdNxuKoA7KpOhQLXsupWc2HzhAyu+5k9tt5M1g9VImxjJSA4+ufdPb07RdBE2usW5FkI3nmOEtI
24VY6P5dYAuf8l25LMqHwxeZHiDy2Fpl1r260duSGGDHU3Zxfet3MfFRz5xRCOt62tZpnETSyxvq
n0mSkOwQNC5LUb0yxBHnHGy96ZbYbpz75p34jGG6EaUHplYtEAUTI2bpIkQf+GiJuZOCexOs5iBg
Inj6OCwE6ZKRUIHDMicZF+7YKUrwLnnVpvP4d8TeRyEr26YbapSYO/6T1J2cfNATj/tP0+B5fidr
tzKVtg8dkdi2u+R/GgWPQ0W1nRcl3fdFloi7pcZbejKmS7JOX4WZAPK2sQyeASByfDrssiVgERmg
fEovw6uNryRwh05r+BIg6x2/MxFtI1nCoh+1W54DNIFICgMbv+7zRSTd04AdpSpYiQd0VgpRZHD3
a8qjboTmAw+JutHDQ1wmydlc6n3r+Id21Rdd+dHtgW2unRBoAdHbePpXYbrh/44Z3TY7WveFuSYe
TeqkLNHaMrShmLnv3FAPKYL0Nfqf4ns7hHI/An7SjJ5jqd36gOTFyHSdIKbY1szddA4EGtX1FpUB
ALaFKV/T9UzMaKgm0Ne5AXTHdTaKhge/CQNh2k2BmH5NbtNnY/3L1iBUOcEH6Yq2K1oHv7FiYB8Q
GsZSzoukJUL0WmnEvyyGgbGIxsbJ80GiIFx5AEPtn3TlwPPycRVHxEV0kz6fe6+PlFAtTBqwk1gc
hlgNy9qXu92Rhqo/lr+afUhCFD2z5UHZfoev1R62Dm/t0X2mQLNVCw8KWRAK+CToDfJNZUp4H6g8
ti2kPM8mDuCQzg67Oiux+Oa0kZ0ForPWMyEz04LHkoqnK8M7iNfliGWO6PHoWyuLFqpRGyIyI6nd
ZO15qHOmpxUKZ3noE+kpw2lwv+2PaE4T6PZ4w9OzqLVHD1jKvgusyn1vO9o4R9QfljlnABpiF2BA
kc/Cafdmqxmvx5rWJFTkhPyGrp8WOWP1nRV5hGzXkQqqhavIHKNYfTZBQS6xNni0dGCQmrXScJCx
HITgccfN4fIEnePemGluUJcx/9MGBOtF9MNFfmPODyqHovWSQ2R86CwyakoCwRXdsdIXjk1xBCxp
ko0Z4IW7LcQoXCROe/JpG7nU9wo0t2z2Jobo04t84zF6fjwjXH4PTdP0HVYUEi6iIQbg94JrU/b5
MuBBAhTmqEjRPaUQ7/y1y141qNkR9KPyrZHz5QxisimKPvy/jBuzP8YsJvySUQ1y/ZOQ03sTU0Eb
L60+mZvHiBk6/Eh+5AG2vEhuYi8ZRqXxieZ0ugn69g/WN+Blu0edvtGQKVxha6SBiIS6vnzimKof
a6+DRbebiWxcKhuNbKqPejZ4FHQPje3z5LS6RJdwNJeoLt+fSPDnt1zHPLYi2S9iaIAPqq6rWNUt
qr5E3UcQR7npXwoe5o5XYgsEvLjma+hEBtj3S1VuEtmlmykQTNdsROI+tPfkofWrGQYiCg9QdYh0
ghLZ5aZxZ1nAj8GDY9Vq/Z9O+m3khl60WkcmZxjwUshIewLupbw+zgwJ1kkGOym9Qwx0i4RFi9z5
x5olcM6/2Uoajc9kiYqo98WJE16FG4MFrPDUkE1gE8kcXO0/pXrEc+86S6flgwqeuqTi4UFtdGb+
oEFPOgQT73lX/Ad+9l/2GVK+6ectlQUPgtsbBg+tmkazKCCDgQkgKqLYeKQu05xjKberjNxcwIjb
0p+AAWRqNKUZgWUW0scY7oiVmLoVPVXGxmUlb2DxIs/0NOY+/0UDkE8fdKmu4OIEjQEE+S/KQ3kL
K8LGbhAShqK/J6YgNzxUf6H96mvVU09LtGWZB1zQ0qxorLRQo+o9n7gTU6Eog2KbyxnBJfmct33H
O1Uj6I4vWCkOb8pDtiNOm6HDX04Kg1pNjX6IwsqMjyTYYp4eP29Tl1K5D8JqEEOLP2DTtQrVuYc5
sB9Ag9Z8diPuOjvNNcEVxIb8Fqaymm621RSvn3+Xw5dIuGTZAFqMnA8koX6rJnJOD9Z4f6gMC4gQ
mLxAicIjPuyjaWubmfQyifMf1EYUvDG6uCi1S94VvM/svDWerchN+fWZny3w3XpqZKXdp6luamSm
NGegtVG+G40atBItfganRaWROWNW6FYASw69LgbmfpGMBAWT1xd7amVeHogHkEKNyBEVIZmJrfRw
Oil0Bb4dg/sVmqh3GtxITgq3eHQiVS9hyiSaGoEFln23gaahaVydSRnh51qQCZZ2DN4ngu9W10V+
3GVTHcgU7sz2GfEJwALt7MQWnF7iMKZUU0N7OrEU/HJ2kv90+ENtTg7R9Ccr6ixRw+Dg0hbT68CZ
q+b5GbUg5JJHpBYGCZG1WWMo13BXEiGsWuDPbzfxrgGilNS9tQOjkK7AxX6/dG9gdTxbS9kUObHZ
UG6EDpDLhFo3Vfdra/EsRf1kg0TeTxSZWGjzYk+ILhFxIj+ENLZpnNrKkJWKIqrIKh/9gpAOCKMP
Cu7PNfFxwwqpE7f83vuJGaBWkfErc/qpg3A+VmMXKRdjJeDAJL7wzvs6loKNU7rnaZWZzq+LEkMy
hrl6/LvevxwtCaQM+9NCJiWIQ4WhwEFDcnDzWg4rYEy4WUh92zrPAF0jSdTrLMpBY2KW4xKw4gQa
BpxePs+VCWyilqKXAMgeudpjPjvRDWJ3dw1dzF7e3D5OHPazYO44xlIIw7+18YaRIH5+B4LPTpBU
noBJaDaIPIylN4xJ58j5JzcDxrmSEd1DWZOkrvQXKOlIBHzVLZYWp163KO0yvyp1a9x23ojbXv4B
G4dRy+rfVvBbg+XDblGjwetbUKmZKqiNmesobUjYpI/fOLzYVaO4I+jFlxjW8Psd6MmcxVLczJeK
5sKZlyhO236fdVTvtwrXPndF/nDMmq/lDpkn+WSt9DWr7c8a57cHW3VCi5mIKEAbwuBM1VGcHHDt
4nW3eKo5JwxFVAsmNbrRmylSTWkQIlyof1TzWIiH0OHqYPLoq+qlXtxDuMwAXu2F09Lhom0cMx8S
BzZpitbwlnCgl4GOxH/cNdquCDpogt67NlBkprl+qYae3QLSSzhNkAto6Bwz3LcP60jp8YVp9W1S
3S8HmdITclB+8f7cg/Wwhx/C9KAJ+LBzbRx7aq38TEOrqqT7OYuNbDPe8TfkX1YYsIsw1FgOzz7g
O5eL0OBKEXGRC4OfrdB5T79wRsSdr0+1Kqs4cLXWFHR6353d9LUhO6OZDxY1S83KHt2YGPqthhYB
JsjK5xQXiPqV9jp2mscar6IZtlHcW11seaQXkA8wAtMxLaDwuSQ6DvceGGxgtPWPx7TU90aWbtfE
act1a1kTi0RiLTLqjqnBDzYRb7D3WlV2e1USB0Jqj++oFtGqPLWSenQTfPOEXU3wd1i1CXV1NwOL
i/hYPYRWHZEe9kx3KOGmmAMPX8QNlZntVS9Tr6vxD68/dsTez2k5+awtTVacr6eb5n1xw32Yo91x
MIIEzMED2J/xXj6Eoe+xn488V9efc3WNIW/sARLs+cACKUaDfclQDZD2JVjuPvVjLCxRlG1DAMFt
NbsQFQfwDVQEsmipFZqQnBd4UpGiFtie7mPGM0Km/itXmiJtUV1orlQC6c4yUAKZal0/Apd1HclG
hOz1dMW3E77F9Cd0DxJ3C0AbHvKt69+BXvt1xL86x4Is1rJpJV3J8fqFIz6oDTA+UUY8ShupMo60
QXkQbp6fOMVc28uYZdZqNxjOoY0zje1qzmASmz82XBKfgsybM+twpIj9OcD+GCTSrjUobYayMb+Y
YUF+8G1eicp2yUyMDoAO/Pxga01ZQQ/LPVZ7zoB1JTtKLf0dsd4eOdNKsOfPC6s6su9jPyiROfsU
lf0znz2A23hTTDwoB+Nv5duCKBS89nackwpnQa8HdXHe410lsH2lGwjGJsNkBnxAOlXAd38QUwWV
Dc+/ubr/PGv5w8D2fO5VWye+FrEbNaum4H6Px9rcR1+KJfb5W7eshTCS9tzQu1l9YD8efCVqj6RY
87MM3hfqhjbNQHKZ7Z+ihWsJ961pVdzGbsoxaYyXt8N7/h4YNXrKtVgINZ6Z7tulnsl6BTJYJFEc
gBWOto0h8NvUztd1fNR/j+H04qAqg+l7UkLAyEDm0OpHztIVuRH0Ez8I59lO0Gmm+kRsLZEE8j0F
4hMkLllHpA/yND7gXc8T1uNz33NAQGBUt2RG/ECJDTF0xETrIUyNoh7NkVGjeBQkijwBGKMq8epi
bnvZA3IJ6J0SSvuwD1OOuxqleDww1qfH85I9RJfsriKLXP/VA2eXmbjxrd4mZ3SJ4NVGpppz9vnG
BRodbf/BgiROrbbSbwwqwgzhujwLlYRjL2TD1vH1tHmKF/CV+ZJfHhrdoWACA3dvR5YR/YKgF1dE
bQGlUe6igcg5JSKoCWQBMuWM6uI9m+a5EIFpo3J+bRQ02yC9pTj4V6yuEq+3xR7AoSuK6Wdf9l//
TPRaUKCseUpcEdNoinb8Ec/o3Uh3DhSyjH3nY0O000UVSoHjYJvAqHpt371EHHP2qhqnn2mKErOH
7xToKNBE31zsqzuTJqNjp5yJc0WWddlvQwtEyIKSUzIMbkQTWClUCj8CO4dzT6ZX5e02oC/D5+un
9vyV1j9b11jDGvB+9h+tpxUe7O/IYze2jupD9CBiq9UMrUfGJnli68DFJlFmo6ExlgIhHm1dGXtg
WfYhJF4RXNIWYA2skVTfIEg7lj31B921123FZ9/OP+BZs4DSMjcWrzcugBxo83gdCNV5FWTwOpXL
KqQYhfLe619t6amfTIyrBomQQyHtYciK7MXu8aR0VRkUisubwFV6sW9LVUa2n/Rbm2rexvfoHjrx
d918xg03wRwg9V4QF51Ls1bdnHAuU5oF1sw+0q5KuMj/FdixvKrD4cvObgG/7iFSY/4dOBFi/lGK
O3Ok+wdgBzHfcYQVdDYwKeqjLhQDCnhvozxk/hVLeOF8p9TTFbi9BQJSW7coRbT5++olzUezaPqX
dkKyqcGOKphTA0+1zrhq1h6oJjYGHh5UUYotXOW8EtlfNtVv0onHgDYkoM65V8ZPIND11xZN39DN
RxI2tGseh3fdF+064+UU/6e4FtUL28OEVh6XekzY1Ar4jKmbsNa1bnCNx8TGKa6CF+z3LwbdgNwt
AbjjmDK0kAE4QjVRqe/I6t1/otlqbOO9JMxckjMSugI5lXC9LBnAb8LATTV1MGVhR9V6NrE7vll9
NORCC3UtQ6JZrf0hSQR+J6x1BZl0Z7+FyTSLVCDMMfpKdBlu+9MuIIWTzb/Aqiw2FTqHtG1sA31T
Bshquv7CW3Z0k0C0DtI9c+DbzOGYx3nYTDj7l+pwYmGUjtlLgIQm3mEYd+bzuuf1nRxaI5Zwiv6G
hYwuI+SsDfutTaRTTcnVFB2blIaucjOhbXYn2VEvqhzKCYmB9X5wcwkZzX4Te3In6R2cddKnym/8
WRe24c2vTcasC3SaQuPhh6sLC2vDCPrS4E7eyWENjYXBq3d3OWJd31ohGcVJCIabTTGk2SbS6NrJ
nM4ds4Hst2HgxW0BfgjWn6yKubBBJIkrvwPLnpINQj8WLr/LpmLhVGxO8o1BTEveuuEtd9npxDCU
MwLbp4CJXL5jfh3R1r1Zweiev6zqLy3+7JjM1u2vhtF8mbmwGzUDQjjhhIP2xxgHX16/b3qpMdhM
d1j7ggeibxctkG0j8+iJriYdiA80dC+ZaTW3D+EPLAEbLs2Q0Da4CZ3VpGvjdJWvP/WMJ3ZnlvfL
x5X7b6V2wSPVfpxzV4iE5UTBx3R91T5D7pVSRQsnX8KTM3NKVnulsg1tvaYs9p0KTOl590bLR8mo
tAMtzE0843ue4qYaMo2qzJRf8I0uYFo4y0fIwG6Gf9GiHO+9sfVKFanrtJ4knKUCmbI2qIe0BAmn
PFi3kVOP5baQsf+9aQ0cQvEfR3pAflwOHX6HmDWejDOW5o5VnsJb+CgYNjkAjc6F4zRLLPq1nvTy
HaayAMSKPwYINmkwidvttoGXFCyUWh39dIVBDpnJXTgHOeADKW+Mdp6W2qiiD7mWCUd5zgktnCiY
SThPLaLTVoClwfYSlbmtckdyF9fchcpGgYdwmXoko2XbovjiL369v1XsmjurdxcT3nhwbYFNFcNn
49pNzUX9sf/q6Po4YbsAmLXkYtrAV/JR2ColWMOGZCT6pS5y4sjurLZNAizHNOhHGP+jvvaLLNaE
r59QLPA9/YT34NI4/MuYyQCIpg097w6ZtbKO2vPtWtgDscS6zHM3iS2PX9eoMjomInW/TowfybA8
hocByMD9FFFkCXe9PiaO9joBEZ8bujgXOjcO/DPe0nfnnDsgPFJtRXFev5KeXsakw6SelgjUqWX+
fqr7E7pZEx1x/4MPJhioMQLLh/pCM+MXHjcUf2V6Qqut8AUFpScw9+rKzVHy1eSmOSLmOUN9T45A
0DQDtDxXdxyLjHp8xMrfPKmys6/yCu+1EE09o6OFW9OrELJg0XI20nf4nZP3mMOdEqC0Hbqyv3gz
y0C6LRQp4Eeikstvbr1P8YKQi2VRftXt+YbxIV/Qt1IOEAWIYEMyzQtKehJuxVtsTDe2w0sSmFMo
i3EtB2Fl+fA9iXdUe79VFU+g2LEB3X/ZpKPn2kyY9OeIWSRavDrYR8ALASdjZn/445NoRou6j4rT
INOYpOyZb0Oy8+JgzGqCP6JIeraN2tFDBqb+64MpAJl61TCtbE/fzT0zuHzX+fhWk07HZDIulzB1
46f2hx8l8Af1JI5/FlqVHPeCZpbaWIAP2UUEVRwlsJwxX2eH6pUIV55knOEvpHBXqMhFOB4vXltc
EYcIg8gVDhvb20owjXUb1eQu6BP7vEupEglCrlkekW2pWGVZ4k1NUA4CppmM+vK4HxXZ8dwKSPbD
2Jp3j6/4RuI1lvAdBXUEp9c04CgffwSe9Dnd905G+C0QROjKd2HTptJQ/+7CuI96qf/05IQ/3NvP
z3fwYxczOUrQKmdXhgbSaXs2PJ2eoRQq3JduFEj79f6UZvOQJ8yZTrGl4gUpKl5wrRHG7NG8yN0L
01l+X6Rg/Z+v0DitGXWYVu/S/s8U+NL5wXRsSPCdxU1bZYTLE4cC7ccHc6MehAyhO5RlAgz/92uV
YVjWAO3LkIgm/02saKufGb7svUklVZHgeA82h5gd/CSB6pfqo5M9CGa7Y/hlLDk6U7sUiiJMa2CX
FhNsmoPxKaPLyiHh0ZrMMOZmKIyHrbTnUb4wUHLBuznpKhP8etIftTh0aAJ2L3EEb+xTlCjn5hEa
n+KJlw0bC4p8stiiODFV6JXzJIKT8k4mro8t0ELx2atuxZsLtl5XG88DWFegZsqRFzmkJZw52JHk
n5kOskDkQkE601Q1s+opAGYanVhOJiBe6V6XxGBhNbvSNzJ5u6G/a+4w0omrZWGj/1anvdCb9rjm
osOhZYRAPOe/ga8HwnZZLHzaCKubzQRkWuvuG+aTg88m55VlQ19GPtZINGJI7ipySuR4XKngRyvi
AyQyuIUi/P7ONafDWsclvntlNfvE7GSjV8c2zy+dH9tDxIgdsXMZgmauGt0ZNKU66UOOwFc22XpE
2+Hsg/zdLRrPRJ4qDjweDasVLqaYL6B5rsxd2Ytfzm5BrgVZtqOcte7EkFesluEGTtyQ9dvsbupC
wvyPClVezEOQhRR+1hZTfkllro2xvivYBIZ32nzuNYlIYfGmhk/EvpEdox8JlLH8kYYrvEzh/yWt
hYyKSVamnPl0wutqolceX5Brw6diE26uMomoFmE3zHXaklFi3ALZ8c08/eAefgBf38XHBLdn7uNJ
RjMbzRUtNlBHnB33TDfmmyo4yWzY2+FNTg3SlXO2y8tq3FeXJFzl0hTlbJ9n4uxTtCIT7/3M3fO7
Qd1OQgtyoT+/QcFGzReOG3V7hNqyKNM5S/F6WG3dWp2F2EY6ACSVqwjXUWgNQ9xXKMbeFdkNno0l
VDnz70rNotD+wbT/kREEPAv1InNcuX7krwWzkOcIfHp5tZphXbOmnxOa926wM6qGDzajAIp84mo6
Qq9GYhfABhyLGQcHi+E0FdSSdUTmeBVNn1ayqbmGeOssfrS6tOsDZWY0iCcuMq8X56q/0FAAx5BD
Xemh1sA3iRzPdo8Y8Y2si5WGLf0ol6eEuQoR7fnrDsLMYOKV2AC6tRirXRLzASgJrq2ku/Szv1Wv
97G1n2b/iZ9TXP77rJYgnAyb75Am8UxLKnJPGf8uq0TFRZsEJy0pE1jMM1vlKeviEdRFmHfvu1Yw
6/AGZpFb5Xm/t4o9xwZhbD4fpMQA4wLHDCUKz1n9vuGP+wrB6IuNKdpkK3R1wl467FDNfh8/vHE1
FSRnnZKGtjb7lM2Jw/sWiKmd+U5s4UvC5BRMdOKXTXOtn2LJ6bhbjjd8SwF0ekmh7s6TZL5xwDhs
26/XCL+dKul9HPBqTZDIRgmpDqkXW/PhmrFQ+91XGwxwuQRxTGC1tEAZg4axBE+YqOWosRP4QGyt
lzrjGwxp9Qf+3kzZvgzIhKIKxI5jgxVvt3uKmQ5RKBNdXzJdhXVXNk9Y/nJPjNfwPO/SgxarFX1y
pW4LSiMNaqMI++GHULSDdQwCW3jecNWwEoz7V+b/T621Fnqi6Da0OR2znPsSTj5ubIiBhI/8yXVw
nhVkF5uQjzmnsjyqfR4HKvV+2yH7DbJz4/4mTPk6t/yDyJjSa6/+ArjCQPblStPOQdw9aguYi4vv
B21jeGis2PAizzQFDRl5nzw1fZNTigZ1U5HaY6xKj7wvWESn4+Nb4uaO2HMNdzRbY5+nsg2+Ub+y
gnIyy4253DomhDDYMYlPiOSK5g2Jm3PJTGZBGWfuZdJ9SAsS1fpTo6KEGDHMJeTc0/u3Y5f6kwKX
7pp5/JrDJlcraxtnzOJAia/+kHwN93PHPZkGD5YVURXiVlz0NiO6Ul3BMAoe9/N5JFnrLCZG/1JV
d+U3gWKIpT/3xWBGTG5Yi9op/VCnIWsohSbZ7vMq0c5+yRXgywcHOXLD6LHFKtckiivNzGIUgbuw
ksfik8LHOsjhmB9H/BfwTX3JEkyMHcz0LHdufd5haV+UZVpZob6yDiNnvUIPohKnMSTS3LkkB2YI
s1fqyBECPBoJq8u8FOuI47qYkhwKXJgspn5UWMAuUIKn/uHRJGOAJMgC/QmX0CrGBSHTlJPbc6YE
l4nzaza8wxYOgUXZw0QiModPAbSW7xKXeYPBxT4Sog8SCxuuXRdgptCvFtIh878HxiZ0XO8Ncjuv
VKirXbveId40R6YehuOxWsbz6j+bf4QY6E73MSaVO2FQFeFdzyGL/0vjnWFTVFfPZT7G9fP1zF6a
8Quii1XQ+74ZHOH/BshrqEu8GBXQWkMAd+4MBBORcXwQ2BXtOI72Rd57yPed1WZGW9TpYd2f8FBr
DZJ+vpgtDamlvsETWKenLfi7Z5RcZFt8BRY4wWmsGGGRDVsPYx1eeURD++J6LcR56cw5vhvJjejy
/bLUvOfAjGjrkS8JZI5q1TN8Myd7K4ci0spfplaUFuVL8v34ONnspBQG1NustJPx5acXh1LdKDw7
YEdWPft+IIs/JE8y1rpLoTn7o/kxd9hqSbegTJ3KE2tAkzQX8Xgebp3NRaulXC3houNG5pTo+6nz
oGaIqpTeOPn2T71UGYOsicfDxVF66PB+TbgtjlDi8lzuk5/iWeyRgtXQZDKMz7JQF3nrBuNihkwg
zOUrrhWnoXZnsa2r4djlxEIO6zl5IgBIRrbVhMz8hwjE8Hv++2BTEuGhHZ29hvw3V8z5r7JIBq7G
4/BWQZljEnjV9XhIqTwTydkJN5bwVoDJ1Db4LZkHy5EigyiQbIgL2jPPZpN1ZG42xXBv7j/mBHcz
v2OqZYETbWWgic3eu8Y0hfvWk/TPI1JqCRVONlMjkXJBEgzbXBe0aTuVhfByyVO6ui5K7oOC3gEB
myMKz8RRpJzjMFXyNH10sEv5rP41Bh5Y2JmxWzsUaaiva30PhZns3DOSiYsHcAxrO0VonDbKhg5Z
M2Fld3Ki91aQ3acuhTiuUMitdB5rWKxVud/1KQUm/6llFBdJ5lcD2K14Ow0GFvTG6bE8/4LRIvab
60+c1OXHG2iYloKMQ8S5r9eOFOgVaSYISznytBH6jHelmD4JVTuo9jdBpjTlHx1w7RgTQH2HxO4Z
iHzpQlzNThojFAKexBi9aqy70khS6ttF5W/xFEaFDP2FORz2GDkDjxN3YZL8yp2ioCgcAVEwPm7g
uP5jLElfx5UcamEdLmACdq6K+kzSWRKet1vFj3nwonw99vDo1jAlHKkUVvWGO3NqbdXzx+dAbjS4
TdLhb4iuusGPVlr+bUAbsA/QwTJm/QCRWVW1G9ffYy/mn3WvM6RaQpk4NlYDgRUtqxrecN86gDS0
cvtVlSNUcFVmuc2iaWj4+DeCrK/QZpjmr/vp8pEbUGYFn1QTeQ6FvN/p0gkeElafAyCC1CRl3nKU
sL6dgTgxRLZA4N9Au1ZgEv7iPoswpfAWcQbVhHTcoh/ELryK0Mj6ODo2Ki2DMYwz1xA1qUEVFBJV
RSxpDMMQxNKJHhIncX45K8eu16qJ3iJAAg+DGbL6UVaEhODLShcvXnzFXDysbIrxWzdShWhE3x6p
1vn1+pGmEgesqYZSCUZVYpEwc2Xi61lu+SULUgEVHeeMV5PsYiJudanebzS02soFwicDMpv8Zgrq
vKC6Y5frtbIPStEn9oDXc0PWlTDNorsNZwPRBgHxyepEQkQLPviH+DJmOwL7KJXyhjzffixV5H9z
skAYHl0o+A36chc7WSFnSCxmTXX04o7Qc1wGVT9Be1tAS4+JEqlTTduvmiHTP5iDVv9/efYObcy3
6vljLkR3IrWB2mZBvkhyS6b1VWSA6kAV74Q8h37hkVNTX1Xm7/Dz6QCxy1Mc9H5wSKl247G4O6al
ku29mpGQFa/he6CHovGHqJkrHK/QExQbq+IvEXhsqSv8dbVliVZbCTuJOiTRzWGH5Rx4TwlZ3AFg
qycn5sI+AQZWqcFWj6tpEa95uruajVhoEsVsFEvx78gB7EYPwSNKid+vInKM/TVeO6uP1u0rXRmw
9HA6UbXZaQDnv5tEBFNQyzcCrflfHP+wvCYYXMoA11MllN4UNDEAHqdzmob6HmFG9/MRpfiGC3dM
amN5l2dcRt5DJ3EuR+rpHvrvcww+rl5qrAD7fRH15ugLl5t8CuFiyO7p3DngOJQWezlf1h1a9Q7D
wTKCwrCoiYSNL9J5BtiCCqKe5WufTP6eoI0hHQJ1O9xPtp9V8iQd8+73e4EsFFlyFKYC2etMDvHX
V3gPg5TvEllGbsUAh2hJ99qQNm2gmwr/OD3F0ozNh6UeO9PNA+cG74r0crsCKrTIK81H0Magsnkk
Xh5yFddaudgddJsrhV9mbFANjIwGtpyzd4M6jOCAyT//uEvcFJxG/2p67N7w4ragDV2HaVHLrlhl
/RjI35D6Is8buX0jQda7fszYV/sEe15ke4ks3cqz+d7y1dGBBh+My6o1701RDDwCLJKucea6A5YG
BwjB7bEmtuib44SKpY5wZhJfMi4+Fb1dfsei1Xqm9HVNvkXGHKngeBya3bVPSeDr0L1Gxn73Z+7I
G5S1yHK9FyJEn5e41w6hrH6ZEf/8//5uHe42/10sdSGm2fLzfAoYWN91BojfaNAS13C+7zLLLjDG
VaArCrgdeQMSKcQdXn1ws/RcWeLGTDWYmY5ttzrFpYCk9us/Tdlr0874P1S8xtPMhnE1cTfUzys0
qtmvEgjzeiV25KcItqmfy4ITK62ltrkp93yRL3+riij/RpxEQHRcmD/UGEoN9yMGTDPr2lriaW8/
vdARwVmynzS/IbutevcQQHD4iZcpLIVJ431s6CMnQldusDm+mrB32AyJeZS2G3VSVWGPXQ7zmha2
ccUMfHKDyckDbjoiWmXeGmBcLry0PoXYry1ILpa/7RRWr1My90Z2YSPpThEoK3aQL7GtP/CTY1AO
fsk7EN3Twjj53miBmgWAxqHRf9TSUrOzuaDXW0sK8LThYisRlEbVBcevVELCsPxS/RWiPbNZ9zyj
4GOAiPvtgYegl4yRhZEat1sMY7DlbByujsVRCV9MnrtQyI8DwV+GnJQ6kDOI7J5vnLo5Iw/LDYBC
XhgKjI3ffHqakiPcYJhqrFl8twD41VzKAXWOTK573C7L06bIOEZ+Gjup1igod1C6OfhTSB46RGT0
MkO8zAfGiPprxWirdTAozdcrnS4YD6tJy/zpTMI4hsiEb3AWWt/b8Y+J/nTbmtxiGPQMSnO5i6q5
nWAWuC0FWKnywWnQP5YbZqX5aDwbl98hxQDOrNmVXGWdFKpj/tNF/IqTj+oOTCHffW0UvDKE9zz4
85hzJYymvvyeEW1oy1FZpH4PmkRLM/SWq14Z+6pFX/lAxIggbs82zFYssXwUmty2XcfW2g4kSx5G
3m72ycPfoyAl04+DFnyvW4wiNgR2U7zhDSYRxPxPZVCfyaUPZOUlKc5sGJiYyM5N5IHpuY5eqsKX
QnlVgtB5/AzRv4X48K1a0FJyz9RkcY6ZfhbfmasA8GODQf7tBa84xCiNNJc/BXWZ68tINH/GKTMB
5JI8Q0MnFhyxKC3XdTLpxc5xrUdq1Xcur8S1ZMEbfEE2v5qSzPsr/RgUI6ffo5DjABGnZ+ssG556
OVuthVlHxKC/xEDtA/8/kSk57nwS/WFLJbNRFhA6zNntUu71v2do05vxpHoWRqRKcLNVho20SoDk
lygI/J6mBWZuHQG0WZnPyXoG8rsfJscdjF/wFMv/sgV7Wc7zbvNmv0i3QFcMqNl0z5Fp/SDpvqnV
R1SsE5G4zybVWY+XLb7neL3UiCDf+pPn3TQ/pCtyqHKzlp2Cc19c8lbXCXIQPJPY32ch8ckG9pb3
jCRPNqv2DjWixjla14QtscNbzsuf3sT33/Xg66CPQeo28dT3OP8aJmp45QpC6fgjlbnfKGReqz1m
A9aebIugESCMMYcAs22Pgoh5G8wz3ReuCxbfWGf1LBmvGd5BBfigC5+67zW0VslajceLofM5QzqI
syuuFqjnB+Fx+N4oLlK52BkaYKeQhU3fIbNjkeW80czQv2a4SnWxj8Me/U95KePN3d7Uhgw6R1s9
0qe4JFAO3lNIXBwe7Caouc13iNF+A3H5acsvd/mtyEA9CKlu8OjO3e7OrM9GAJnF8z5figab50Xq
faF7n2jw3MWIC5y8utQ4JhGcj0RGOtM1foMCNX7oRJESwZsljxidMfni3cb/Rq9Utm5FICKwdnek
ZvSZZCD5QuM2c6apFh60DReCaK/9ILKeg6tlgv0Li+YCDIfo7QL/LJBfj0G61OmdpnIRUVSY4mv7
y8uQuxtHX+/5kcj2hG4BZl1EkG9v0ndpdVALbHv6wySCQjWhnGRwHyl3D4V92tB9Ug4d3hkBFAwT
99qhshRPFzi6et4+S0WoeWwJ03eAoeLTXquNCO5g0s9XDuheYkppVrEDAEd/FJK5wvXy4rnZmOpE
S/bpxuNfeK80MS4uS+icw+CV0LDvDN1nsLMkYCNNfNLuIYWDR5ysbElUZ9ITkL7LjJhAzWfGuzFY
PEfjMQCJmVkBdHhnT5giQEV8ZECVbB0el0m3dT3YN5NB2FmiXt/Yf3gn17wecc9kPqd1rqH78R9h
HW/PvmFcekwNee+FyJPNqvF53U+4tVGgLje3tjGsRR/3RVsTquSrn8LVj+R4TtZtPtZd53Xcfvz8
95g6OMR/FOJukOFJUunoVVV/4X/5abVVsrOXq2vURnQESzHOf5IrKTT+vUSPKqnnBmsKSx1VwunI
4wxIVGu6BT+mEVm8ZDWJE1zomSklgQ8kJXHFku4V+snAVz9pyAediUtwvPkAmpXou76zBowtuxTe
GFsdZwxPaYouWTV/QRCm4e7PmMhnyO4qz8BnzwOA7rIqqmIL91XffqMncvRPKJ1QEQLNzvwX6YXP
jqD/a3Tmxx3KHmA8IDRKZ1ksH27KfIfcKK5cVDXv2McpnBekRCzpzNdpVE7pNxz9vPrr/QSbKiVE
PfaW/gGP6rLf7ByMHpPR2ADRcHrmV873B8eEo2W7PTxpn+yxX2IiKXqRtlKPoI5mJQVxj1EOgusP
aC1s1BDQsKk3agjseI1wDCGFXGEDrEUNCeZRqKK+uuVL4sbypJgr8UAlOwRdAg88eTbeK7LOY1V5
2k1FIP57qFE/wK1Eboivk8egQAg6s7oJOO+kXLiAAgkRz+bC2eUXc8Bm5y+48m67GpbmZt64sTiq
/PwJN/KsnJPqvLqZuWYLS581jHRANJZ8kQLevgusjiNxAp+uvWrz/GiLZoqkD+UIIjzApkn8NnZ4
ji0kx8XADolWM0QfL1gz4RlxhdzeSRUoI7yvvAfaW5ficUpbF9YtArg2QDCaittFfiz5CIUJxjjZ
Wjt75oK8fD1ajXgjYOQJPivRa/99MWPE+1DbuxU8sY8BupeEzUJW57CtjtVy6bMVACqYbRIXy8FG
MnumYpwk/xsoU0fcUtxvtH36pouAq1KpJZrwkvjgkzYOAmrBUttunhP1ng6E8gCz3V1WWqMGA5pY
RQsEInIV8W1EmOhF1cPUExeSjt/SN+38lIWDF2EbVFyLJPQnKRwzxbl9JC+FC0VzASY0+Rgkt6qY
c/V92tzL7J+KQ0ezR0PAPkieSzacAVaAC/HxmJrvG1wo6TfpoHV6Fw0S1D6fJ6D48MqXJihWla+C
6EzfZ72+N8WTIaUGdY90NhYu83rIQ3RuFhC4wHUyBOQOi4m4eSxwFUI5q/Almqq5ptqZjb6gQtrM
xg1P2eAWoCY4SoGYdpUCRkZqxRR6QR2kKglHvFICvRNTTheo+X7x5G8byu7HLd2wwhmWwMiYcBIR
NqnlRybQhOpLzr4UrrNfP0JcGvc/LYkn/bQa/MtELRU/4Sg3s1vE3guK5FAgyavu8UP7TA+N1Lyn
gI3K9JQw05Cm5BdTUQVDbyT5DF9fxcNwkOxxZhFLvi5+LQucRnCq3Qr5lyJfylkcSuuGpzzuAbPT
oIR2hTy3JaYodBRA1a14w24i3lf2Cx028kCRiC2BDii70VHgGhyXD6NFkLDTMJoSRRXfs4w5aM9j
kwxh+F8CyoPJkE7kuSHIhwQQt9AmmCE3LAmS/8uQhlnwfnh6f5f8PFqQ7p22gpNgnzAvZDq2Nbn3
vzQtpA3+hpc18UiJG4dqjzZMKL6PmqdcC2Uppbx3c5CHMy2HAoJZMWd9wE0e4lu4WOJ8t3Zm94+G
RGijIvkzMe1wfOkYaRtaqzTZGcgEMH4V0XLh/fRMKtLw05r0sJuBWNoZxXKeXoMpRJKoGYRf+pc3
+HB0nN1plEMF6OOb1MmHFd/2mx5+6nzT/wG4R4g1G2eeWBD36XfsiYxwR6czeiclw18F3oh6M2M0
bKJ5BSjsaDm4MJU1226cCJmjTChkxggp8OgiKqpr44JF4cAYieVby2nHVO35sNickJNXNFJjkUsG
q9A5CVvfeeCuD++RJkkHd2m4Vwnv+qTZCLK2+cAJMF4iOuGjX71InJvsfu6AutP5G89EyA2Glqfq
ejQF4i9H7LrqZM6edr9VnUpWFIjwPn0C8Dw5Hp8Rv26sGYVYQvg4pn9bKhTxYILKjBJ2BtVi7Zn3
yPIFMCSONTbIV3KlvKKR8C4e2RmJ8v6SgC+a1Qsvi+HUTluNI1KQcHXUEWwwEsm6Gdl7MsHxTia5
WAeXXVbqcSyRi3Q3hGAKfbM3RJ4AuBzs0EIaI5DOFrJ8ojbNerCDLM0QvBcadTrH4PM03PyDP4U3
XdfcquBEncxFgyAQwPp5CeeFl8FZyQMDPtYfc2CUbbVFGQKqdEwBYzhuV7cUNx2TfsHe5oZrmdti
Jq8BF5uwwYeWahHfhbiIw0f4IG6v9It2Zb75i6fplhGXDgYK8Iw6mcKnvuO8kmHFr/Zzm6IrMi+f
lVND3ORKc0mPKPukFOm3rjItYUIE+FtjUisVTT7r1DnSwHFKTEA2zkOFhLuJ/b/7q3JXL9MRwHYI
915EyDWiQzbud7WMwq8vBRqcQR4jtSXlJAnYs9ck/zgGlwDHpsmYpA2C18x11YEZdxDNKTDn1CAm
SGVbRyUcoadD6WG4/tA+Ejmutc1RilT7MDQdrNnxAQfdmaokSxsAI1EABXsbLBAaP0ZY5YGM3fuM
RDFdXdbG6wT3dnAVy5MsV0f9Ipeu+jYU2eLzK8Qsu1vKy54ws6JL/woAMwObhFOWM0vbbeQxWnQS
dc9PCrie2m3BkOBgdmN1cQBrfUcYoKPYGody3xUKSXXo2C5Hjn8SHlkHJMrK265dU0pmG1Mkn4YV
uk0PbGBa+LlnwWeMkZNk0f2SimWKx9wecnuxipYRpkUMGkJTYRRuhIHYGyQlz5ataHBkdBozaZgV
ORI056QCp6gEL6D6Eu9POvUuav9f2jb+LdasVjDxm8Ap3Fm1ypJg5eckSOd2Tayv3yZTJZPZakLS
NW+Wafb8JtQHubpXKp3miQNTQ6aTzx/lHZNmEXs4IyZ6oLCt34/GWR3RWmkncY5r2OH5UdcMiYcZ
26n4LdUpFkiPERyUPbTS5g/ykByVqyqImYUEi6JMRiBe54mPGGkompa0s2nWCH55N0U/IAYR4/5g
qfu+xqmz3vH45yV9jkUNtYVjIWNmiFaEbu/Gmn8wtwi7qExcYHKTZwMEEdH+qzUM9rbSb/MYEyxL
o0CHXkpG8Vxc62To9maVhWyVOzeb3q/xkd90c18vcwp24Ze9PdozSeJBl7HIhGh5Hcdrdt6UKgVV
akPTF+9+WcRoUrAIdoDBkmtjTOO4DDU437CUKh6LmU0+ME2IbfV1VrQWxt64dGLlsWdqtFWgFTJl
2Eb29acq5nW9MMM5dwNP/WWjdbKqgrc/NW8hZ1bIZKbJ1nvkIYNqVDEgGnwXrqIEah4z/SYwIwHf
W+XiEZZz9H50LoE9pckr43ggkCnlRV6TxlzWYbmbAXJXMc56XjtKBrW4dpGFs80La7uHjmPhHcRv
Xl6z5drz/596DCn2hlNcL7+biQcJw3gj2nqYRhanFrJF5hgUq8ZwVafN+fpHlLOGiJLtvGGR0YBh
k21yDRXoeztnBItX8qWePDfiLt/SCtu6jwuQ9VOEfYM9VHD/KfqRibNYnsgsB3SmsM1uswqgItKi
ZKoAINblD3xurfdX17M+fA9a4BBD6ME5vc3igSf6NV3abZinIgYdDm42xsd4G/0SWOwlrwMnO3cI
PRYUqf2qPLPbbz8GrrehQEsyahUnQVcjtBPAkHItysNoKGsb2Qx42gJM5DDvYuaTutIhuUaMS/IJ
rnmPknZ3m/Q4xhByJbs35E0lQW/59IuzIDsIQAkqspEEzgVm8YniKjfNeHl2Wl1+gqhdtA1sBFA/
2ZE1AcaXSL6lz1+hOc+Q1Z9vSXOBcLc9V7NDXdmsqAy/T4J1/nTDpOoX/j7ELVfdfl/QV2ke24MB
m0wbN/zQ+7KbHIaN8JtHnMpy/JJO7RqNOk1EO7K9HHrofdzn83OY5Bx+W6vstCPTvhU9b/s3eQcc
vcow5XY1QUZicmMv12YBdJa2ll5mWeNnqPTM/m7Rep4hTzAXITATLJc7YxXQ1TXvcrIVQcL7OBS+
dFfNL7ELfCwc13SLVJsAvq93z1jmt2FCSZwZgKiHDa5mbTfryVIqJIATlH7woFATD44P/+yef3nJ
K77RxgKH848yCY9tZBfZVnSqVmK4Lyg8D6VHBdV7wjrnySYo6yb37E+4STG/IdkzPe5WQ6ac5FgR
MFtAKgVzLpxMWY18xW8fR2Mo669fxHbKV6W/IeIV4Y1GhUr6L4V8JnOdwONnhWC+b/3ujgYM7Uni
DAuVFquGAayKnG1MNl8SUTftooj4Mh68UabH8F0APsn6jf1AeXT5zJujv/jilZCZStgOed9qYuka
Bi/Pjr679jqhQ3WC8micpOI+4efQO/8hLWnlkIDPdpqdtFryGk/7AdU0Q2rgjdWLVfQ7y+BlGdPS
Av9IyyNnU8v5gcG/S8zyoeFoARQmdI+VlZdWcZSMJqKWKqrgf5MAAXepMHAGBEHJMLU1avCOr6t1
1+R4RR2rvLcoK1nF+sXw5w0KPp5yDkPtjcPTtvjevNODuLmIbWZepQYV5cxLncjIpBDLvUTXbOpw
8Aq+nV3LYuJELW4LIJBnrhO7mmW1jxxbwnHgol7d+ei90iXSOk2yRO42ZRi8ZX5+nXh1AMkP3zwJ
x6WvlgY+/wTJG4S3maeb9YW/wjbbhgDZRYeL4raKFqFVJq+2t/6PkjC8GWtxYkAYAjUf/bouGQsH
RrsZX0Ud8RWU8rOKUvo4lUGH/XIWy+q+s0V7u25s/M6Hts49a8ekRJk7GFEAMTFG+lBEeSLAs6kp
kYSsKAy0JdtfDpPyciKQzPFWVTu3qGRzAlm9iIHhJmcR1Cu6SfuXseUGUEqwcW4C5tcyUxHhJuAN
eaGN4nCGPnjwvzhijxAWvW+iWYKfsSxSizuAk8YKzQcTHB43RaoJL6PTSZbrslr1mzDFqUSpEmBt
MNn1rUclOFOQCnuQWJB9vMj4eX0uwcSm2QR/UhznVPZIizu/vLLJtEZufglc+AMX/R4GyyYqdLWn
O2kQkboCXrH6vhOXdY5hHIW/cLDz3q47gYZJRkXX9iKgZOM4Ii/1LIFzBrOtOQRxMQjmQo1mv3pm
XeLPPXnEIqK1wxZJZRSL/1P4jjHk/cb8ylwFXlwGXgwP1O2usncz63A/bZ/3xS5MYy+ZhA3SENlE
s1UM+6eaRjYcatxCZblbGpZHH9WAAjzp0arLhLXqqY+d8bXAxE9jysjkhNNXh+NmasrVbAl4eEMX
s3uTdYsZ5Ig3mhxGArQJjQek/30YCnr99dZH+R4uLQeIHvGdyUiHT9WG5lp6EaTDJylVDjQqZqV9
H0Gx+YMOeHjAGpetBbXzDAKvffahfqkiwX9VW1wi7bUfhzJ/FU19Xmf+rBTrPZCI3SASberj0Zrr
3FFYuiB/rG/nSLYHNtYD2EEi0aV037KK6bsM+oyuNP2R/mUzpZro5cynhfpjzDYAs1VUyQaF6TVv
ulWXd4pVzzDpZxpKanCx0TvjHwW04DVvImensZ3rZuwpblKYL533YJpK4nEmaMk1xKH7qLzvgCXI
RiPMJhfcW3f/APCl0POXi2SBtYBoOE6oUtTLSa2jc6xEIMy0JRMr4yuHvr6MfMoRd5pzmzEvBTJx
hSoPE1eMWaZGNz0magG493DuIQHrcX/Y1QWgfJs8M3ZQvZ6hyHgU8YqucRsF1h0/mqq3ouIyclny
sLbF2Vz1mc9LGYvQy2OSdB5ZxgGsALoRAfSZUsqrn+kYxu4uFzKubm1dyhn8U464IfXTm0AugXWk
Mj9YNZNUGIziaRhWsowuccNrdOB06Ghkm5uXF8/tJIeVblcJgSEGqx1HVTLcmbPFbKBuHxji7/cf
V2RIZXcpgdzCzNoOj4QDIH24ZFl6A/FAGhciuA1x4FSTWiaMp4yLZ54dONz8Z0mPN7Ewcc0U2gpf
GTdAEzrI0f866pJeGUhzC6DFFFLliBbaYLrFk8+xp8Q5fQ67YX+zbUK0uoV7NCN8Lsuet8FLkI7Y
iVy4qvpNznHmpUL0B1TBRZ+mgNhO5o+TqkQKq+dATscfNKB20WS5/arEB5Lwb0pWUqEbVKp09lID
Zqo6sjYkBe4XGN7Dj0SCVMqap3QObWHejpzIDbJogWkPnUfxUab9W19aHLMbLG5SjQBUjO5/lZ2R
4Y27Dx/1V2SehOj0l9XqPEz0xQRueOCiQEKRVvA91D3jv0xcQUj2+4+G16iJ4e7sjYX3xys9yekx
yrkBLaE3nY+nsAkVvn5q6mhEOTwtCWmiavHFVRWaGt0iNCKEbIUL6bllp0rjBysqf8CzPtbVEPYA
NOiin3gi2ZdStE7Gqvo9fkYoEwyuAtpX6vHgBKV9Oa5Mvmj7TB3IkXGs50qX6HIosUd62GBYYoKF
g6cpXSK2st3B6RYWh65XWQDhd2XAMt7KydEJg9LxVLWROYMBzCUnJwrarLagZ8EwCPVV77P8h30L
28lW446E3VaDfEqNAt5EtnTOWzeEuxPNo1AInXkO3k1AH/kugEVTuhay09lSlN5Cadtb6NiCCip4
ySf6kYkle9zNNJFdEtehoWpu5mdgGCsFIsT7D0g19/Mt7S2FDpASRQD2U8vB7YdHxD6A1NBcqIOy
Pqu0LF/25MovZDrklOZTO8pZa4cKN+HEo7onQh7r9CtGNNpXdFUYir1RdkqSBrJfrAiuq6XWT374
qTYNuQkncTjctbf0L4+r8Mb6YVYM2Pa+FNsveyj4ptcq6G2niJFZQ5WOW7Fz72hkCFtix3RLhywu
HVr8pIiQIHLwkgo3DoLey9I52FSJPcmVU/JbBiOB65jszon831ztHm+M264gfGsU68pRI5tu/pUF
h5sazFrth/DXhTvjkBgdZbs1vT1kDBgLU66jkMNXppo/Z7KpRiKI7+H58fn+RuGbqmdwjVcm2Zs4
BGTYcGRCMBcKq7sTMZXShb68G36H4tJMFXn6Y+21V6AQ6Y1Si8gBqlWKJ++fKcRo8d3+9p3zrMUa
f2GHlIB6OVuHYoCsASEKwhi8Gio7EBaLbYN8ugWJ3x/w7/1CEq9tJBAl4hLRmM7B8mnL0GSfTLZY
uQuPx4la6L+ke1cnHoAeT1jg6sOVVU6MHkGYjbkMqN5kEzbJ7Dx406I1YQstfNWL8I5RiOAx0FfH
qHOyhYblE8snF5A0awuPZ8NM4Bb9nWqlyICAft6Cv6KSUPfseoBg3/HQWAChK93rLQAd1hDsdT4k
VM518YUu/xfsILfwTGurfYCAvQi7Zhx6XMjMGdLG12H53CFxu96f0ffLdOeRnl5WH+nyLfEVmRI9
mz8pyCav4gWFA2JFrU4uWfZD/cDkppIVnjz0s+41EvkNFwlTv9bTx1Jy4bIkqArDF5WzLOsAQg3f
Xqs9qU14PfJaQJp5CDdUuBCHtaYSLfNESyPxpJsVkYanqXLQe426eOojU6HhK6vfODsQ7X7OjvOq
BR8G/i3M/xTO6RNvnYad0LqCIGA/0z/EMDRVMVj710ENqgzlABpmmqYOpyoG+gs20zp5lmTTJYM5
DhB0X5ctM9y4zUrsdINX0D4i6WaUB6cBetDEOfN3j5XO3VMb9JZxRzAC0fT0C07MbK1wZWNvkOEl
rAhYSt+bj6EcDYqcn61+f+l88uzu0MdivlXQtsajBPRPynhshAWNMKTw9uYwu0ZZM1ZZg2vJXJlP
RGt4pdnAo6zqHLr6XdGcdR3B8Wvazr+tkgGB8qF+5iSzREFMbv+rnQMniOOe219Tkan6RMTFg9+I
CpxDcxFpYdSWn8mMMrMLkUrmXJ94aEKCbBYErg7BBA1TdK/A5HM+KL2fjMCDJmrdY08WAUTu/odV
R7IF7cY+aiZWjaVwuQkR2VhQdVW/xML9D+T2gBG7k3NMGblXkAPl7B9z33SBzY9LdmXdtSHSDfNu
z89k3ajZlaw+hcsfP/vYs1+6MwpCV306rvxMpKVVCHqBwNwjYLYdfpEdT33aHbtpB1WwW8KvB8qs
QJ9XClt2EqUPp/Ez55GqpefQyGbj20bOg9+SDqGuJlZNJHPdPtSCSfRYrD1PFH+Dqdd0jd295AmD
RMsQdK2PPYIPNwitIhP85O9WitkgHnO0LqptUdkTRToDHIkL6WqJbUhbj5JjkMNiN24e5vGNmukA
2h/5R2znIMrkYewheEQV0EE4qrIlGnfSho6M4pLOf5xdMJhCgFC1n2JjW8MgXolDd8B00oN1pPQO
gTmiloyndqev0s/bMmHIxbzf5s4gc6L14yzPNR7z/MQWIvBAJFujlBrSv7oczAGpZLQUPriJb0fw
t6W1e3X/IhsZu+gJDaEeeFRuA69CgWHH9JsEHJhpasv74ZsQjvRfZ8MqB9XjyKoiu1r4DevTSF84
uy4KkVV+xzBCgWbQp5noCY3WFiAJEXh0VG7mL6KWqWacSE5nfMI8t/wzWZdziGO0YwdF+9818xUM
JTQfmEy9j0EuPc1XWVYwNs7NyW3rup/r6Qv/rDysa2FDLAJxZ+9A/TgzDgqKR0IR2uyVXza+DBef
FTnw9vFjePzrBliBhnf5bjV67TkZ5BXXUk7DSNrt74bSAbdY6buTBccLY66KuOw2u5BZ5Ggd2EEQ
yMsJrzQFr0Iq/r97FeUf4yOoxjxA/rsPDZV4lNcGts38TpG5KYc4hWKL2y4F6IUCTyFvXqE2s7Wj
Cv62LrSayfUuCqRI6ViQb6NJi1DHWLHXA9ZvaV67DNbo8fDauHedUvegOAWcpbMOTcVUjAPgcQYM
WVefuovqty7AxH+6FW5cKOI0Swu02Z2iND2i5p+6yL9fFPJPNcpQp7ltC6fxnRqvJGicVMGLZ0EV
uaavNFBYEfFklUcJxoHfLPJ2vBGK3CqHSDb0EmBNZSdOVPi0wCUGVQMh6foN6g0QIwLtEYGq2Rak
CNXSwH/6YgMiKGwyazzt4b3xDvV6aHrYk8ZJ85EhUUdl/IzdWy7ZLoc5Hr/ati0U5jEHiYvpshz7
fqNYtM61FKrbjuOSlPi8FUBn+ld2gDaD8mGuCaOcEC3/nfP8B5cZOhmb+BiSErkeCbMuBUaaoQqg
G+Uc9MrznjIkSJR5tnhufs4NFTMiR8228+nO+YR5iIhCMr/PYJnlDmDg8z0kvzVmLProShWi/uny
bfiEkTcDt6KHtFYU5rkgBKOAHzwdqagwvrjXy4mFtnlMJ8uPyi8vaN3oM4lpVskbExVhbnWrQhKW
Lw9dCuTX18qZgcFZNW5r7JLmSORhKTQXX8wvlaJCsu2NirzcBI4Serq4EP8qOw8OuT6Mcz6+FTGK
ogRFrqpkLMgJHsoobVGOJEwN0/zvBe3VmIKjFBDelHvk5rM3l78/XSif+YqSk3hmabAGYpaSi2LJ
TanNdNT8ZyNgwZgr9G4Mv9qHUX/3HJDuPhlzJgdbhbvp9rGRCFFANoWeIlwmCjvn3ts6wrwSUJ56
kLlAGZWlhGbwNlB+W1CBVRemvJEbqYRSleH66DssoPoyh2SltfIcE1GQsNS6lSHt501KySaiU/eO
14O2Uz2AbBBuLC6rxQVc6yQV9OuB6aymRobpDSuYOQIQJjUTKx/SzloLpDzxpzwoQ3Z6gg9PcHsZ
nRxWlG2XwEEaLD6q3GvsB3JD2eHa/qQaAEh/C/UbCfkCHiAcHOYTvkMf4LBddtgqsPYf0dwjEc9N
w4XUHuWgY55KxSzlytWts/70TgfD2Wfm2x0uZjvQZjCu26C/afrsuf9YMzcLmAHtAb03cgyKJZZE
KwG5RjF08b1OBedNabJtI5xRCb6SIQ4tXEkva9Lpj7JtzfCphTPrbwIAJ/M1eog0xvUiMGCiyW1R
2N5pPcXXzbcsQkq5XpbKoHtPv7FfiQ96+6+2ih9Boh+7Sbwgd83ZnlluWztJqMKlYOpLduP2aONT
TYS9PZmfTLWaI7GW4S8yuk1vzJ8uW+ikAvNa0ZZ1kcPgehqF5UVKFrx9nITzy8Hs0e5Uld1ODb7F
UumvlCfkfa31Fjo6rmfaHoqBbaZDR+rfjQHgNEnWlABqIsU1VkGHYg7HD22Ri6v03oKwSFntU2WN
X3nDlh+U3QGuduWKQN1dwe6muiW/xKUovJG8dQnHQgAu0OTnVrDKefm3CnPgkywNktGZfhOn3qYy
DnzbNPHGVF/8dn26m/iMUzY33dxq3vJCoGReIbewFrBbN1aqE3EpPulg9U8Hozr8gnfq3wE+HvOq
Xj6AM4IlBKFVhwXU05QBw0eE4ATsDB3Jk4U+uBsEYhWVjhgU5BgxVX88JsykGoWAy6CrKRHMPVYk
ofETjOjHceA4G/KUwSsiqn07hTNDrAmReAaf+GBSFOcT5eMB/3jiobVUkD4DDpSRt8xsqymqdl5p
Iz/yxbiMUeeqkwHKUUwF5E2bigNK0S77zhF2Zr396f8MASfXx7jXmdIS5FAOnNsX6tcN4jYFKhkv
qjytnUer8E2Ym0wCq6yzUDctWyDB6ERouJs4Y5lKHuwdLEw5MbmC/eEgDJuizapDPmpe58ZCUXKt
elWIzcI0EYvueRYx9bkw1ON1bbvtDc4K6q9c6IcgRttqNzg6VsAOaaGAe3EOtQKCetWM3y3M8+20
rBtr3wNXCz5uiC3gSu5gRFTZVbMST8x4lcv4PzzRY18Q8qspT+mn0xekSVX4rebUnuulEEgsS7jY
ublLW4Tgt0+oFe0En8dEk3nrC5O1F9YxrZc1zUgKNIbUiqdk85qYIsOoF/dQabxhZNLcIOaNhknw
9HjGzrIE4M5ruBGuVsPXN4Gi5MlkNnJ+ljkWKYwk93SfdVSHE0wd+P6HThKQ6tUdD8Y7qughnsql
YeMHs6B8xEIVVtkN+sA0Epbb1Drl29q+SYuC1PEqfO6tbjJzYfPGjVLAMOKsFCGnlKuevocpCSdT
5o/1weLixOz71BzE4uD69sPR/yRV0h8yj8xZ1QLvWm+ZsJghJbYVr3btg7IqSr8wEoDqkyNcgMqh
xaK7DpIdU5NmnWjukFTCoNq5pmGSpYEgE1JnwSFLX7OsjNqiHF4RWgF2HGsOPKyFLnWV8+6dwbIn
xYFpni85xiFxBJnOwi6qV1u9zGXHbMk22XeCvdjJcvqIbhtZ4auIHcCEHGo1jMQRUR5PhCPfXFY4
dEnjirRrGxo2US4iWaJIjGF9ZARiTTbdblarMqf2Pbb64N56r/69TRM4bOqgcItYZElYKhqZ4OO0
bJIQQbFr2EYc/QpE+RKpLoShzaW+EnZrSo1WFWpSC9HcZ02gOgkqMWEoq43t9b8iE1NjHcfh+LdQ
VZJEK2LbIlzO1THOSA3l6MxxVuJnL4jXAVKybcSOcyZWGrXKKkMRSMwe4tHHpG3J3kzYpwt2n1w2
fG907zeNz1dnOfTzKm0tKKv4V+5QHyxUmCBksNJ1jG9H7vSj13Cx3+K455hI6atBNM3v/LhKzZF2
DEsJ/Q0ERNJOJCZRSSZ+/slXpGC52K9HJAjjaWIKFizo1r3Xx10VaeCjj6zZi1k1N66EAuj6j8ql
19MfukFpYQ8JRM6gX2H0ceaR+EUVcCQFmmx5ThonIH/qyRwVcU6Awkc1/Gg6RU2qI6943tKsuc9y
xPEHx7JWTamRGsR+Wo35neoZ1b0b4TVB11r7Imh4Rti7mtNCtGzEqLmK9HItIcaWepdwPqdNifQ2
4w8wY0V2kCosFgckjl0zUtRHlKd9NJ/1IDVCJ8LNAUKBPZqhodmXqjDzrs4gNrVqQS1gf+ePukhp
omO1BL2HLDuqyxYNJ15bMWOMwXriwppGUKqZskIIFuRAV2TxoF5htGpNcQtwvZInH6dtlAJUdxyF
pt7GXe6sfSBQ1eLfuyGtSVJ5q9dE3JEu3Re3jiXDXG9CGHkPThDazbNvDhx8CNHshxtQkgog8Xfj
SsQaUUMPNwHwjAZH2vHiqQwxEWmF2gf3k4B/3G6l89L7/yY4VR9yn4VfiaYhulWfXiZwgfJl6HvH
443XXsXB8loew2rpAs18HCDXOPYjHskT0VIPM4JC1tx6TYSyui4hfU+rHBPflaa+FRa+KlQz5y6N
TSwUXuHz59sZM4E+dleUwrJFgikm5ftV6KTX8ZC3kXil3+/8NBHSeoUwF3792Lp7Qtrmge7+X1xf
qYlkTl1PEIRzkYEZ3onqMpvoRrWA9rqhMJNbYeL8knT2XMn0Y6JKsznjNYc32CuwSqowJc9pz+im
pkJDOSwsMzmqX43LIU9mVCiBAYOiQMmn6e2cL/GSewmU3p7keU54BKSgYnSBt28lZpo9lZNoDb9I
i7/v27KHzfZwEnMryHVksTCDOk01T45NZJF04BViPIzydoLGhsyhrKV1FGj7tNysZnB5t4N7/aRx
F+xqgz7Jt6aMgmA5mGM5GS9NtKJyO66h4WN1CcTJXJ4F/1lf5s05wbJe+do7R39u+rR0iTjoEi21
DCmRHEnzaDC5TWPWGbygoZphMxC1I87UFWjevPX/NHc4C4SGkAHWZZQAu7/J0Ex8Jup2x8kpMmhR
fD55PfyFyZD2C8iCw6QUntlvkAFmu0S2IKZjANL2ok8xP5ajo6ZsHva85tN/NSuwyA10PV/1ym+L
GPcgOuPKpbwr6GP1Kqrd2zuheMd5CVNgtEisptHAZVrznal4Zgos6i/9MwM8mslbDasYM1Lk3RBr
PMb6oAWfqMYbu/IVAWn8ODra68+TJyhiSYc7+bnYLEiSsnWaz7gljZI5zTWHZq7GzVwZJ9up9+hO
8FaWWlJd3TGsfdLvrwpdWX4FP/1e9LN8qEr7dvnIgmwjhptrNwFE985OA7UJJECaa3NiUY4w38eO
SWWC0FO7GCgBvrbHDfK7qL86wf41WU6NZ4EE0nZI3fD+apF8he8oSZsM811pWjW+9OxGGpPNQ3Cj
MO5xWp8djdX21msTBnrE9P2lDOI1yDmOYFEvInYqNxSps99sHrj0RcREx4q0KohBWkpYtFJcUneV
wIU0qKGy6veh+BRScmMvkfzvGu1Yi8lgpHp4ShWD6CncUvIVBeKC1qliaV2D0kTP7v+vjWKzfMYT
sR1/3s2vA5qH1I39isGs4WpenO3RNMLylKm+d02C5INte6iwj0qzZBAoSm9hq7a804H0zKASt522
MwFCY0eNoDuipMcaDT3E651LYl11LPdTrBUtvv8MITIXtiKDzUTLMESQV9HJEADSCBVJjGXHMr/k
tw4p0eSVEG8JvAjWUNSKVT951faFqwMWIBB3oIqL6s1FqG7vYQsUBsdgtfekHbubsTh6Vf5cBjpM
TDsGH/dlLwOjTBgbeyMzTOJckSUY5LQs80RB81U55MKJHzyijG5i9jNp55/pKhz3c0nRSDM96KeT
rgikvzw0vqwsIZ8/ER46GDL+PethehmaAMB9oZS0HXS1Gvi5PqcVF7nvIBCIJ5QoxlrgtHYDxEw3
K4oJPhD1stjXYaDpk1FcyyQSJ83k8r/c82FaHcHgv1H0FKsarIujiNylaqVvjXx/a+YS10XM5zAS
6eiGaUzGSenNoPik4ohPgjLB7XHUsWvKE1M8LQiXvPrWLZ0E7Kp+qKvvt90mh/eqmuBGCGU0xL/l
1DCpl1FWPttB7iPK9CfkeXT5w88PisBkLRz7jQfm5o4eYfAagODsWCEp6IX7LvlE3nSzqH2/dDVn
OCAuGbYx9UvffVW003b4W/dfoeS21y4KAU74Bl3xF9Z0GPYlWaiHYMyiWerLQoB6KlNv3jFKQ688
hqasDAbX7BIO6LwJSwEPU9/8vDXWNbkafENQv8ckn6kDR2sYij01pI4ucuy3NT8y8ANprRntiGfb
Pc/IXgZWcB3RYNTfP3hqh899IA8yINDqS3c0DF3PlSWlYyNyE/txOs3GLPRt+I4eURW83s4RLDgg
h1JvSlLpofanvoSYRkCiZh0ThL9ck4DCmVV/uPYs6nmvRDsffb5HhQlfHhR1OQ68wWIMpsEcdA0q
ee3UNTcnbWVP616L78EzEddL/uOstxUD00d5tDCqE63eTvc92jPdC7fVfNM2jNWixS8expnPx/Nn
6jTYioz9PEOdM3j5lXzSexzzov+KAkyV2MHFIpoz3ateWZFCnIt6JViHs9+NEHCZEuAvUW8IWsKK
nfm+iwoWHumuNnFKsgLq/MtKQD3uvoDUJGc4Gf8e6+6MIS2gpih34iM8wbWh8DjZjHORpdibv78W
GT8dp+vjocNWqX/a3KgGXi6Vs1OR/Nr0n3grtSxPOauAkWSS2QZ02GPAO8BN5ntoMs6k8AQUutX7
R+xBox7+yUealFFgyn0pAmp8Xih8GPS7itw7VyOEdyRBjtg2VvrcsgoYD6JLswaV3O95w9oW6sqc
Xn/fqM5ZPd8XbgtCUmzwN6d3Wxb3pVjpNFIHj0cMcJwnwO3t4sH+4c6IDwv7e3qJIXuyWE/e8S8r
T89it4SKXCynuY2E7S0tGLHVgRg5hShBHeIt8i7e+MxhRHAsObM0pAzTq9uE/5rQ0XIBCv4Hr25v
5W4USHjI6PvXz/Q1Rw1efuxGNoFrZlvXymrGpRE2JZ5uehmAu21CMNY//QAOvkoG6kWM3qUqWFBb
NosBepVOeJjmD2JnGraq0Dyz0tNwCXjWOrePZqoDLDX9HV7Ptx0QVLuZKwXOSOydUHij98CElNdM
KqYa7niWvX+aF/sB2/nVcWE27NEOqFQ2h+Ra/EXstXZFeSfVlopzULhyocbn0L71sAWb8iIJprot
lj9c+qyMaYxjElQa3BIm1Mfv09KkCoOCgsfFx5hYbP0ng3VaoC1R2JaNJEmpYzuCNsT0c1HK4Llw
mdAkaE+/mzoQkvjV7tKuTNeBI/BAXDYJ/F9bQuOZgZzIOthZZensdDgQjuUh9a1XHMpTXXhwTwU9
EyYcxT7Z5SVB4+5nuzUFpYdP/csJ8cCxxxtP6hLvZbqGWTo6ivWKRnViVegxm2c9TwO8OhXaIkbO
nM7M/HvYSike/vEWRdQStuawUYmlfJIThPBbFudfrvnhXN9TQc9s9dlta44EVU3GXhXa1+Zp92Q5
RFPLfYSnXFMvQScn6ClWq35jtQd9B8RvEGJKYwY0U6Y/IxOlttTmvD27gAs7rJq5fF9KBFJtnxki
eKLC8c6YKHWjnwveiD9PrpdPmHrYt3Rknm4xhwLj8aE/Q2q1QG5YRtws6jbLS9B/9tiC60LWeptI
w2LOGKD9xjpqT2IT33B5qnnkh3uRWhCemMSTG6Ai4QYKSMq+YUFbr8js1o20ATHczD0wsJblFJ7r
CZ3ovOKBL2WH3LJ05LBFt5883QPFB1YR6tsniiDUIN0YoDSpVvRILscKapIbJSbdAohSBaZ9MTBA
pAJ05UYlvH3Hkz7faACqKwCT1Y0YtS7jWqe1NO3DyiFZIAe7ALl0HsrYktHgiM2fuxyi66e5AK2g
yffRXKlkLocCyaIeiecjYnqD/oUU642jl4F6lWGS2V7n5N0TewKqPCr041GwioWYtXVeU0mE8vzK
kfNjAZEABnAxM+mCcn3CUBms7kDFKWEXAwVoAZH0CrjxnAiSr5KYb/0gP+NleStoRoNEUdtvaa7N
cwpTSqb5b4poULAeB2frNvXTHkOp3SVaYMg3IsdH71mElMTKOXVJgfnYiNYQLgy4v4PTxyoLOGXz
wVBNf27LtgU5mGhD4bynvmK1IfTgZ+OONzSioGQX05kcXyuWSqQSMB6D9bhSYyzLRQfOt0vPXnNB
G6wbgtwFayIzxxy5FjWUpCewZYFe8iaFoTbJaqQSytuh36VJ6EDWHlk9Il97krjewiZNnKDqQu2C
1bRykEJ/o3LR3HIEpA7WRPrODXAxu8PzBKUxLNfMDe/XDhVY71wKK8SLay0BpE4xQYP1ceVTunJ5
JtCutpQmZXzGEAEmsKCmG1Pnm0VueUH6Gue4fJKTfZ6sWPPYpaYTwvqbNnB/yfD+pQjCnxfsc+N3
IVbMs2Ksq4b72WHfj4yEMM1XpArS9vFW8ZLYdpEK0E8pAmOw96I6iw4zmrhqwcI7dEPKrsPdc8My
lXfPXip4mTWJiSWHUnCSGbwNxFAc3b0gw0kmoaqTdFwI/+8enZRqI0NSAaNL6xzSRY4zeTCNrLYT
ssyb/zDT5viCC6WMhoDaDmrfE/1s5ow8IXJNLToARO38myN6hViD5xDKuFWPEXmo1khV47xch3GP
boIt6s48LybHqV0mBjhXUzDin/7Y8k4wzqJMbmtQM5SF9/RkkpePxpmD0lWVFElq/iY1SfNEf1+L
6xitH/qDYeT2H1Y3xL0Oaan3DtNpLZ0VR5sZtg/j1jqD7pBXxrPyedfHfQJ+WxNB8zyzBlaGVof4
nnxueYMw7IrqWsh2zeiRIkizJSuYBssmLfvlB40z5WwOD5wWAgGmatTzrF369Yz1nX9OlNFkzxVT
m1cm3Kw5vg1Hn9QRb4yVuzVnx6XMSQac61ZXs4Zu9La6x4pMr1gnlAHNbzIjs6sOmR21cHE5vHTR
l0zIRRq8PUGjQAkmrO/IhuKZ8D6OQsVk/B8ef4IG/LtJBppZ4xtJd9lgboiVz/HHfBGnTg44uj0g
hz/mRhaHdLW6CrZRz4xRWrUCMJzcJ0I2rmsQnAk+5Z8TvEYXZaFAkw/AycpHyHOzDqfcBezbR26H
4Qe6orzCCt3NowsBgkw4B+SBBOwE+iRxwPIyCOWumQqiUI7YdzHpcXPADKFcqTMzI98NRZToNNz5
JoEGXwSfYBewlvE0/BbMia4oUnCRg7LHNvEawPQi/mmq+siM2G7qY1bjIiMpKa5i1q8P/Sigrot0
7g6VKfWAZUtvaU19jkLTuliEnM+mVKR6g1kTmQ0arPuF9qwLyqspbilkVQMlSsXlVkiDJiRY7F4Q
dXkWMdIap8f8obF+1Tyr45DCRu15IpOMCgpWf4IGiZChLU5c7mWXv3fLiyiczS7h2HV2/YqGhhOM
OVh1a8+/4SfRTZedpcu85ZckbWBtw39bLWOCEnz3F4ERATugCMffd8VFLWYD+BXJ1Yi/KZvhrKzk
hk73QAVXeevAWgxGX8qga1CM8h/aVZzlbN7f8RXoQlbcF7H66M4Pcs2fVtk1wimzXyLwtenp3SNd
MiRS5ff/pSBr+3B2t3BERzSaQVGy2HuOkbl+NEwJ0D0jMuS9GET34f6SGo3Rf6ObHS/3OIxCxt+1
ZV7hu4BO69m0RfBNFiIxUroR7zC3/C5YQPCapkR4jX6fdkdxjMFN79qqQLoksOW9kbD6XYlDOR+9
w9CotqSCfGlN+DJi2d64VSlyD1jxV0i860aemigwD47h7kzgdL4enFQ7PDXQIYzHqtdpPzmHl144
tU34u0kglubGrYD0CNBFQealutS52A4ZhNElnTClqMa2VZGMQQf5PnptMs9q8MbyQb6Ys2mcdyR0
plA66XAAE5EpDNHPVT+ZPtN/FOfZiWkjvW2ralEOaLrSFuQDzbs/oZsM29/T6Kbr0YUOynakOxbP
HP5qZ2PsEv7cqxE2QPc0pnPWuwwGMeiwkgkBUDFYB3ZUDEEeqkeWru64gb9OnlN8fkvR3cowh9vs
WaYLNjkVLVTgJ8aQVyABRfREa7F7s0JQMO3pXaMz3KdAn2r6FgywwNdMap4wd2jilv2ec7gFntTA
ofL6LA13nddMza9EXspx+HF4J9jWipzsJIRvj+iBdneOQyXSsXLKOafK8nk/QtlXLg1rl7rHnJKU
vCyyl+k0d2a2lKY5xUgH5JVgCODnTn270PgynkR2RZ4BDobWuhCHuz/r2yLD1hxZrl+OEX7aB/hC
E5xmkCq7FEqZc775WFaE4I7t68d0FkfnUJB49X5f4KPqFz7kSrELvIuhcrcA4Wf1RxuhmRwpb7UX
53XVmxmxxlLaoHFaP10ejSoYIEggnbZNNuzwHM7U97ElEBoXI4ugHMZmicYL+9sFECPtN3dHIf3J
FZccVg9l7LMI6/XBeGGi4+WUHLTMQKst0Mn2qzBEAKB+FgXCk0zG4ZsDndE/HPHPnDRRGAlM2+TY
/if0QU1t22OxCt9IwJojs8LHQwZuP77Hw3gM0jEQM3goK8iQDPAlga6tnzl582SyJYxkAX7aEC3g
p89F1UC0ZlT+1ZW4vX5242FSE7MUiudC6BohKBnG4AdXtaz1p0Yhr4dYDVcAYRpj3mAWGfflITkX
2t8eoct9h19QSXxVzxrQ9WKbXe73taQtAgumtHxYdTe4dwmyj/eJnsPENqMAmXsSw4Zz6EJp1T41
NdNDHzP6Yl5q7+8WFxXNH4GkHAbVQkYX0F4zdF/kqTE6O9yyFR6m5JVDFEXm6mCOaX+JQv8UXRaU
v1JmOKLpxfz8MkN+PvdKU2Qz7DyXY32PGrSwlO7gGd82OKj9KFadzkEq7PTj4DRwuvDN6r7VjW3L
25iKEEDtlGLr/rJhhT+dayqrpIrI1XRQXwe5b0MSAsoNTbHIWbCoT4iSGxysrEBheysDAww0dRsi
wHjQz1js9tMaYLf/1iMB0l/63G83G14Kis2vPguh4sx6wGweIFfsnWmaPNbn7RjzT75RwIgt7m3r
oAEiJpozT+lhJtaf04Gn7cB+QGwJz8YglAlhsFzTpSIP7d7hi8/7yDMErLuGdetaULa0L2n9TTxT
Fa/OPPsPvlpmIBivTf4o7Use1E8F7LxXoIctFt9UB2VKAtRWOsbaJoQp6xtFVxXlQnAk/oC3wtmj
E2+ZAY5A6s/Pl71YKQGu2A+yIAmKlsmp4pgc3bmWeVTxfYOA8lF0f8maBXYlEZ1b6VWeNXlAVc6+
NDIF/w474MLBoEgAGUKRTFJklvYF9L479ttdEY1MTwYHq7oW8MaRX3bD4L77cBNm7wXDjxQZ3t0x
N+/AP9Z3ZfROd6w9GT2b7ekOSyijF6jrx4l8mTiBIMnNQZnRorul4xEIe2psGyHvE1Sb5hvhYwPj
oPL186XycKNzl9jXvlBlL6nN5lNvgHGwTmqtNkmQLD1WQzx5ow/cb1qTTI5NUDWzF5sJoDL2pWlp
WYFuevICT4TiIw2S5yQzw0PHdkIOgf/fx5GSIPPDcc8F9naC5xEwDXMHt87H2Nx2XNGfodaFevlj
D0P2XUBa+QxwWolZN+v0OjntboAzs5jCuySe0NwSwu9zZi5623P1yB41ynAtg7suuskYmJ3fhqTg
15Xvp3XSuGO/AgXWwF17vg9i3izvBmZes0rF4I/ndFERcH0Zchl8V/HA3eC1maS3VQCWkvI7AUAe
y5ok9Wkyrghq2B5bC3lBJyuL3LkoN7CdSd7tOU1VUqu3EldWe1Vj9HQ1WQMKzamQpj6ILq9HinTd
rPtukl8AcOY2o7/pn2GdUQu9CDclyGEu57ny5VrMVlEKXqa99pfZ9tWwd9kxaqbVE0XtWN8mvhRR
lkKbXN+pWtkqMNRjDXxPgbNt4iU3rGzG6GZ/WZRd6FjEOorHCdd2MGUADTw8R2ZXcy0yh4IgZ9Z0
P0BfCfEug3Ja1AZrLQGx01x3ASAi3ziNDLB4cFmxJFPmPQ/jug0Ulvx96Xm10JYv0ZdpqGRsoZuk
KTzQPsbRNJ0jYsYOzj+GpK5nauyhWSDxi/OQZ3kt+ZZAkDV3vKTuJz2g2G89yK237sbRW9COTTO5
IbArkYY4D2y8H5ZkhePqWOJ8hHSKxG8kQZHax1aU2m9Qu+AKL3lOHTc+QXM66z8Aoc9dOSoH1TWx
Dt17R6lPDqtOR4wdkKC7Q0291uuiQ+yY7FURZ05c1v/sRRxB+tEu2m7ZoGuf58gFeUEqrMZWoWWA
GyqiAZ/0Mz56CTdJdN5lljjGK8ggfIRGnuV2jpEpm5WmkYKKqpc1rObp3mBgwo8DfzvaYnI3K1zR
w3K2kxejGm0h69NEah09kgZr9LZlWfr7VGI6v66AWUMUO57r5fEu75YeAUdxbNEB9ZWeIAVfSBsn
EQZy59mZLz8lR/5JHxBP4qHh1pBqYF7/CaTGtroKCv5LX6MvtA6b4OsZE+/RRfb1ClKVJTosJsYa
AXfa/zXF3YadYePxhjWe+zoPTti0CZO0idIB2nm1yVg0kGok9MjjKQfl9KJEoqj6HVffB5I+wfyB
PC921olDIwCjuWoWElN61lrhrY1jC27NcFKn+1pFo979F+M1AlNfm5TSflQOND4b6f9Ei+/wk+zm
7le8MTwv0+Ie+qz8RFE7qwWuuonqD6FHDPh8uxQEOoov2h+UA2WYezCuArySTfjVBtXFLvXg2Sv4
3e7EN8hDYrQEyEnFVi6wYwmgFsXxY4/Wp7MGgrdY4EBmtm7pur+LOGz/A6c7+yv5IQusQGuhSIsk
E3s7jGhDyFI5dcWYrGmyEXZFlXSQQtZBj0uEDr5enTQGU3wQWxKl2bR9KIQYzQZ1Yx11kWL9+JP3
cmaNDAxaIxuxkuJhE/0sumJzaYrVcEagfPIKfP85ErpPPWSC4tjsuYnFSKqPjPoUl7hDQM21DLcb
sVe+yWS5UTlM9pD+PReEnRpcAHQcG6kc/KnymFqHqifBJ3A54F3Q+LY/5RxWp5BryB9BPunjGsV4
LF21Nq42++5FnEhabn4j8eSxXd67H8m/dnSw3ayyOgya8gtIuCtASguSa1RiDIXrlGfAPIHb+H1V
yJNd8pjmcN1d9RtG1jq5tR6Tn7aI0pKhMq3ex+MMSipR2YD0WgrxbmkTPZ0MOuC8p3Ll1Ywrqm+d
6ZERtF1JCOMs1RQrvuWgBiet85z197lzXwhS/Ynmspn3iJiI/mkEz4xkn3SLweGaHCUnr0RTbq45
fDSSVuq8uq2CPxfifB3MUaZHIKR4VmbHepCGo1TktnVwIyYF3Bw9vXckwkDwu1JbxBioUkpt987R
Fqsvuf7hg7W4JIV8vNFAr+fXKC3lF43L7Y+9eyq+64SbNINyh+hWomOdHFDhZdZ102CrPdzjpKTo
hAZdtdHXvoknrETaEmz9QiiSjGUx76oP7X3U68RMFNmrqHfHpU2i9fp9OIAz6QkUSaOqgshE5e9k
CWxnJyAndym45TEQ8Q+SChF0ePLeeX17Yx9RY+wfnL9nAt8oz9dP9zuER+D5OvMnZ2qTU/pY7dUw
FlZeDRVpLF85vYIr5y7L0DghfrK3GXtMrV1KOfKLS8EusjSwCKaRfQNx86dwxvcy748OV+iZkPBm
9ftWLceW6leIreDuUz0Ilgs0G2/rUpQd4NzScne1KnfBabuAKia6KDQUYOFqif8H6b8WuUFb+Isn
4TqIYx2qO2WEpfX3UNanfyQzHECl9Uqd9ZPYE1XvRdgMsKUBOwpxnQ0PhHLv6nMohcUwtP9dqi1N
yoA0VocB1Vca0ZeNwJUtJRpQSMoOUjNvBtnevztlX96YDgjLLqGxCKg+vkPfQWRiDcA2rrvX+8YI
Z8voKgdJ5ZJV3/Xi6eG/ghrqxfjZ8qY0eVWUbxS0/gVGDbDjEPWthCqAIVQ9CpC7VaNtFAoRwATv
xJ5cznHah8lEQcewdkFKM6drt41Wb3NgfKUejhiqSs0E8mk5mV9K7AsX6VmCOT2BNz4+GJJBPnMx
rJ/AeDgjjBwiJEMm4IlkKa1JXRip4vvrbFWFTd79TolhXXm2+lke265jjHzq3XWd7usNsOjUrFH7
ulm96bDZ88rT5NzrFJ1k5wn+K6+DQLKHH+290JkNSwvyDdSztz+8DL4X2PCG3gpEYAsnlpvJJSyB
pTSQWAT7MHKQWUsJmSuY04/uU8bq7Xa5BhN/cNLnlZud3bFF5IWXeuRRL8li7B2cmj3cCfPxAwKo
kAs/LN3jma96Wp5NcRcWS3JRDsHPVGnEBYnBaLeZPe8DR5zpnDdBOF44h/072xAvxfD5Hc5ofQBS
DF16N2ZDS+6RXsOPJk5C31YUHDc2bHzV1BqG3W2xuZZohBokQ/fyMvoGJAu2AKTi1Ta/vleupj1C
K6l0MrF+5qWwxHf56SQSY+I81FkpFPNHk59nHmibHJ7Nn1v+GmNoNS3dPUUd4ImAN3JgRgm1tdiM
6TufmRlfCjSYrrl8i5PSGlVcQLmAWKiWcck/cNRgemXpAg8HXUuhaHm62JBcYMC6YzjIOKXglJpT
jfhyngOyJTGroWeH0fyLyNJ5roA1LA85YnL5y+MMj5X4UQqQYbH6VAFQ4D0rejDUCQUNrMpzIxoy
o+HnLB+CVEt/EWJWpFuan86Y/69z//l+OZwuFvMI8brGdlpvvUMF+0+SNLUwjuuIVgt8yaa14pNa
JW/LCzWo5cNTYbJKuZgWG9VyNKvy9juAlFVDFsiZN7tXkAisStn/dAPrv2fovdsScc98Wo6prIrO
r/nteNGsAszLUar993wtWxQbiAs2tcuw11VR8dSIJ5kA7Sxs4U+vlOCSBPynrfdVAMwCVeJvSrEV
ZSAGoEINPdvKetmHdKnxRAEBqpKpY4YIIcAiGXdUtrK6zqbdsNQAUT99SBA9lEulBLJmQV13O0I5
+0vFnoVGGeZqpU1Cp80K05wRKSwS4TB4wetq+OvkvzXuRjDIQBJN9ZP4XkBCamenlXe8K084NPSu
eRdwTC6/H1CfEKwDSQnaAbwQL84mKttPvHIe2UFeC1yPFPy2CoPI23Ct2hBfRvZ767BmbtsvfA8N
hmIfIooMLlzXuvIxpgA1itHSX6t9ekm1Y9Nd1D8gm0iYOJOyA4csRCdzmUqyUqqkEF5ImKBSevaO
GqC2KECsPh13if/kgUXhj1P0xuhqLtyaUhhZB7DPyi0gxyb+fV6JpXe6/nv0FPthJgXPRTTIajTM
dn3zY2L8byVs8NdUfuUXyBylk5ohlkk7WHJScYQ/K0lrprUbvjsAPvriyXvnApVSgNmVtPzPn2MI
g7KBhEyeJ96PfJAZtFmTyOf+VmqgrcmXySDllQ45LTjyO11Jd/sWNu1+CFAeCY9IINbKGKWqStf7
mRYP8yVwgnUyXZmy4uTyVXSOIT1bqbk8DDH9Z+e9icxyhpxQq9keqmphx+MbMzA3R+6Cz6S60rfq
Yox5+0tBd5cDlvqFZYWYeH9Qjj9n8b0QDHv4EQjiVKhQWHmTeyEDBPSuoo8atM5/x0YyiHjwt9//
91AsqH4FSYmROpcLidE+RzhoPspAe/rx29EeXodmBIlX0ZbpPGlnGbewmUgPIlDuTdFFwqb9k2Ga
7YmJuER5blWhY+KaJQBQn8RTFHRlQFbjod0X3FsB+7SCxXlYES6qyFezCUmMwoSq7OG5AvZndEum
i5m8jOQIcx9WfIH6lrV53yOrd4aDnBcnDGywOge1fWHd9JrMkEM0tQz2TgEAhcZ7EridWfdVyVF+
jGBy0sONBd15JnX+971z7XUeda/4sjAzvbQ0mRRDae/HUaqz6Jtbbg2iKuqHPNcUsoHipfotUXK2
wXvmqnQfK89dejfMp//w5xCiau8G+LStxNxT61pjJlnjB/UfegS6z5WGFDTv0yq2LvIyCQ60uJ5a
XcASFUYBjjRvAxbOZZmTkBJWCu5Ht3gsxuhnNXRnlLS3YfSuxYMe/hTCG7O7xnUk2ZxQ0PU+IdPP
T0/9PVTat7yU3ygvDoSFgrmbLs8kf/7ELUW8NYulX+97uFdVDp+m+EK2G7J2KxflbTHONC4HiNmc
eaGBd5nZt/o4SEA1ZPISCmW93QrVB5KgPzzLRgCvPmegVA==

`pragma protect end_protected

endmodule


