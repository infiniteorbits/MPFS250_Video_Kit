/*****************************************************************************************************************************
--
--    File Name    : mipicsi2rxdecoderPF.v 

--    Description  : This is the top level module of MIPI CSI-2 interface.


-- Targeted device : MICROCHIP-SoC                     
-- Author          : India Solutions Team

-- SVN Revision Information:
-- SVN $Revision: TBD
-- SVN $Date: TBD
--
--
--
-- COPYRIGHT 2022 BY MICROCHIP 
-- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS 
-- FROM MICROCHIP CORP.  IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM 
-- MICROCHIP FOR USE OF THIS FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND 
-- NO BACK-UP OF THE FILE SHOULD BE MADE. 
-- 

--******************************************************************************************************************************/

module mipicsi2rxdecoderPF 
#(
    parameter g_DATAWIDTH         = 8,     // Width of input/output data 
    parameter g_LANE_WIDTH        = 1,     // No of MIPI Lanes -->  1 indicates : 1 LANE,2: 2 LANES,4: 4 LANES,8: 8 LANES
    parameter g_NUM_OF_PIXELS     = 1,     // Number of pixels to output -->	1 indicates : 1Pixel,4: 4Pixels
    parameter g_INPUT_DATA_INVERT = 0,     // Choose to invert the incoming input data -- 1: implies invert the incoming data,// 0: do not invert the incoming data
    parameter g_FIFO_SIZE         = 12,    // Fifo Address width in Byte2pixel conversion module
    parameter g_NO_OF_VC          = 1,     // Virtual channel 1 : 1VC , 2: 2VC , 3: 3VC , 4: 4VC Enable upto 4 VCs
    parameter g_FORMAT			      = 0	     // 0= NAtive, 1= AXI4 Stream
  )
  (
    // Input Ports                    
    input                                      CAM_CLOCK_I,                // Clock from sensor (Byte Clock)
    input                                      PARALLEL_CLOCK_I,           // Pixel Clock
    input                                      RESET_N_I,                  // System Reset
    input [7 : 0]                              L0_HS_DATA_I,               // HS Image Data from Lane 0
    input [7 : 0]                              L1_HS_DATA_I,               // HS Image Data from Lane 1
    input [7 : 0]                              L2_HS_DATA_I,               // HS Image Data from Lane 2
    input [7 : 0]                              L3_HS_DATA_I,               // HS Image Data from Lane 3
    input [7 : 0]                              L4_HS_DATA_I,               // HS Image Data from Lane 4
    input [7 : 0]                              L5_HS_DATA_I,               // HS Image Data from Lane 5
    input [7 : 0]                              L6_HS_DATA_I,               // HS Image Data from Lane 6
    input [7 : 0]                              L7_HS_DATA_I,		           // HS Image Data from Lane 7	
    input                                      L0_LP_DATA_N_I,             // LP signals from Lane 0
    input                                      L1_LP_DATA_N_I,             // LP signals from Lane 1
    input                                      L2_LP_DATA_N_I,             // LP signals from Lane 2
    input                                      L3_LP_DATA_N_I,             // LP signals from Lane 3
    input                                      L4_LP_DATA_N_I,             // LP signals from Lane 4	
    input                                      L5_LP_DATA_N_I,             // LP signals from Lane 5
    input                                      L6_LP_DATA_N_I,             // LP signals from Lane 6
    input                                      L7_LP_DATA_N_I,	           // LP signals from Lane 7    				   
    input                                      L0_LP_DATA_I,               // LP signals from Lane 0
    input                                      L1_LP_DATA_I,               // LP signals from Lane 1
    input                                      L2_LP_DATA_I,               // LP signals from Lane 2
    input                                      L3_LP_DATA_I,               // LP signals from Lane 3
    input                                      L4_LP_DATA_I,               // LP signals from Lane 4
    input                                      L5_LP_DATA_I,               // LP signals from Lane 5
    input                                      L6_LP_DATA_I,               // LP signals from Lane 6
    input                                      L7_LP_DATA_I,               // LP signals from Lane 7

    // Output Ports
    output                                     FRAME_VALID_O,
    output                                     FRAME_START_O,
    output                                     FRAME_END_O,

    output                                     LINE_VALID_O,
    output                                     LINE_START_O,
    output                                     LINE_END_O,
    output [g_NUM_OF_PIXELS*g_DATAWIDTH-1 : 0] DATA_O,                     // Output Data VC0
	  output [1:0]                               VIRTUAL_CHANNEL_O,          // Virtual Channel Number (2-bits)
	  output [7:0]                               DATA_TYPE_O,                // MIPI Data Type
	  output                                     ECC_ERROR_O,                // MIPI Packet Error Correction Code(ECC) status
	  output                                     CRC_ERROR_O,                // MIPI Packet Error Correction Code(ECC) status
    output [15 : 0]                            WORD_COUNT_O,               // Output Horizontal Resolution in bytes
    output                                     EBD_VALID_O,                // Embedded data Valid
	  
    // AXI Stream out
    output [g_NUM_OF_PIXELS*g_DATAWIDTH-1 : 0] TDATA_O,                    // AXI Interface ports
	  output [g_DATAWIDTH/8 - 1 : 0]             TSTRB_O,
	  output [g_DATAWIDTH/8 - 1 : 0]             TKEEP_O,
	  output 									                   TVALID_O,
    output									                   TLAST_O,
    output [3 : 0]							               TUSER_O 
  );

  
//-------------------------------------------------
// Nets
//-------------------------------------------------
   wire	[g_NUM_OF_PIXELS*g_DATAWIDTH-1 : 0]	axi_data;
   wire										                  sof_axi;
   wire										                  frame_valid_axi;
   wire										                  line_valid_axi;

//-------------------------------------------------
// MIPI RXD Native
//-------------------------------------------------
generate if (g_FORMAT == 0)
   mipicsi2rxdecoderPF_native #(
						 // Parameters
						 .g_DATAWIDTH			    ( g_DATAWIDTH         ),
						 .g_LANE_WIDTH			  ( g_LANE_WIDTH        ),
						 .g_NUM_OF_PIXELS		  ( g_NUM_OF_PIXELS     ),
						 .g_INPUT_DATA_INVERT	( g_INPUT_DATA_INVERT ),
						 .g_FIFO_SIZE			    ( g_FIFO_SIZE         ),
             .g_NO_OF_VC          ( g_NO_OF_VC          )
   ) mipicsi2rxdecoderPF_native
						 (
						 // Input Ports
              .CAM_CLOCK_I       ( CAM_CLOCK_I       ),
              .PARALLEL_CLOCK_I  ( PARALLEL_CLOCK_I  ),
						  .RESET_N_I     	   ( RESET_N_I         ),
              .L0_HS_DATA_I      ( L0_HS_DATA_I      ),
              .L1_HS_DATA_I      ( L1_HS_DATA_I      ),
              .L2_HS_DATA_I      ( L2_HS_DATA_I      ),
              .L3_HS_DATA_I      ( L3_HS_DATA_I      ),
              .L4_HS_DATA_I      ( L4_HS_DATA_I      ),
              .L5_HS_DATA_I      ( L5_HS_DATA_I      ),
              .L6_HS_DATA_I      ( L6_HS_DATA_I      ),
              .L7_HS_DATA_I      ( L7_HS_DATA_I      ),
              .L0_LP_DATA_N_I    ( L0_LP_DATA_N_I    ),
              .L1_LP_DATA_N_I    ( L1_LP_DATA_N_I    ),
              .L2_LP_DATA_N_I    ( L2_LP_DATA_N_I    ),
              .L3_LP_DATA_N_I    ( L3_LP_DATA_N_I    ),
              .L4_LP_DATA_N_I    ( L4_LP_DATA_N_I    ),
              .L5_LP_DATA_N_I    ( L5_LP_DATA_N_I    ),
              .L6_LP_DATA_N_I    ( L6_LP_DATA_N_I    ),
              .L7_LP_DATA_N_I    ( L7_LP_DATA_N_I    ),
              .L0_LP_DATA_I      ( L0_LP_DATA_I      ),
						  // Output Ports
              .EBD_VALID_O       ( EBD_VALID_O       ),
              .FRAME_VALID_O     ( FRAME_VALID_O     ),
              .FRAME_START_O     ( FRAME_START_O     ),
              .FRAME_END_O       ( FRAME_END_O       ),
              .LINE_VALID_O      ( LINE_VALID_O      ),
              .LINE_START_O      ( LINE_START_O      ),
              .LINE_END_O        ( LINE_END_O        ),
						  .DATA_O            ( DATA_O            ),
              .VIRTUAL_CHANNEL_O ( VIRTUAL_CHANNEL_O ),
              .DATA_TYPE_O       ( DATA_TYPE_O       ),
              .ECC_ERROR_O       ( ECC_ERROR_O       ),
              .CRC_ERROR_O       ( CRC_ERROR_O       ),
              .WORD_COUNT_O      ( WORD_COUNT_O      )
						  );
endgenerate   

//-------------------------------------------------
// MIPI RXD AXI Stream
//-------------------------------------------------
generate if (g_FORMAT == 1)
mipicsi2rxdecoderPF_native #(
						 // Parameters
						 .g_DATAWIDTH			    ( g_DATAWIDTH         ),
						 .g_LANE_WIDTH			  ( g_LANE_WIDTH        ),
						 .g_NUM_OF_PIXELS		  ( g_NUM_OF_PIXELS     ),
						 .g_INPUT_DATA_INVERT	( g_INPUT_DATA_INVERT ),
						 .g_FIFO_SIZE			    ( g_FIFO_SIZE         ),
             .g_NO_OF_VC          ( g_NO_OF_VC          )
						 ) mipicsi2rxdecoderPF_AXI
						 (
						 // Input Ports
              .CAM_CLOCK_I       ( CAM_CLOCK_I       ),
              .PARALLEL_CLOCK_I  ( PARALLEL_CLOCK_I  ),
						  .RESET_N_I     	   ( RESET_N_I         ),
              .L0_HS_DATA_I      ( L0_HS_DATA_I      ),
              .L1_HS_DATA_I      ( L1_HS_DATA_I      ),
              .L2_HS_DATA_I      ( L2_HS_DATA_I      ),
              .L3_HS_DATA_I      ( L3_HS_DATA_I      ),
              .L4_HS_DATA_I      ( L4_HS_DATA_I      ),
              .L5_HS_DATA_I      ( L5_HS_DATA_I      ),
              .L6_HS_DATA_I      ( L6_HS_DATA_I      ),
              .L7_HS_DATA_I      ( L7_HS_DATA_I      ),
              .L0_LP_DATA_N_I    ( L0_LP_DATA_N_I    ),
              .L1_LP_DATA_N_I    ( L1_LP_DATA_N_I    ),
              .L2_LP_DATA_N_I    ( L2_LP_DATA_N_I    ),
              .L3_LP_DATA_N_I    ( L3_LP_DATA_N_I    ),
              .L4_LP_DATA_N_I    ( L4_LP_DATA_N_I    ),
              .L5_LP_DATA_N_I    ( L5_LP_DATA_N_I    ),
              .L6_LP_DATA_N_I    ( L6_LP_DATA_N_I    ),
              .L7_LP_DATA_N_I    ( L7_LP_DATA_N_I    ),
              .L0_LP_DATA_I      ( L0_LP_DATA_I      ),
						  // Output Ports
              .EBD_VALID_O       ( EBD_VALID_O       ),
              .FRAME_VALID_O     ( frame_valid_axi   ),
              .FRAME_START_O     ( sof_axi           ),
              .FRAME_END_O       ( frame_end_o       ),
              .LINE_VALID_O      ( line_valid_axi    ),
              .LINE_START_O      ( line_start_o      ),
              .LINE_END_O        ( LINE_END_O        ),
						  .DATA_O            ( axi_data          ),
              .VIRTUAL_CHANNEL_O ( VIRTUAL_CHANNEL_O ),
              .DATA_TYPE_O       ( DATA_TYPE_O       ),
              .ECC_ERROR_O       ( ECC_ERROR_O       ),
              .CRC_ERROR_O       ( CRC_ERROR_O       ),
              .WORD_COUNT_O      ( WORD_COUNT_O      )
						  );
endgenerate

generate if (g_FORMAT == 1)					
	AXI4S_INITIATOR_MIPIRX #(
						// Parameters
						.g_DATAWIDTH		  ( g_DATAWIDTH     ),
						.g_NUM_OF_PIXELS	( g_NUM_OF_PIXELS )
						) AXI4S_INIT_MIPIRX_0
						(
						//Input Ports
						.CLOCK_I		    ( PARALLEL_CLOCK_I ),
						.RESET_n_I	    ( RESET_N_I        ),
						.DATA_I			    ( axi_data         ),
						.DATA_VALID_I	  ( line_valid_axi   ),
						.EOF_I			    ( sof_axi          ),
						.FRAME_VALID_I	( frame_valid_axi  ),
						//Output Ports
						.TDATA_O        ( TDATA_O          ),
						.TSTRB_O        ( TSTRB_O          ),
						.TKEEP_O        ( TKEEP_O          ), 
						.TVALID_O       ( TVALID_O         ),
            .TLAST_O        ( TLAST_O          ),
            .TUSER_O        ( TUSER_O          )
						);
endgenerate
endmodule/*****************************************************************************************************************************
--
--    File Name    : mipicsi2rxdecoderPF_native.v 

--    Description  : This is the top level native module of MIPI CSI-2 interface.


-- Targeted device : MICROCHIP-SoC                     
-- Author          : India Solutions Team

-- SVN Revision Information:
-- SVN $Revision: TBD
-- SVN $Date: TBD
--
--
--
-- COPYRIGHT 2022 BY MICROCHIP 
-- THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS 
-- FROM MICROCHIP CORP.  IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM 
-- MICROCHIP FOR USE OF THIS FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND 
-- NO BACK-UP OF THE FILE SHOULD BE MADE. 
-- 

--******************************************************************************************************************************/

module mipicsi2rxdecoderPF_native 
#(
    parameter g_DATAWIDTH         = 8,    // Width of input/output data 
    parameter g_LANE_WIDTH        = 1,    // No of MIPI Lanes -->  1 indicates : 1 LANE,2: 2 LANES,4: 4 LANES,8: 8 LANES
    parameter g_NUM_OF_PIXELS     = 1,    // Number of pixels to output -->	1 indicates : 1Pixel,4: 4Pixels
    parameter g_INPUT_DATA_INVERT = 0,    // Choose to invert the incoming input data -- 1: implies invert the incoming data,// 0: do not invert the incoming data
    parameter g_FIFO_SIZE         = 12,   // Fifo Address width in Byte2pixel conversion module
    parameter g_NO_OF_VC          = 1     // Virtual channel 1 : 1VC , 2: 2VC , 3: 3VC , 4: 4VC Enable upto 4 VCs
  )
  (
    // Input Ports                    
    input                                      CAM_CLOCK_I,                // Clock from sensor (Byte Clock)
    input                                      PARALLEL_CLOCK_I,           // Pixel Clock
    input                                      RESET_N_I,                  // System Reset
    input [7 : 0]                              L0_HS_DATA_I,               // HS Image Data from Lane 0
    input [7 : 0]                              L1_HS_DATA_I,               // HS Image Data from Lane 1
    input [7 : 0]                              L2_HS_DATA_I,               // HS Image Data from Lane 2
    input [7 : 0]                              L3_HS_DATA_I,               // HS Image Data from Lane 3
    input [7 : 0]                              L4_HS_DATA_I,               // HS Image Data from Lane 4
    input [7 : 0]                              L5_HS_DATA_I,               // HS Image Data from Lane 5
    input [7 : 0]                              L6_HS_DATA_I,               // HS Image Data from Lane 6
    input [7 : 0]                              L7_HS_DATA_I,		           // HS Image Data from Lane 7	
    input                                      L0_LP_DATA_N_I,             // LP signals from Lane 0
    input                                      L1_LP_DATA_N_I,             // LP signals from Lane 1
    input                                      L2_LP_DATA_N_I,             // LP signals from Lane 2
    input                                      L3_LP_DATA_N_I,             // LP signals from Lane 3
    input                                      L4_LP_DATA_N_I,             // LP signals from Lane 4	
    input                                      L5_LP_DATA_N_I,             // LP signals from Lane 5
    input                                      L6_LP_DATA_N_I,             // LP signals from Lane 6
    input                                      L7_LP_DATA_N_I,	           // LP signals from Lane 7    				   
    input                                      L0_LP_DATA_I,               // LP signals from Lane 0
    input                                      L1_LP_DATA_I,               // LP signals from Lane 1
    input                                      L2_LP_DATA_I,               // LP signals from Lane 2
    input                                      L3_LP_DATA_I,               // LP signals from Lane 3
    input                                      L4_LP_DATA_I,               // LP signals from Lane 4
    input                                      L5_LP_DATA_I,               // LP signals from Lane 5
    input                                      L6_LP_DATA_I,               // LP signals from Lane 6
    input                                      L7_LP_DATA_I,               // LP signals from Lane 7

    // Output Ports
    output                                     FRAME_VALID_O,
    output                                     FRAME_START_O,
    output                                     FRAME_END_O,

    output                                     LINE_VALID_O,
    output                                     LINE_START_O,
    output                                     LINE_END_O,
    output [g_NUM_OF_PIXELS*g_DATAWIDTH-1 : 0] DATA_O,                     // Output Data VC0
	  output [1:0]                               VIRTUAL_CHANNEL_O,          // Virtual Channel Number (2-bits)
	  output [7:0]                               DATA_TYPE_O,                // MIPI Data Type
	  output                                     ECC_ERROR_O,                // MIPI Packet Error Correction Code(ECC) status
	  output                                     CRC_ERROR_O,                // MIPI Packet Error Correction Code(ECC) status
    output [15 : 0]                            WORD_COUNT_O,               // Output Horizontal Resolution in bytes
    output                                     EBD_VALID_O                 // Embedded data Valid

  );
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="author-a", author_info="author-a-details"
`pragma protect encrypt_agent="encryptP1735.pl", encrypt_agent_info="Synplify encryption scripts"

`pragma protect key_keyowner="Synplicity", key_keyname="SYNP05_001", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_block
OHrTRdB42Z4n8CLuO+WZyUiuiRX6Jcgs5iMBHr4ySD3RQKgcek9GU3hHrU6h5pEmNP2cq7oZ0l3W
SpsQsVMaIIHsIln+yn7hcB91ltZIcSafu02c3RirOk5LhSLWVTy0RS/f+StKeP0TqhHyC4NhqYVg
+dEzOmhM+0hwQ4FR/rpkVs32jW6txmlPwwQLQkNiQENmfq8NZwNchUq//4X/Pv/2HF7hrUTk9BFO
PMI7dbNkJTJQruxv0dlPkslcPCeI3e578JVbZhzBFSOJ/zZ81Aprn90soA1wVjv8SQbowqRR1hY9
tf/hcCbdm0pl//bDj8XDgJh9qSElr2Qua03umg==

`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_block
psAwEFDfNw3w2rWTysfJzx6JLc4XUWnGMfEcLIyyCWykfnaSgnn1Yb6n3lUFFJzpzKPZASdmXNpX
wO6VT0Chs4W7uoU1NL+ChZatw30kIzSzIKJW6P55Jv/kxRwqM3L/Nw9APEI9ccA104CRxtwvaZUZ
f935hurXmo7hftULwtQ=

`pragma protect key_keyowner="Microsemi Corporation", key_keyname="MSC-IP-KEY-RSA", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=960)
`pragma protect key_block
HEDVucqGonGkbYG/ptn9IRiHFpBvWaKFd+dapwTQKY51abRNofIym/X2Onrn+VD1dr9NuuzGUMVD
2FSQQ2ORdqslcHM7ekN1E3pypfYmTzvPcvF5V/9blIYw+yz1irk7x5cYfn6nDAC4LRV3JBGZeUNu
A3b0PgkiiXyFJO5t6HWR791W7f1eRzgZ3J/IqP0n41reJchsRisKG/BBOvdQQ+8kxLJ2Z0949cRt
iZ8/jsLSHmV6buPL8Qhn11y3E7GcDho/zFSTVvLqKDN9gtSIKZPVhXadJypZYdku2wjzaGRnKXLf
BB5AksR/gLQ9D7XAvZaCe8wPek2gslt8Xf/y6b7RH7/gfftjkEo6Kr9AuTijTPIBTM71C9gdKU4R
iAx4rLZM8FN0kOjIEE8xLzpsxmG4Im1+qAGaBgp0akTIXhxs4ryA8in/mCNNN4iHSP/EEMU9qZIz
iMR808UwLD/V0cvvhXQbtjmsdVQZHy+94igunQ7zULoGLyrFxHtMfaoYD7EEy5LcCd0d08JxU1eh
/2NkhAiDO7pt4pGgcc91qIfUa+v9u+w2leJFBcG2McAdEn9/KVmRNrqxIhrWAv/m3B5hK0waRYZ7
rQAjff/qMQYUUYj+s4AO8FUjM7uV9NeLZna1wEu0WWTlWMA1H6JekwSst43HTew0goM7rBJ5rOGg
qpDS4U6i5j8YRfLTr18VQtTdK/1Y+p9YVWoUpaKDqTTuDMK1SYi9M9I/DBBjLmCxReyPYvVZzxc9
+zdkSB+IiyMhEptq0u0awR8O+x+775mvMsAIIe+QpjW24EKWCCp2qC0Ny4Mk99zXuHhoPV9jUrZv
KyU8vG9pls0CxdhhrggTTS6L3P+cDqzapQSgR45KZ9GJi2YAVktDszLgBK1iBZOKaemucGf9fBa/
DF/+LmylgUZ/caAJEeLDs/1L5yUeJviDG+E+u0eJHb9hOSfMbVAXSSQ4+lmmrBoi6dlrkvt9TZVV
OLqplCYtaVPkljhb1bS1q6DLAD7HhEMGmEjYJAX1HQd07bhwaJYiNfj1WG+ysmP6C1akEuSiphF6
edi+pm4WcQgD2jGJlp/BikuLR+fApkx8Ln0ash9izhpv56MUIXSkkIxBHio1EQZzEThuzP8sIDTw
j3dTec6PSheqgFC+oPc8cwqhN3wiOwn5xSOVQvyvAdPYauHKuh+T+MCchEHFrKZxWXlcgIL7pfXl
K9eTyC4EeSjL58MDnZXOv5IT6jXqsanbVnkH6pJdTkoScyLol4yxD4y3+UhvZpC5

`pragma protect data_keyowner="ip-vendor-a", data_keyname="fpga-ip", data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=317600)
`pragma protect data_block
m1bC52glJfilTjyVV/RNvJCioa7VYtP7ne9H0oTtvNqqRK04Bz4xqLlBys6ez6qy+3vnaWyLqFP8
E1YEPOG6S0ehdchcStKQlAVTcGE6fu+Sl7Q0GfrSQAVzgJ2dD2jAXIcRccVg9gOY5TOPOvbGdJ6O
Ad/T4uc9nGELsL/6yG+xi6ZvGZbkllhi18AzgwNR2pYN0e4MyIL7FzYCktKdaAlyHrJbEiSAN53I
Rb/Wx3o/CmD5OqRmq2bNXlTVYQMdBZxQYmq9VTPjV5wXtd1mSsUMJYyYgTvOHKwM4lkSN490Hh5X
Aa8OXI7zbwL6pEgBO4rkZARQmwOpLMcNzinIySdcwl81ghJYI7If0EkLvFr6UoP7SdJo+LMP9cVx
Wv8Yk3EMwRg+2L7+Ut8rGJVGdqX7grfHI0zTamEqs5RagA0qUEX6JPZBflcCxYsEdaANjLO+SU84
dMs2kajNZuVqMANSOlGoW+JNucrTbOrsYfgcYDnl/5n5FHewTfoSOlV/sSyMvUxmfGL4IlfEExWC
TYKvu32t/HIjUP4/dDWVv/dBHkpPCxpfWfDEOfluGGL6GQ0GX71AdAsR8G0ULQYcBrNFpJ9jDDqF
D8Wi8wuAn9tj870rZ7wTP0EgaXUNKF1KpEgsMwLScr3A/NF1YUVlkcZ+MAFsFTIoPw80kGcXYNIA
vusKCbf590ZQy/Z0Fxeb5LiIDggF/YCaVq0berzLj0nOGE7+G5z4tIhjcUL5DWWoy1e+SzbMso65
axg6DzxF3EFG43hZEG3K6zHLvcxtGWR14VKD6q/sGpMYc2+OQOkLtTxYelzWWbDMrNjbd62tVaJ9
o9TcxgsUQPTFdj1g43rqx2M/3Kifbpz/W/w8MjrOm3dzV/p2yJ3kQ52Hu4n5cP/EscsEqr/pVMYM
JtagWRNpLRNMobPMoHil9mLqYXE+aNam8Cp8yhnRba95mbyXDhvhbUzQx5devnJjBwnWoUqyyRKf
A0Lzyi1uffDlxbkyxu1EtzBoIhF/tQRib2gCSu08AZWShwUhXugv2c3tXtUO3zmohBnrWcDhYe0i
rs0Gzy2KFDc6HvmMfsqttVY7gaLV7CugJjnW4/QFsALRtSlcZAqCZdHRFw4ywNsTR0t6jHsUBUCC
LQhFdkV/cr83k5pgxNp9tI+qDyKmsueJ3wfMWczAPSV+oK984RCR8+iEjRKtbwmTdu676CxbwU+G
3tovTqUo9xZ1mxO10df0db+n81xOqoOkuEwdmgbPf/OXxv99ONuboT2ZpNrbl3ZN7whJGT6igWmH
FiVkaZJmKmUuOIszsDFohMdos843JbRAUbr8S4D2O2oCoUnJZVu8vr2wUI6COGaRMtj3lOumcYCx
c8ZoZNLMa5wn3KXxCtOM+U8ixJZ64bv9OfgCi50/R4JqP4lk1nvmBYU8EBYeRVprSOBM/FpaNzgk
p6DTTGCCYyZOF3T5TcxxlzjzdJVZr6KNDGMVUGJ07/ULVvuF6xk5Pwy19eZgXj4bb0aq23ERZF6P
7F0p8LavP9DGJkMqMvO4OX1K2EZY+mIFa/QzXtQApkAbsA3GZqGU6Y4nkPyrYfQKkdrPehNO58Gh
5P+9NS/SI0OMHs8luODRPON7/08Y8zD7g3BURIfcf8eFfWQDn/99ilLZk9GbDjoLh/DXe82d6pai
GikukWHJtMpGU7660VcOeLOQOqXtUB4YGBkHpk2tnUwCkqPQZ+UTRw93N1mdrdZ6+QdLyXSkh2/x
6dRnLoad+g8cjRRqVSysLeiuCxlndlRj1mTRoHdYcJL+K7e8hWnr/zrathK9tgiPRFJlFqOZF1sU
CzQhqf6/H+g5UOMwXhTD9jMZiV4SoQ3RPtcQV9hymMHidWYYveXI8wEje1DgIkOcRlHsS1YGtwzG
z9XrI2zUzuGH4jRmg5DZm0wUk6cpSWSqF6PVhmGIYNah4dJOpIETVEafesmHrgjOSpSNLzxAKKIU
auLDAIAq9xQsX0ZBNWuxD2IkaV/MLVlOe9/Ine1xlZOev10vSLydafraqK37GU8WxmxzQXymY5gt
jX+3oGSrHaUO0sqyvUP2duRdhLsUuYvhxyR7U5Xx/yWzUksu7uuhYJJS9YlFGPElSRJn+YfqT45i
auZaEJmfSRkHYhAJ6VR/A3NUaaCa9lJaPcDjtfwg4jBFz2PftDWZkqW876K/g1/FsbHL31EG/eXc
J6lW3cCQUVY5EqotVxkdL0+wAogoRNpEPOeigH66gYPpi3+3yBgaoDMlcBgur89b4dkDSdBDWPzH
qe9ElmkxsM+g3OXw/GVTZc9xyKvV8BEsExMev120J6u2MojfjBq3j60zSP6bLpUmruoI30M7oFL/
Fjju8683W0e24UABL6EK0JCXGHmMwNytdsii6GLE0yPNup2IMUuq7KgOcAlZ8NxyMhC+RwH2X8Id
fXCb0YzikOgsqcteJvXkrEH2/Q4RrQKsCVIE7Cp1iuRH2ngtwApmVR3bnje1xxbjfiXp9TQZQ4YB
E4zhYC8OaZaGMxDl2LIw+GNcZoSF3x+yAxGwr7ZKQbn337ub1P9cOYfsltLEed5BZNXmEj1/Qiej
6hBVpbjt/WTWf5/PkKEuktHqZieduc8tgIaRYY1mNLbNgD7rzT3e09qxJs1G/PFQIj9xI8wrqNzp
HDCURr1uzV9ybeTmosSpD7dCVA89FDVR4jWHRSCRzJIK5iVfYicmdY+EzjxMaTIpVwY+4t7MVpuk
MukEwqs7xzEhN0T5ImuNdcf5pQu8L2doLaJw4lloSv8BL384PeugaAP3QXeSvBZd2WqLk5I/5rAV
qeUmDfge/rEHnuO39P3UYqBtW09iECn8hz0xLThYC/AUrealGC6D/DqqQJY/yKNZeoAEM80cMDKY
HncUMP1PpICjxtfdmQhtM2cTz6AndIugdyiW57QPGSC7qrWl3iUDeJDi8qtUtDfH3zT1K1vr3hba
YOGj0cQgTAtj+YKanBIcFfeVOjslKE2Q7ochocKZxldgScSiCpCxyX1XpZ3uQsbmjE6oTLCqJTGJ
Ap32toMYmglu6GNjJmGge+t65ly03FMJFT8V6xQmgjDuO5czZ7M3zRChOqNZVoiWl2c3YuDoXGCb
YeIrJLwMfIrWpMVsxLdRmegXHoI3gJyGTuNiYj8cbel63uZoXN/ba/lHZHMghU7GqYV4qtMMhIQC
nwto4LCQKOIurRMXA27jgDUjPXeokru2byKedD78Z9x7TkUjZ3RZybntlx18U9lq0qNpCyEks4GA
RSEp+7/QvdLXKxDnDAQe9+RtoksFjH+PIhEigGxOC0yGp8pvRm/OsAhql6wIXqpwPrkrLcQXV/ll
xRlGAmw2oBl75TCAaZL5klHlWLoC6bKfxum2lzpjovHVRHef+KVjpXchBRSIFJDJo+HYqBIU1kBl
20oGXFHJWKYnJZ6FkA59xzOvB929PZexuqeWR135rbEpKOlovrp3rDyTUduoaH6SI77ihw9WZHYe
fJNOkE5LZAVWwmZCoUcwYGNJB42s82Ei6uE+PgwqD63WOqtJI22F5HP2bf9BWgSezqSYOSOtrX7K
bcpcxZOe8CXuyHU+7cuQZ72KmiAgYLXnjesYiXnYCRj1N1O0OIRero5Y4D5wINpx8SHvDSSZrkRt
BgSn/jikiXgiMPb5Rm3hUsqOoEwWRmBkfVPfbKszBXAKyM3rUpH1J+2WXbWNtnFYhiQFx2QxRtNo
lGNwAm1aUsuS/VCz2wsnUJDhExnOpM+9QBiggFqsvWw/hchApduj8yr1iI4aSW1cu+s2tVMGupgd
qmnIGDo4D8QMjvPKFyl9vQ9jiqS1/zBRjsCA80yB993+hCSxhIP5y5bxOieA0mDwz2NSY8g4Iw7V
Wj4WrJ/uwYHjoT18VkVYg7fI4fc6/J6Dj21UUcJfHr1aLh7NS2LPTw8505rIvG2YqFUs4JLDMAvD
MVsm6m/gQwGaMbI0fRPhfI1bh5CHbwhLBW3LNt8YeZV2tp3qD3MuSdSKwgzas9oPcB6bmxyAbiI8
tHpiExfOv8hHt28ZBreD9C6EpnqOn6VLQBZZJre+fX1RZo2NoysOGXk5TuWCEyp8os08L6yh4oYD
3yieJ9eRiK4fRwkKn4tB3V9fWZYqZUnT0lSoJqk/1F+tT7SqvC+X6AWWDFeScVTezCrH24D/Ou4o
PL//l95w6xnUM/S326ZYbvXvDsIllhc2TBmUqiVJpXw+vRtRx/d/UXTF2wZSheQ/wYAIpMVE/mmh
PftbN/ia+0A6XGUoK9WvtGzmEOz74NlfyjCMtapb89Dqr8+YxBdYoXVWvkph5aL9AU++0B7GsRfh
A+1Dfhx5fLCrFtv5jqHnOIDkGIL71OivU5PPJwn+DYzZAYQds9M3uCa/diqgKbuz8oY5RW6M4qVO
HAOspNs/4DypD474D9bKJQGl/I0jwGGo00+al1npmiOYok8bdMu3T0YCp5k7IG2dJjjM4qDXxnjC
c1w6YI3WVmFuwgjMorH5xcbZJBxHuwKeI/QmUQ45UmH3TT0nigzZmh7mkBHN/Vzmrs39g2S139DN
tGEhZTL7l7Gyxj4EirflOwqb5MR2arVHiHYjM8xg0NT1g2QB+FX0U2rpScF8NFN8VAmTErFE0FpU
v3Dwg9Qb2wDea976styoW9sPmSfRpWyqj/8yFaTM+LxUQ9+OVfLtLAV0+8chGSW09l5HsFrL9EeH
OUi00iqodH0t4N9ap2Kj8coe6vYdlQuViJst1vovWlH5R5GgChp8/a674eMKq0/3Vl8V3zLIws98
Ppo1nbLByU8lrgWqHanNliGcwMGGGN5T0BFABAXAWRGt6+/q9GPNvoW49u9hgaNy0veNH3Zn5KU/
C2FdClZqgAHV5FXBK0MD7GuWMIGZaevjZjEJK4fQL7XFq7VWgvyYAtvGiotmtPjsFr8IM5MTzxF0
HDIJzXPcF/OuYk1sVXT+zXK9Xcr/ia9CJ8CnF0glcoBKMCKE1hdWanhdUxi2qfOoiyWzUFPxw7qo
bGhtk1is9v0xsWt5Rsz1T/AiqLxUE1FuVRpqK1lClQumI4dvS1J0YJPUwUjj5BTkwIY5ndEIjKyo
W6o2kpSx7e/J4L7ottnak6KZs/QpsYbbVwNXFpKWnGuhlWzH9MnF7Jcey0eMkvJw4Kq7jlOEdfbU
ZCxU9c5z6riZWO3UfcTzlIKmsOtQ8F4S1Ecj3NcWhaLcH+7kR/5ggfuZvpfoYcGS0JVSuwh2sXgM
WzsKIfPkErdcZPWuZo3tC10as98l9LWUahffi9oDEbJhDJGkJ2TP6wumw4Ekdg38Rzj9h+x67YsM
MHJfo804jsi1t10DiD59I8jeXdiT0xCWas+rSzswdCrsxYxVdLmWmWgpCPscrVCnjroaF8Rx9TGi
dlE2rKmMnF3gs0jNqMHKM8q0g5xOWMF9ctfoi2npy1WAKfBabdXyPOMUFiyCNk691Cr5jTt1DJbm
kuZWrcQhXxyN4ZUL9AubNmXTDFTVPVbQz/HiO1X6VjH/l3Fz2ZJlkpuexwZyPK1DV3sAcYkTHNMK
yKHAwu82L2sRm2gmnPIZg0JsVSQf26uKzRCtLviohqNYLenkBG+7FAgnFUkSte/oc0Lxf8+5NG8d
Zv82BAQTlgIKCqMXxIq58bU7EuBX7XrsZ744XgEBRj7UxG4JFN/dVSmcuRAp84myVWo11Rjr9lbd
x2LdmWq1dCgs4cJvuDgoISmS4hjl1l4DG8uFbhke1DH3KO1vQ5W11g7kaqirBMLwvGuQEQoQEo7f
rxAbSGS+7W7IsTck0pI3OJVGs1NWPI3hZO7UV5l4JD8qhgLhBSVvk1RG+m2lS76MpWLxNBERUMNW
8M8M5gYfo8x3jA6f0PYWhKXw7oEVHS4K4uI5FGXsGfSGKSbcJx4XjAceIOboFB8niCFgfmxoQLTT
HgVv/MsdGr7Jdgf7d97vqBH9AvQUH58h0ukKQY5EU6QRgrhcglji6XdQGsl37q1jwlcaFDAqFNM2
CKJyBn8KHDqVk8B8+3J6/9cnE+HpSMMVBJYA1NYRaxFFQpSpdfWO3+YMLlTFI/hagGY9qAJc97ko
sgIRDG4sunU2u1sC+jD/pCG7t2MQBpep0xJrmCSx0MW/Cu7ZRW+hV/v3+nxzb0qzhZqrT4MlMqIQ
d+9kLH3pU47tFxd/cDpEJH174nhTUfLK4QyBu9YW3Ln9Wf7zuvA9xECdiPlpm8+YuHNzm88EFwrb
eIbL4mGnCsCt7y9WKDwut0thOacXNMZXVd1DEaVrZGL0P77Gx8owG53/RyAAM5xSHdIA/r33II4d
L90GfBIh//deKmDx/I1uHQtBipSgWUUbbYIZgbUxz5r44t7lRMTgm8MbIWZh8WKBC6UNg8jN2tJh
8P0KFU9nFECa0WrTs6jsxoueWhLIYyj5q8JmP4nBFTGu1/nx84TzmfR0sai3Npv1A7qFUhctckOs
cKUX13PL2XTvAr+WUemk4jvxe+9uWpazXdVxoL/YBtkVNGYWxxvVQh1n1GeCV1cxlEICqsd7t6py
wg7bbRLaqPIEnQr2ESvFvuLMkk/mIxILvaRQ3DsgMh/2PUKtHUpXSp40PTsz1HHC9aDUak65iQnL
diDqkHEp7ApC1QA7pK6fEWGDa2FDMS/EcON7eysN7l4qpd5f7clLDU1xZxFOoLecuemfLxS2ff9G
1uoWRjow+0ld0XDPVeZFv9dorb2TFqExO5r/MLmdI48e56SWvn8t3NwHIjPWKPCj8otFiDcL7MRQ
kQCZXpF9+ipWOYjoy828H/9upMioRpzsN9eTQkUoX80+TMhsvINdaHFVqBMjws45inQ6ZdKg5sUa
G+DAR31XIZGafoXaWRoc1WVXroXKVHs1fVh1hm8yJaKc47hf+5wRcapIVpKCk6wUSm0C+0mTPT0y
friyPUbhR+jp+3FSgahAtjMM337oVcyGsny1Hd2FCBittXvumoIRVDWysLy2Sv1HHuMD9bIIydh2
G7Co4jhwrFCuLc/dhMaZEiWEpQ/U29U/NqXWcGdj8LjuC8aTXOBkxAljD0bQAdNdNwEc4bQ1cC6D
ZOUohG/NvxHLolsFAG5eDLFMNMygHClp1EKHeN9KbKyxKeJDEQ/SmkL9rcolUOkfWke9v0IMocTh
01BbZEEzoS9pSYG3pT/vb/sIJKEHR/m8XhGvystOhs4QCWvF/VlNvPd14ZyW8juHK3679UrFbY/W
0uC6Naq1Wa7OQfEZvez9PU1B3xDVUURYwUZERw2Raw/6lMPIs8bCJNUdPrlSaV/wEMr8chYWKruP
qy7Y+3/i8KDpBbDRxKrRRr9wMIsnWsAKODbmI0Fth6eDw3cHqJXO2gdrfi41euqtZB9KCyG2vHKG
7wsqYO1liFeha2I26ZL3qKNfR3uxaihQlxchtO0nbGwjaGSdUv9vbleAxgeZnnCFw8/oYyHHKeZL
gSl5EQVoWVlwhKqqX06duRIT8U5SXDaj6j53nQno23GKHUjfmkuZtJiAy46eMv+iDEtlNfaNiPwD
BLQq6uqKxeVz5NTRVhNdbxIRAnZ3c0PXVGlccKJcLoLSDJS7gtJ64imO2O+iRlzqTRsI00iAqk3D
P3Q42BcKpOFb36QdzTbzbdWztfOFIHiyrClBWC244zdvqBYh2MqUuv97iWbTaf/HDtkJP6I5jinC
kvWYftBRRiFtt+qE/sfoAoX3yO7nOJb0oLyO90TNHmqnmr/Dlqu4bXdMJZMiuRmlfhtDgBPYD3Wv
MyUF/AbyOIeyUksAbXPwd5ZlF8cZ+BJxmr/6X9bN43UZ4B5UXFlYbYHCHG30dO88aZUtGFxi63GT
duKN/O9jp/DpuIgTFIRFDHBzBocCiSE88y0M430PGECK7ETtHo3FL5gEjxfL1q9hwW1Cvp7wlAiC
UQgOZWQkxpKdO0D5oeK5ptxlJtJ4B9Zw1EjuH1o9xRD23liqrsWf1+5+40v4Z7OHA8J0hid3vm+b
HvrHsqSZG7ELpNmx5ypJw3Pn7x2Ioq7mJADFw5TKCywz54gi7an6es0DKtOBJx/RBLtCUdHoaBwK
4Hx5CEnSdw8Q0XoWj+E0dTaC/5IHZTHt8yb/SqVEbb4ySb77zmlpYZyRQU/95S8o/F1dQ3Oa8KWd
OYAA4PEDfF3sK8ZdpzQE6ODn6nGkUi0fdnsoqhhqI5Sv6kEOeEpbISLvw11PytV4jXqz6S2oYaUc
0JSamih7QY1fGy2892b1apoWEz+MyaqBf8RUAJ++1Ba0tArdjvrWGXcrOch1dnoVHNRvGj0urYI4
9l8MDeN1pKy/X/rQQH+/+/u3KgGgZjL5KlchA7CP6coW4OXDiU/bDb/Va0i+ttaUe+Ru/CaSLTxs
zkX9Z6cujxmbJfGZt3DLrYIBgLUyUlRswGn+f+vAJiX/tpCUXjRhe12GvnWAOl3jQqf/zchbSuvL
F/6l0nW7YgCi8Gb4HBkXwmrogQF+TeLDJ99PFal4DeNhJl6dCVFtr/XyG0RSCjksDcmY1l1Rb2WI
cQ39ti5Gggz0sKaQBQpWJ3d8sePyrR3CUvZYLjVSjzahLBnNpx2vX6skrEKukZojdY0APb+D0qTw
P4R0tiNa3g6+eCg1vWL6tiO30k4SWbaxXfG5S1KxqoQdRaHSY+gwJuiBQfY3qw39cQkjFSQtiF0N
haxTgCpm0cjFDy/eBjcQuOzpttMKw2AlOLV3bksV71udjH5+SEkBVTjAdvSnTnMZMslkaCMyWLXB
T5nIWXEjSWvexrIYBz9tQ9s2KgD1uMnTcAO5wlF0AS3ZoiT5X6HJ5EJgA9sRITkrZh81qs6e99GE
vvYnZTMhPIeQXJ9QPA1wehLymuFsgqoHlKuifM/YBOcPv+bA29kJN0EnQ1BkyXorh2IV8F7ZdIK7
0lIM3TgWsR3jcmXhP3alrVTsT/PgTSiUpnDIbqeFJ2kPgihBmvTCb1GH8i2bXUPLibruxQxFhtdw
LshcevHsPpmiZerprW8hVXxNa/CxpFAkILjcaEY5dDQLH+bCyY/L/hwzur5dp5gIHovqcPYJuT9+
kULUxa12GZBE93LaLnzcCs4ZYtRP6MPQwlmjOeM64EUNuPyzrX+UAwPc1og4Yb7/aJ6E9Q/fbhn+
wc8Y5lH02UhtapLFfVyl4pm9jTJbkFiQ5pM6bRkb/D7fhA/tZiuOT6IL7rvBkyD5QjJOM/zt1taC
2PhKzJOvnNL0VQjLbXlNh8hYV2CEkZkxuqvvaqmsrTM6LlGJ2dgoi0TbafpK3mwjQhQys/Y/JWj/
Z+ZLV4h6uXpJv+a+kilKHJtDLnkPkBl00fM6wERht91/tolm5Weq6id1E3oHsnQSovp4G5O0g/Y7
P7ECUdYCJE+ukUUfAes79KbwyxGFzfl1Xo8GRJGWtZNtrieNFtL6K3mojJAfWirpC3lhOoI36lt+
5jiHVKayOBhFsipJJfab30Nc6DAyFsT/BHwTPCmVAzXRemK/MgSwNgZ7Bk2g28T93YNhc+w8YPd1
62Q861C5gn8A0uLkzgeAuz4C3I9KPiVO7edqmfZR0dfY/0j2d0jzWKCtz22hu9zuQs2jkZOYxoX1
3dPQfnwcBNC5LBeMadIIn6cAHinhiJtAKIayS6S7FuaCmF2HrCfT5OGbrOKj2gDodgZRuJ8jKxRE
/8NvIgw9lZNpnBQplfubUqUnpiTEd1MXkfhIiB/D/0ybH3FIsTDOW+6KU98Ba8djnb6o8GwzldwA
wQEnzpgXmTXquEjgQnzcs50rtpIyFodeW+iSRN1ELFZVwzN/Udu3KDWxJ5sWBdwHhE5U/gJlCc6z
Wlfx6g+wmpvQ/UPTe3KBGxz4Ss1qCEsiN8QPjXJU2dyaRokpqX0pGdVZQXFIPJXpfovG/4ZFYC7K
9fgpiliCbWRD3jFAjWpcYd10GrI6G4KO4ld02c14EHwNUXAThdJw5SvbRB8lL23rrd5cIOXOZh7Q
4KxYyDLTJC9/2eKpL+KtVYCkQwFDQLUFhy+fJMcf19aBNu3yBe/GOSCfjYXd+aP5AR2HABXN1dFe
EATSUM6DfSdgCCQCodRSG8nwXx3QFuk5D1hjtBLgyMcXnNmu+semQhBOMF5gueTWdTRHy1QlDxJs
loT1IcwYmESqI51w/nWhWYaHG2lTUIjiWBgFYNcN70Pk2ZVMu6xGE+AjqDXZiuoOATwSxBtkUQS0
lLmcWorQTHtmgsCutE9wvOpi85pXWEhYzsuG4tEXZYte17W177hhHZ3W3s6XnVVglFmqbodOPAI4
ztUFgECbcGVSKWumPKnyzYefHncl2qWOuYgU01mNvoMzoodvfFpZoNxCcwxgYAiXpeFyVqcXn8Vr
0loqW1R2d8cjwr6Vk6WbsJ0Rawy7AW5zuexjB5iqEfB/mpNvYTyPRIrEUhpQUDiWPo4pjwnn4+6B
afmoY9KDdez1SPQi/ptG/+MdWxWvKeY5ES5RZ/7DzHYFSiLlu50fdfa1zQGj+z+/nIR94y2SZeAV
i+cbB++Zx4HUxBd17bQDzhWwD7V/KWcE/lLBWtq6k6HdVDiSGX9hcIP7N9f5Wd8ZkA2dmp+0vAzZ
SUEenNBTN4s2Eo5VWplNFtTiVqzgQyzbnddWBM5Xl8Chx3sZLfd8NMc7XviY8n73Uq4MJucf3U8K
W95b/dwWurwy58geXRN4ZFvYCcqGzE4xgFm6KgLMB+NtitfwBvIU3tpoo9TtKNCYeNFypNrhmFgX
K1eherukzygoGzlCTN+70GsnU1MLf5e08qZtScP7USbMn36N/ymU5x6oSiOSCmzReCSqrxQgJCw+
hT5L9o2ZPtrZmihfmUwKvh3safju5LkkYGcscVXHPkW52fejyDz02OkZVOVYJTNhjDoh+/H3wT95
PRvLnOmu310YQNczwgH6i3HoKo0lNWj8HiLFsWec06t+tBQ4RwYBbJH1GGooWUBQLvgIdWDB0WHD
exPVKWgyC2x+bPlhVt+xtfU+zm3jayP1GD7QL6mRqujTcBvmP4BWlzwru2J7GXbikXznI26KGk26
pzHHWTIp7Tt7eatFS8UuQsbyD6XeueTqcVVL+U13ZiTi2i3j7/SbRCQ8atUCo89VlCYV+5TezRRx
fCIyhwNnJtz5m3pJEGwHtWzuv5oyrkM9i07X9WyNzHBB4WCqXdU8hP0ItgL4unfVBOKmJz/q3J2V
lfgMcILMh1N8ZvWgwV+7O4nm2FaDwKCNgvVNsZ9Y3TtPpZlZqdlkfIdeaTl10UTQ+LridU5ainyu
3bBVELr+CGww3uIKgBcKdUmhdF89KtLBC1YHPHmvADa2GBh5CLTD+C+vT988K8iJJcHVUY5w/83c
NV1M2qbOIjEw6wmpWdQZ3OkprH5vXTcPsLv4fh69R6p27Uu/LauikZY6Cr60UCL0EzenIesT7Gia
ArJBnFJJ/Xwg3gk9lZUDemvxkmYoROLm3c9E4LJIdAHPCFTKI9Oe0Yg91gJuogO3eOxY5ok740pZ
mKvX0IuAqzGAV63QWIPj3WQbuHUBv4Ax37VAqAmSkRMCO9Li2BN+0P9sNRrdM7gGhYdo3NWCF6D6
oeC662ucWq2yF9rUCa0EfT+PPjeJqfogHXl5Xly1k1SI81PQd82+2R8A2r5x5vy7afck/DNdWl8a
J1mQrxZVx0Hq+RRXkEDI3i2+F+gUC3mWKUpgH8BizjkJetf1gzL0fd0tzowyCgYaYmxNwqamVEXC
PURF7z9xONrbFGWH8R+vDq4AyU22lXVouePRa4IFuE8bNJB17nJz05500U6hlHA50CbGnEpViFq9
uEOQSQMNHQZbsOL1fN1FSLuUBSzPhAQlnIuUVt5dxIbV5QjB68ZycGVzxqw23HhwqVg+ZPC+HPkb
PV0FMB7kyrMe8TjKbUOAPOQHydcTNTqEv8StonTQDW/VpBTXmp8ayCk1xmtiqZlgfaR3Ojx5OP63
3Bkzx3ZZpdXnuAx3T3MQDDMGR7MeZmTXHwlhW2MX+eQAZZ1PiYT6f9RY8ayBmU36K+rG7QOxYE23
Q/2f41Nj931Bq4TAwjnLH+6C4/NnxfAW2wTD7XXVeYsSWer8imtKTgzrPxMQu99/OOfQk1pS13oG
k3vLzhlqtyVguVzP1FfJDyIwHnqJw5gQtWQispXZw1UWFv8mWZMDe2QhdV2yECx4RN/3WSYkfv0d
7/7ASiJyCqcY7qZgzG7UyuGGruLHhilgam2EgNgTnH8nTRH792+GYo4uC+b4/i9mZYUuHvT4slca
CRN4Z51W02mfVTHG+vR54PgLYBGqyik+UeHkZcfcaIxNi6gs6XHfkPmflkNex1l7ya3pHbShRsdm
zZ1xqXWJDgrhHG1M5k9JGWYDq8uY8KpMedHbPxH5rw/DL2sjpx6oiMD0TAx+68Wua5VeVQx6eGRC
siTw2GE0PNcaKmV9seLkCB8wG2eiBjFuzwYJcGii1DLFd3azhxHpnTEJ6dHtPeWKaIVZT+WvZvjH
JTa3D3SzeU+UC5XcqCQcCGGTHbyNysSRfG7LGD+ZBzxUNbtwED9LhMTPhSOxHCGhCjQDEkuO98yw
OtCUOQEZKQCBQkYrmjknEsCk2pq9CRPmi56Dm3p0VddzsxLtBZr5yijkKyOZloigA7ytg8E6u1CP
/ESVtMRvX82ORwG49afqVjSDfsleCQYzEmU235/NM+rBL0XhikSdb3TuWYPrvJVlEabGD5OacnZX
AbVQcMCsh7gyKKnDYOxw3CC5OHXSjVeB5jQcFtuaDHnfas7yKa7BHgh60j66w/Ib8FytiVewvEAR
ODFMmeEfmGV/c9gS2fhDAUbaECdngSk1thM24SWrj3D3dc9uknuSDrEu7CTE+qQH4vd/ES+t9aEd
DCak3H1OGvCmFB5crYZbb6Ntvvf/JhDFABQ/t84zGM+mff7eZK+sIF8AtsQM/DtWqeBxRRMImli3
mpucmxlVruS9IOwS4DtLNJ56ofuKAdh6njXi53CCZGYKEs6/Fg24NdQCEOmNzoq7JludVD55djHQ
0FkgfaAne1dHcxJ4sjxE8GbCQcPUft8baahEXWGG7f3fYGWRz5wGsDm2JmnBhm4PXqHdcM6rlfvx
Wp9FYSIKoII79yCXSjLP5Vq556XEEFeImlxOmO/rM0D69vn5FKGnprB9kD4p2TdbSp3zGOhNZ+o9
z9gC9CBn8naOacejTZyeO7Beyv526q7WKBISeFLZbJXIeiEzaynr4Fw/Lg1aLP+cyVCenej8BviT
ANAjGmvBN6Qle6/YVhK+J8zIIlxEb6TNi8GYbRrMNnRqNN7QvWl28j1/mqHV4KLHlX1MbGjUBnLl
TPS6ocr94Nv2qtzUlVLQCGHqr+4/4QglcPdZHKHeNgN03df5rWR5Y7zjxM5QY6ikjLj8GU3IAfXp
V57Rv3fa8nowu4gtA7vd3kNpFRZ8+j/jeRngNhKmj81oufeiiloes6Brufip2Rt0nRv8lwdoseiy
2i0ByoL78aLphFZU91IXTER0XdZWkd9hl1g5ATNn0+gJoiZ7tatKeE3lyILmCVzIv4uL1dhaT5x5
6brFhvrIHKCO6xYjFWUhei0oeO/zMgJV1v6w34L9Dk97tLchik2jihzVzoS5rQ2kSCjf7wg9CX64
JwHkS2RHlG+eF+oPdVamZeawa1/ljWQ6oMjWhJApd2D8fF+rqCN3yVEkK2evLCUWz0L77BRd1Prw
jv40+wcAhtg1hSYrUrRI5DtxPoh+rLv3K4xjmI3e9nTvB0YW3dws2Qwv40aqrEItjlpoJ9U8odZa
PsyNLZ/oL833ZkRJH3VV+YQtIC76fV5n0tMVGApKQYcYv9wHFp31/up1DFZwTstVwxHRCUAAahLO
rZpMl2jtLS7aQyy5sdhtd1EIYW0LvSXPll//eGdrD1S1OhJ1P1GkjlS37K3N4UXOZsc8wHvUfDvP
gKHCXZznAJJq4XShx3BS2kItF5kWczzZJroyGe9nMJdNrGxsWrVmzrLD1Y0dW2AckxgLLg9eVO9x
b690zkewf40pmNDM6jRo78HgrA/+BzY1csplaJpsPRJ4NWe3n4kw0JkYDjpbpq8iWhS0DvGwj/oT
NG5aymNUcjIyBpEUuwYe+abkXyLDo+YEF26ydje5MvkPZshqEmoeo//DoVUtJE/kpNaiotuK5Y09
BNN5eydP9AoBnU0fZcuUlXDP29YE3jd4tdM/zhpMVRTmkMEubS/dbe4mTQ1E1MlMnHRwmzplAB0/
I4fbLwVXYk87kcPidl6gRYWzlvE+eKDyrMfIg+AqwxhIq+5HRxAwBF4xOaog/LeypcehnbUNj+y4
GVV2IC93qmVWlhDeT4CTtc+8qOHRBeTY8Ll+wON2UHINEzLZD4qBenfda5cvuxNxmtRDwK1vD174
vo7lzSih1xJyrkQfJaip0iso5GNmXd28zXi+eVZV7SpIIPsDiKEpmRidIbG48gONVuHuN7bouAiY
a6EYd8H0chSBaezWE8LzQsDW7D2sr+edNTO2rB0osBtc6u5lMWsOYEcYseLbUrjPMsD29sooz71Y
Pykpbr1xwlf4QITApDP5iqqQi9Rl8pQv11/NcAdrMeOg7o+ewcdz8MlHJNZigCTBYQCLopSefH66
R1oWb9HVeUvtQKVhugFP3ROQwszWRwwnyPsExDhe/Ov/cT5jEJG6picdsagqtamd4czQkm9islmx
sJaGaZKySngNEpa9c9xXICrhJusaM337DoWE+E2hqnGzVPVT76IAiBKpF0y5LqAorFveuPv6VA3V
2CcQaIkcYCxWGFdsdscDLN2cst4pgb8zqqB1z+7sZS1dIDo0NzXTulqTLuKhO58ucOwLRCrp63rs
Kxod6PtlpczZJDYbn6y6slnxE4MLRZWoB3OeZPxFlH7g5Vj04mu55mwaORZj++pnRhprtYA7yoJz
fsFGBW6nlMfTfOWFPLCSvy0d1SFld3loGKKcLmvxQRpMIvkSXHR61xkD/oolMJYfCwPC/DpJPunA
gWc32GdWFq+jjfJd5CF9r+V+ryqlkrsjWunB0dZarvM/V2tiQQEVx3UWfREqewWGcWyD8xzHzfwq
jDdwHWXblCDaf71SKb9Oip3o1YsW+rFyJaF1r6S8jVqxAL4+Aacn/Tf9jkCodrGzONKn0cP15PX4
F7qfJ480Rbfdyfeclxim7Gimti+YC5opnielYTXVIqqVqYl1gIGr6/AGEG6FpUuEcYAiaxZZUMz4
fJAO+ELLUAHy5I8eVsp450xW5NTxFNPZb+tBBo4JicY+5n6IWWB/Vxz5S57B7H4bGEgeTbsUxN+u
LNKuRue775ak/hm4UkiN//Io2OSeizH1zLQnn0nj4TQHr9sNKUuwJYhKy595nakjfROO4VIdTtGF
Grg/6ECZKf4bHc+E53GknLynbnhmUCXtH75Q5HPjKBI0k79OaEH3ZYHP2oPb6KYdRGhAsjf7DWVn
U9JS2qGkETzqmIMTEjsJhKGg3NevA9nVyBHpKXnTF3/PdlCZurWiiaMtnO7YMIdl2sKIZa4C5F0l
lKbJvFfTVQTz0M19ZaP2NDuxMShC8k1X7ObfQIJA080i4PJ3h9u7ROxLB3TJu+bD8kxtTAA3NUKL
RYegaYw9JS687zcUkLXGkRD5BJWQlFTSICUIgiBLKeZmKQQx8zWt+0st0xubDMWGF1rgm4ulGJDb
HFs5uEpB4z7jIO3w47/2af2pyBNJAb/Bc6NZbBkBEzgu5bY2LDDtCGY1ydj6AFeX7Z0lexKyCOVk
d6TIU/x1xvGScK9pDq028o0Nvy0m4EPknt8tj2GbDnIEo9nDj78lermNRCx2PByPPQFRfzVQxffO
/HQVuJfnopU+vnddNYfsOfxi4nTbZYc0lcOfALMPO8g/Wzoe4EyEA+4AUYNq941VSJR5bj38aSEp
eQO3aIcxQgmdNYPb7c/UBwsEkJswwE8qKMGguOpmipnoUvbfEEooCeAvZv1o3mqCsuJ+Jp0XgDC+
7hXNiZWZnO9Or5sEkwCwfIkGfo8q7hhMgag0SfEvIoZj0GdIVt4UspHPGa9E8VZ8bkOEUhBEtRs3
qaaaR4bdiMfx2zx4WuXFe/UrOYJrGikE67132uF2TxfauwGrzRleOkqs2fMfKnMsgg5UZb2Yn4TA
aVWb8EsH807Aa5remClsh5slApSg7h7GQO/s6SaBPMUhH6nyEFe0gyJYp6KbR6sitd1+c9+HwuLk
DfaQJamIG8QEToKSrLmvFcWqYgvA5cw2uPsvzVmX0nBx0zWwN/7hhF77uvTR4WCCwBtvgUin1r+V
FgiQMuy9vev8u6EbcTO8UibtqH9OlR3ur40UUOIWUmV9Igt2mxmTdO+0j9lJPcl8T9d1dztsYAQu
B+t0KefKn6f7EYkXyd40Q5iS26myOFwafzTVQr+6a+SEOtc8urk0Tcw4XxKN5IY6MKIPEVgugE3C
bwme7Nhm1XkLI/OVmP7QajRW9so3jPOcAMhWDUOj8WeUn+2ZIQYH7zqJLgoPCfWZvJN8eURXA7th
inR99qLK4JXzmkbl8QOJAZsChnVQvUvBFjPlazwGeORSpXIW3LF+KRmRmdIBDBck0ZvL+6UsF3R2
+OKrj8o2XuVJNIeC/g9gQGz/M6sFVUpRznwJR3YnkAp8E+k8OHXXSsOGFirhpOSm+joBRTddG4HR
k6bqO+pBlf52ILrHLjO87YQ3C866rG0O5XzrCc1/GC/64EsSURDhaDpksPpP41HVOjhRklfpwppK
2tcmBfmoc93Etj/wK5K1Iw1RxcD8m8o9tNmJMdagqIAcei9cdwSTy+2Vn5tBQ3IO8zIKXHK7LuBc
0ic7YryYK7UDtv32FXRlD5CieqSGzIgf2NIYcFpHBoEHKtWZRMFhJNhekSq/F2VA2UngsTYq7N5Z
OgwJX5wOLSBKGpK0J7Vyylhndy15EJFaxNCAfYWCTnNHrqsBE80D6owZr1Q6zmJqOp+ZsSztnQgy
R4d8yLWt4c8PNhAoIP9MLfWQVXis48AVnjyknVdoD4FAY7G4bJTI0HO+I7z4XwGMZKHhhoiJh2al
/0PYvc17ReN7m7BEbvSDjiVd32LSXqRNBxCE0b1PIS69A/ivnQ6kNjakXEgM51gCTTyOYMTl4p4i
aXQ4on4NzDmIZrO8KGaSPGGwpYDEcMGzF11YyxQ6NkvgRGIo7At4VWkcTgzc4dL3+sHvCd8I/z0K
JPOusKKu23QI+FJ2XNkk+I9NMj3DsOwSoZrq9sqBGRwJN0fNC1bnib69reTWCFtkyfyYTyCrzq7x
epmWAENMhezRk9ebuSoc/PyRiTpQROVhpZh1nSNGkxUaH6AcFBPKZ3HRJXlXAMQnrZwjJIXi0H/4
TfqWEIHwWp3Td1f27sLCk7iFoZ0RyT2+tJYziPDJtLJ9MZHg3k/X+VSfWjlqKWIlAUa03CdGASYu
iB7N+Uytzr479nKxAs1vdW9rNNhkIqtKKyiv5EXFsit38fqBAoQTZ14YV9TZXAWG9R7FtAyi0ULZ
Svg2ePbAP1WwTH7OrGmUb/JpPFWmQeQu5g1dpdb9NxZ9mYfcTsPRcLNd1zAXjm0uZuvp+pLz89yn
CyRgUohiyp1K4UjZfLa2i7vL+oP+dpbG2IgrnE5TpmFXN9QxpKG6Rvhht8Y3T0I4yVaSmqr69xSE
7CfTwwpzZeEAHQWaRFfeUoSmTHxZVyamxQjL2iEjaszF/f3RAShU1GoeXVnuSL+5xfEDhi6X5wa2
zntn5kL8Uws6pi+4MnuIChg1i47dHhq0v9hnBz7Dpo/ZI1Jhroorm63bVMCe78cLWRWSNffbLeqL
oFsZHKqIseSoNHYglnTEtRXzGUA4DDcFW3Wuc2hEoVra93YVirheZPYDHHD1IH5kkF5WY9d1gBBw
ovxe5OSblU9gL2jXa/JBLKvA7Q2ucYUJq7Vte8ipQ4wj5zKPL1qpRSNQgdgLmYyqg4ZrBp5vFYbm
NEhMl2ANvrFtsLzzjPm35XHWM4DUQRhNrbPygXdpEPD4kSKk+deAK3JT7XAhHiQ8CJ9FZyVWfu9J
Nxgbt+7dMaB+lalqFdvU8D3c9MpwykMsbSWOEyzJWVuXFTakRHA4HEMAWJufDvpTU9G5+3GlL3Fv
THnw30hzxPgOD7WhIvQjCnocDnKoErjsHsjnUcN7IYISm6veULgP++/Ja3SUwrUf8lPET0BbiTXz
EnYlTg7dNmk46Vepa9w87Gvlv82+l+dfsbuf5ANtRO7TKlivauMpXbL5cb9cpW8AogM29b8CKYiW
tfsJ9E92vjX5HOrSjkwHmAhnf3I62kz/fs4gcRm8uhU4EDR5JX0ARKylPHVjn6QWc2PW6KPIzRm+
VQyRBEPZu/XZe1gke7Fquqfgay3ib6X8ojC76xApBO/8yjTWHM/kQLVBT+Sn6r1NlMb7y15uNd5v
farvY1weaBa2DD2Bc7L1dzfvEIppi+2hHISsUhhOMtdIHw3R1VS9KtnNm67OPOZXRO41TA2JkIyW
uomoiWQuA4vedvuphjfhVgOGWt8envnoZzMnFjBF5PR9o8X2FLBEH1b001kJpg0zpxw9FUYS4fqt
GS7hX1Md8++K9fkq/RCMlNq/hsiYy9yKYRz7MqNI2VVhKrFW6YNjaOW9YMep6em/A28tV9AWCnVQ
HEGF2IoM5LBMYjqTov2qcVZdMPfdYewy0AWG2ZT01evEEjfh6KAuDH+6eHFkMD3qAKYMXRrDYpre
jPbCTn+xb64t3BpLhYd/gDzW3THaTnlVf1UGqIep4LZANKA19Gve3kwxu9aj0TsHONoFch69D9aE
EN+3jLIVWSPFFnVYzsghzhzl9vSFekJcdW9jRCD+vuZXYTGka0djuBqjlG7NcRDxtcYOdHyGSBOe
6roQ3mDxNRrniLGWC9duECtd1ldTHfahIEeKlaFkSm4KsUxBIg2fpinIaQc8XI2i0sZARg0mqJG/
hKCL9Q+WN1QFIvjRlqMtjqI7oNJxln82y/Hl3Iu8Ccn4K12QtPEC5p2KQ4S4fQwZ2ybKKuo+htD9
DPNWdSeGWdTHKGuLrJQ4+eBLgwBPAPbCCDhY0JyXZSE7Z+iuiwgzLnnjjETWo7z64gYi1UZh+bT1
q9+7AnLIPJronxV/i5FAyA5Tku/P2pV3ivRueLOpvTepbGEFmEw3i4klT++Drah+G1disO+aQRVR
WNZxohaUhnu+3Dp7wNJAMBkhjd6B+z9kZL5ZkoE44eSJHhTosMa0nuiAoV7a8mux40mN/PxPnGoJ
ggcxn25/fphz0+l1RSgWtgFcTEXXH5AtfiPt7mw0U8NKgrPf8F1acnPaFB1qgoEkF1D6bcon8ZZ5
nbhASA/ylybznx7vcIAzqT70DylLRdGhZkHSjIFEx7M86u7RzgjDrvdvJERrANg+Xtv1i0O94zFx
Etthljsxs8OmydKqFW2biPvxEoqj3Q6yoPqBF1mJ7yYf70HcPr5ptraqgDjSuSfrhbAa2oKy2FVd
i65/A9oOdWr6XZEX1hZplVkzG3dfgZgxe1Eb+4QESBwmK1RqB0AoY5HHxLZsJSUFeL9VhSQ8RLgV
I/nJp3lqMeqwD+FNb76p+pP/igxg1++2D/aHzgQXEjlORQnzO9UF7Riif3k2/4YZwM9uNRstPFuI
rJITMlMVVPwVDQumC5nQWor5NBMiFcnGzWYu5GdZ/7us0qtTj65Mwkz/sos0bUXzFCVfO8gBayow
8gYH51mAP03D208xKYhFqAEL+wvbmDl8G+R7AMuDFqU3GxSnBR7Dq2sjxWpOP1DCnmnGyxLgTuLI
Kfedyrd0UsEHzfwGVSGbv5C1LSBFYVG29BQIZKc7xXI49uV77ohjv8Ym1Wr1X4Q2t0sCmcL9GW3K
xgunKjoebJCwR+AOKCdhOONodhYIt5V+OuypL0T0NHD/ebM3dGBr6Z8MMytmHs8jugZp0YfSVDru
U3aMLMg3E5MjdW2/j1PXo6/O1UMtp1addwCyWjQBE2kRWqiefUhkFBv6pGqOHfm89ozidMrj1Y35
bMA05zl0HJQU7CptAbnd4s9PWyYU/yDxSJtss1mI3VGafMdUVL6yBKXD9Zn2XY76es/zogfmVrVt
2Gj3Q6mwbwv5eyrza3Cyt4txeMzYVg74P2fmPtP0qf9u6ejbNc+jeDyo/DhJlqUt/aybmC7vtQzp
RimFBhB2IkCpRsibV0OLB2jMWgXEEprf7a7vv7H38kM8mq8dm4cevACuOoo3gJjWWx3jKYE+qKMb
UA6sQMsM6EuTGHubpSqR75YHwmvw/OROr2GLvtZ+UoYqupzODF8DoNUisBACw9gbfptTv8iHoFrH
dxoEWTFpYihqgImfBJeJEdxkzznkO8yzeCmLeJE04AiDBvCw4P2XPClkKAhA/udIs8fDr2+BoeG6
+QD84Un4cy942ZJxN1cf6mjuvlPpBYsKX8aIqDDl2HSr7Bzxp6nhy9iZQYjqDmiGE4lOFygqYrw9
JxeYC5RYW/OPByaL/oisVJ+tUND/WALHd2Nb0+mPaRjmC8uGM8VkFK6ahRcRtlD5l6JnASHiD4P3
rvgj04NqrsfgA8Eec72A4ILZEQuxHJW0qPC4NeC/bnR9b7UFllYh5cnsyn2pAYP/nO/vnx+Y+Pph
wWRVWYV9RrKdb4simtF6fLS9db9PsWqbAsHIUMMIeTT1nna52ekeFb88SJXZANdt7zaycndA1Wn1
ZEGc4bxGcOuefAb7XsH4CgNdJjU5pelhoH4SNm/tLjGCoviCvv33b2BlXn8DraeByLqkOziumUQB
To5MVIN8amSYw8Mked5KWlKScs6Jk+ZoDdDnQow/hb/Dlt8SHSmyOiWZl247e3+zU4MCVlZpCaJh
TuRrMrUmbA2B96ViJtjtHTi9U/Z7NvIoXaSX8DhbvKgfcR2Bgb2f/B/MKDkgj6cU9aQ51Zh0icM8
e4NgQ9ybEry0nhqfA7Wfbwsf9bZRp8t9EEDjJ0vF4G6hZ/q5TiqauCV+2lMrcV8KDKpbQJCEOGv0
Qi38NF9ZPg2DXTtM9tC1fzqZc0XLRBMuk5v3D3aAO8ORn8hjfOddUd1vKLBOCsQz6ybJeOY32+m+
bTEWe6QbyFsOQ1BNaiwyUrTJq+0Fw/TaQ04NcIVsbnzMYJLk1RPGoYyTtXvMYQ5DatoaMQ854FMV
P2+uf/NLXW3GEljMHeEcnaesxz42iShkSCOWWXqryURYYPkxZQK6sobFj+RmAkwSoAfrI4MXvjng
qpZagppmKsqW/mj+eYsxJoEjfYZxuSoRIg8/mvWHftKy5Domz38afsSUl4axfifderwU8gFkRYUJ
Ce+GjwcdqgbgImMDuxTWdPEvrhEmsw8wW+IQpZ+L1KYCsmsFmOZkLNWMKq4sJxRyW98pp6YMjj6q
a6RBf07suP3l5/HkjqdzqKADRf8SH/cqXVJ6xsFi40BFWoC/RjDNrZ7x/69e7aOzDsqngLlRme0v
jTr6Fr+cdTRD0kK4+tqqZW16DY8M/OjhgFbyuG7GAp1LNnEqqW3Rc+eYFZyET0tRrcuRztwe7NEh
zzJ2G/CnedPHeUk9Eoep3n517FsIFRyW37BEWYkW4+NwPcMG/cycEzUgsRRDT5RgY4vJprPyud1i
NQyMYviqvxPgjMT6BGHfjE1u2hJvHe+Cym5vtPeU5rfmoZ/wa2cFiUsbgHRI3zjJFPYIjpvKi+hg
Q7ZplsZeXcDqe5fNeCwiuHUsQYaoMl8/3AxHBQAlPhDgYFSkCIknsh2qv3vGZbiRyCwQeS2Kcj2h
90u9VGYYlF/S5c5+j+ljuY8bFdNMOl3rfUg34hwEuXrLvdZleJSEZ9GHJ9tL3X6/A4q1L+Ebr+0V
vgheJEpU9oE2+UVCRB4LpS8jtxSoCY6ae30ZoJwrqBj/Q6nnCTiQXSFKGDkOcrurLWwBIvFJFp6/
qXsx2Dl/eH2fQbfEPin8zLUXpoYCljtMXWkBx1yIpAmEFM1UXs7oEEZ6fzgb1yCoSWTZaWWm2GXQ
23A9j+6swhKVMwipi/NI8b/nWtM2gxZT87pIN9Dj7gDI2O8GsdKYv6f/LJh/90/0S5F2ubbul7Y3
htOxCWGwSbt0Kfbls4s4Ip260CObE+wtdctgIgc6o0in2WSs6agm8uS7+1jH653z8Zjw0l/vK4EZ
UbAYJfLYxCvYn2Bln3IHk5G2PF63mc3Fn09868DJBc2/1k/FGbBIiwMlh8pfaYtr/az0ayvwMSXY
0NRCOqgn/IL1/+74h1JVsvZD8z5iJxHnDtZaGjTNBSOokCLjY2KDaRxZyNtwFDKUZdy/pFJHoczT
Y5zPXkxo8oQ+LsbbGLIGGPCuqzejT7jpevzvkxwDqEHM8CDsnwK4MgrfUR+5TK69wdLzQwVkFddn
LGrMZGDICWeMaoeTR9fZiFal1zrYCkcLxYwBuG/uqZ8vfkVAYlLjZewAsm/TMBfm71oUBTo4g94w
goxpzk6009WsCxdiFvUcH4CEdDTNqg2rPKpnn2sFCV95XzPPoPvJN7Dq5JxrE4zeFO112WSeHtDk
eM/5mkGVmzn+z+FIl/I2zRrK7h7DLLU/V6y8fgJhfr0zP1YE44Z8mqGF63TpzNBXLiET4AAJh8lw
raTinwB9xCee8lMq0+ai37oe122xqwkW/ag+WW+Fq8uS6OGtT1T0ElP0s8Fgge+EDCn0OjfeSYYX
837QYDtbac6vIkEKK5CSjiEt6Jqye3TJ2heQ7NKl8PEdjHgzyb58m2gCifvBnMpW3MzA4xIvn/Ha
vWQOdakknSs47Qg0YH6MJ9NnkJS4YA+n0JYOqoQY3vv1tk14nNAJVXKSH/gJyF9HJmossQ4OYPFh
jrWrKdUPp1idjpZoVbnlkzYzXXUwsheutP0ROE4HAcXOuoFflLBVGcPqZcQgpJOsFRC0t7id7GwC
CHqnAaCdW0gxS/JpQfabmSoODtDBoO+bJfB1p1GSgG3zSqWBan1MNEO1qX7HqS/1BuJ00zfTDobN
hU9sXmRowMvOO5LrjsMobdthFVhKBcg1PteZEO4oLoaAWuSJB9xmWs/IisHIOZFA0RuFV3NqN9v3
tHLCL2b4EDMwctFUJAfsidqSh6elAP2VmvXTjVBXlC5uwxh8urTA2A9+PGR7T1vxCRbBzodt2RJa
7qtEPaq2NAxjjgwDzPdatFfFMnr0qphMIpZXOPoHoy1sodHv7zYjnXRe4hA4xDMOCc4CFADf+Ua5
q+6KpdBdmLKbVc5UEqVQ6UgGrFlwDbDOYs4GARBfp7d0pNoY8rLp1Yzs7w1Z37uf/KOlWmkvygwj
pH+mcpQGD5MpBCzKQmf+2eo6AFBtIuje8kjpqmyzQaSp2IIDkiASdJh7XiMhWbM0ZrhSwwl10mvI
IoITPmj47uGebKGUEZU8JhLQP8U0qOG0wIEJ30sS0i9/zH2oSJiZjLMwC6k7rQWZ5LIQXzjFfYWT
ydOU816anwsU8wuFkwJQ866x4lcOFxYt+6QzomX0BUrgLwCMkFflWjVnprO3Yuo3sFNPGrUOSkZR
hlL0Dc+y45XpBkAiwbuIlLCPu6Ble05Tya2i7+ayGQr37wtNASjC9lNG3N2jLIjyUHYRQRFEFbkr
e34KYoy4qDXxtLCqlWk8Bs9ZwPVoEUCyY1PAYwr+BPpo4M2ks5vV1I3kTjL2/EtRJVKGLU66ZqrB
pQS1SpCsXYVU2Pnux7EQjz+7Tj+zyizcOl5D6ngqfOCNKYEhdvt+sbyYQjx8nq21kvw/B2KuPsXC
pNi6ZfHeTWwS/LFA5ghh934IpxUCKlW2REzfdXeuGo/ULYTFwCydeC9UYnPtHVoerLcoaIWg8Hfw
lfTaxv3yt1k6T8Cd9hflRBi6EdSx21iuvG4+jKhltBf21E32ctxuPbDEQ+8iM1zi0yZnOnuy+nrw
x+L3HC6N7AdQUvGEv4rqIsRwtK4RvS2zpi3P5+avZJUktJ0VSap9/3ueKYgNxoAQjizaQ58RbDgi
sq4q4tB08CJZPG5D0nBugZFLMkjEaFaUQ8uAcay9zZqDft/afI3jC+NNbg1viXbVbLpdKCF7EOUA
kKrAZNbQZID6tqhT6ywO449Z67eOhiq3YJ3nZrYpkctBlFBDJT9Ko9Os6AUe9W5pS6yIL51f8D92
ZVr2FwXN81MrthwZhq7dPNaTy0hBmpCitCTxeVcGQ7J2nC7T9+ME2xqlVzDib6BAgcxvURcQ+/tP
lagVLrXIzLlaUuXpfM4SErLd2N7hIEa4wCUmsdHYzyDMSntpmnfauWMk+3C5cJnqZH/2DSjGz/jc
V1OifM4PiCwMUd5jZxPvFE/rFYEp3PJoacViSsYsFJVzLh6JLP4v+N1syloQar7Q++goS3c+ZUW0
Xttsx1fFNFabviEP99Zap/RpOa9lDxTZUXvZ5o9Wt1lnvUXz05U/sHbhZeJzYUbAuzXExTSZmvKw
CJmftDInDrQ584OsDvdFMvrK56L8xaqIjdz2P8b1z8B6Bs/wzxoHRYPkOpSFB0fUtnjIicJY9iF0
P53CJAxvKt0uxHShmbXJeND0wQWMtfpEgDcbY/PQuh7c6LqOMBZX+1NQiIu6Oew33BHrwCgy/tld
airs688mgOJq32oNTXwTnBQbQpyqXuB5PkZrqjB/bWi+YQmSpV3C0iunWpKExdmKIS6RL4gtnxrS
NDnYzVJ7dRiefLMxGiVUp18DY+syZ14qncmIHTBuRX7OZIWef5nPs9BajlFpKP4XW7qvEaX1Uecc
1omUmOQqrk6W6EQpax0mfjDxvJBtRoN3cZeM44XaxZE8TqckeeferKNipZUqToL6NKVIcXKpNJH0
Tsg9RjO5dfZ6KyBLMFEHTwqFvR9F5VKsbGVA0pgyH4R7iPQ+4Qqu3zB5utoyy9eM7VR3GHwGSnGx
HWtY1/mAop5hCycq/sxZQA/HH4luRWbnsMWQKHd5NBclU7fqG4Yeb0DcLhq1RQfI6n7wOsla+5iP
RPu+SDyNZh18qrQpqwbuNF26u5BeOoox3rqspyEVvFQ/Q09BL6pKGl7OIvIW7SYn51p3ITTcmn7b
sFT0fM4Adz+FQfSRuc+AwC4r3wSONqEdbQzHJbd/HHELO3sBzDKyM7okQea3Lskn9DgHRuwekO6r
pNjeQxc8ri8oqsKKXccVeILbK4gDUVz21cQj8vVh0zPJK7H/uONT7R78BKc+HdvxvFkoFIM+XPuo
EwbssDY4bDhVWqyAEzKaPZ40S8js1OdxHPGXZQsup4ioasFpDKRSvr3vs9IQUcSywcWfByM+F6E5
dEpVdwJo4MsBRiLjMmTmDw3gjGJec4G6HFs7YeljsmmzpHpP3aSpIlbSEINLrDIkUey5AaYfuTnw
BK/GQKMuP1aozGoHA/U8VnCPGRcTA/VGhDlINx+3CFse3krJVB5KQd24u3kp80jDd1vAIr0nPUyJ
EFjltkCiE4HA0ggHv8nxA8WQNZ5VVPdgRloATNVydxMPc+TlJWjXj0Tr4nYDwIrg0ibkt85RsSe/
vVQx77JVvdUwpc/PSi6yihfzZM7FbvPeHFutdyqPHOixgxtYnJlJoantVyMlV6IAoq0BsuW8VL9k
kSagSPmYtmVmy6ltwFVlUg21siM8gOd9vIRjkq5fjPzMKVQzr3/C+tw3Te7m7iyC59maO5GR3oMV
o30/o8jrDC0duOVITLJMZnGP3kI7s9hzHWqgZGvYTKeE+O3kJWkBOWgND3/Ax6cesZEBjqRknLZX
m6DWsta6T+SsInM9UnIdFMwR6DDUxIW/g0lUGMbks318S2yOVexxuum7gcjcuwCzD9f1ztNAVlXK
nVn1CnsARh2BMAt2cd1dkQkk+WTJw3cv92fZAmlmvO+fUHOW4Ip6gCef8aoJ5MJjao8kuR5dm2j/
r/NlQq/nNdjTy+S1A8FMPTzBmeowTjHdNKRKUDowVhYIROznfrLESUUYbCcXP6m3UHillW7hX8d7
vCmG95wlK+zG6qqOb5hBZfUO/9kaxFwDoBLCpnhdBswh/9ckYT+rDvzTs7+L4DMVsx+5HzsGs9B4
lolXwkTKtlrL2j4UtuFKZlKjmoQZtSc27+vT471hgXi/OvoPKZxhmIKOz9FredqLjOd9CmwkiRgi
XNAAWv7SPbfvXFRIbxkjfb3pmRtiXz75FS+VRRrB12SfcSHLn/mPE2uFk/sVQnw5b+Bp/FON+7JD
FEJXWiqWx05uTWx5mXVkPdz5bh9EajKozj7e8qX+0te1Cy5kSiLcHCyDZENbvOk/PqJrXHX7paEj
DeO4SEY6CQsc/7jCLHim6Rstjg3aoy4OafCBbkJ2MnZmSaUq/fuXxl6JXhFpDhD/nQ4NdF3VKm2X
fcRdputphXRW0+wQ6tWimP6cTGsR0a3MGwfpx82H3LWOz6KGlcIhZIEbetPbkXObsQ+oyffWo6aP
JRmQeXYq4O9txtP2ejiKEj856kTY2sU8o8+xbqFljHKlIf7R0MF87fMh49H5Gw/NTn2XIMrhPImE
mJB69Ch284L3rRs8Nv37AWGNs9gUfsr4N6YJy/ZV9Ba5jGVlN4qBCKl3D3ScG5qH4Fu1+IaojxBz
jPhLzT9CxcGKIARMN/Mak29Zy2VGfto8a1A6S9HB/oKrgFEhcVVz5wAWdT/NlEnhfb3moOK/PvUS
SDerTgsdvmz3qn+LfE3W0xMIB/U0Wt3IJLH8RUOKjUqPDYu74/sPZ4fLwgLd0+e6Zs7tIbmgJAUo
KRrKl8QGBViSXgS5PB0+Y4rf7MF08G+Hzb9I408LRnXV9/sdAj1bkFw4jDDpistAS4DbbdoMShSL
6XUBgu2+fDZ2DwbtEjBt/C6foDGXU4kA/aiW4zxfd5lUHwaC8DELnwm5jNvISCvFKASbXnOrajes
YxbZURRza23BO7sp2mO0RO4EK7/E7G+lO0RVM/LZ1MKLTZKxrr6r1F/qcVODYMY29kvSSSrCjqGj
Jak2B70ye3XbyrRac6WmK+4OPQo0A3wqpKbl5/GLpi71eS/eV8gcNOY7wwdonm3HgzELm67ZE0LS
J9DbtlPufBJb+mzfOIykplVMwToYAFkR44eEG/hR9S8ZBAXIlnL1OD47TvfL2XpkqTHZ3NPYX6DO
QOolV05hhwet6XgkXN9EP6Ubw11f1qetGOF0VjDnIkyJJz66NJl7fbnRfsfIsDRcOQdLf7Murb9F
HztKpaGQirdgKJqlnlvfd3Q0TvSOyuGQ+suCdGmkaHeCZJS0ElcmZa7sth2TEWnLXGZYpG+zKHit
YAPyReTAKddGLVZIoiP2zqudfoskcW3EI9cXvLaNW7wCS146xib5WzhQM4oooZ3BkSeCOdWGpEuz
AZDZU0ErlMVFfPz3AyDUiJINtocMAndSzwTpDQt7xRzQxehxYheOebecFvY67YO2mpXDQLj7sbbB
+L6Y+MqE/v6fUwm8bdu0nz4VuxZaZAcYEeJXCCVeQJ5GlcRwhQHLRtw7hJqmFXoCkQ9NdPSxikCZ
17i2CuSpxdPfF46W4vZj4qVzt0IofzS52RCnzvVwMry5G3yX9/6dWULGPPFlqarEnEJwUKnOMZXt
b6fyCHEt0pGqHA8tBWbzTjQCyS7fUlkGKdcdmR8hOpJrykLilFnPk36NgzmnPBb8gofJxOlmi8NV
dEcPw2G7BCMmI58dX7R4RCMJWO10wkGgnOog0baUiiPiT0iuJ77+G3wFGSzAeANJWjmWBaM9qPNY
nwkd/qNeLH04Rc4VbNSpJuTbBd5TFvyL4vKP2LAiAoXuejqNxw+Q1biD7wMt4gpnPVTakXardr/3
ryaxXhX0s7kDWz1G5HZivPBISuZ9oM23V5PeYMegmvIux+x2Sq8XpeEaIZ0bPCq8FBOSoK/AjPNa
tZ+nuHs91yUQf9FAxteIGIhtqfbG/1XxBkcdpi1qUQSUX9NRtZUs60cLiwNQ8LRhpNdSduGobXKR
Qz3HCClPdcbgDnCW4bt27nVh080ZydtVQJ3VBbEHnDnbzDnqexI5zs17b7hXBQICtMFTO2kk6t6V
+wYujsI73cbx2RQf5ZFJD96Ein0tORYRn+sWvyac7V/8sr5NrckNp6FG/pnGam1uzo9wuvYKWRee
sKG3hQRYFyA7tGCN9VT14kTDziLiJllF6koNLaq3iWzTswS9qiOYLYPjQijbn+CNaDFwvnllZIS8
6ZqODJ349bs66u88s9I8sxaa2USRKhuL5w+zgzRQgr9g3O5BxmN0caifAGj9E7DXhOX4uhCNFM02
9En88+lc8pB2EkjSIKe3FUCCeBa/6nlqQdfTmWxLINopy2gA3AagC9/0y8xGaIsBj3ioXP8p4sX9
Yzz3WZAaZu2eme5XBVa12Xoyj9GNSaGYoaY0s18M1A0d/mJD7YnqrDgSj3vj+Rbfk4Z7jBBkIEIz
BCx2/zZJPbWuceGFDFQzmrp0h6D50GOZyI7dtVMey53IE3mE2egiiXjk1KYBvqD10yAkQvwjpo25
z6XL54wzZCYhJD3tXqIMzDJG/39hiKqyHHaL8Plquwc2xZ1VyXVykgUGu8oRHxK7wSyow0ud8maz
ETAqM6ug8fFkUlK1Svnd+8RO6oBjpMs1pLDhe05yyWMP+JNWYWq21VACJinNlv3RZHG/FuWTWXOm
jE6T39AqjtVY0k7zgloZ9XfOFZ0QFaW59OkeoCKMLGVtsMvmHUuYnFsEUPxAUlGnd+Wh0dIUxXLL
xohoDdo5bpLqDuNySRCRoNn4rx9cL8dE3lfRzy2GLbhPY+SkpIYA8ZGbe6IdauU8I3Nk4C0g0NUn
e1lPYC+20FWCD39647HjcYmWSRMRmRy02Kut7wx61nuS0L5bcntGQ7sxExoQBFj+9+BfrjHf6KXi
7LNaQqea4z6elZ8jsQ6Qwss3VfEhWMH4FuVaSyKimCuu8y+6yKvLr2hPeyvFIwg5tuQnA7ykkvv9
wgZtuh8Wa8LLb1kn3KQCEhQfD9VDJtJdp6NbaEib2Q1X5vT2Hv9RbdwiNvRzZRTC0CRGSRKwkySV
dbd439qCcc3I3eulFncZzcAchgX1A2x46DM8RV4ooykI3E8Sl/b7VUmpH7e14AzectouXe6aIfxB
8diG+0fY/BDf5a1NJ8rziIF6NWZp5IxikzNZXRLMSXESNJz231xBspyUa6PULnSl8ypTTEVRyIES
iutzs7TFwTBZf/dI+6DBnFp2VNYWbyecKsVOreeA7sb0casg4TlPJlJhudTQTvC1XOUZJt98bJq9
/rwxpqSIpw0c+KVRAXICaoUcGkYCHaUX9uRdDl3acpUh8XbIHH0StdvS3GMpgF0073ma1OpmZl3A
hszYrtdIPHnH/ZU4kTbr1bmPDl4BZzAQsCdmROqDdq9RQzDbCEaQwRGe3SHpcf8d+lTjN4Cjuwu+
2/wZFL7dEQx7ToSxks+shdhJN2I+iqpSGoqmGgWBnfkGDvDGIETmDgdAMZA9qO4wyydm/bpMRt5P
JDZSq5kfmOxAWYN8mPns4lxjM5EyFKy3N1I7R0CDOpvDen93gD/VnBmKyIhdQvC7UOHuXHXowqhE
v34cxUtXcndPUISlIQ3lraTKNuppljTktZ7k2ZWUwQP64yUjPlh6FdC7BQKvlrglJWdzCnTrvi4I
t1QhCeLc253Y6UnsveIknC0NvA0Du7W0EjuOnH6H1NLqYDCpXsTk0KW7B/ZtpbOxWCWZ78EPHQ5e
IyYzY81epsULKDaG+2n0q1WKp+NpIOt0YjNeCoaNTDAyaFxb/eBmnH3JwEfSLS6gXhRMOQxz3UFw
k4KrPOINEMGSTRMrjUUo3rS6Jl9VZ+ngMejvSAJ3lOwsOyyIMuI6nhFvOy3rwivEIEriacaOfs6D
4fjfDiQ6wMmd0SNi0dF2AjOR/dwk15+W5taiWRwoSRZMyKOv3WJ2RkhboTtfmJ6JD2YKYhX0whTg
B4q2EL+4JGRimdYgPW6SePuR9jFi0Dxiu/rq3UYuTEp8lhoL/RplAFOcCP6mmqYWscRw/v80dyhU
hr0547bLtoTxtSUl1sxdZ3P+vclF/gAvEHgCB0LyZY13lmN9bO3vO6IGRz7dHsLrdrZ2WGJWBpFA
Iv5Yjh04vHLL73etZ4tHtO2Va3DKWu4FjPSoi69+DRNiYIJcnG0TLSq6ed/Sv3AAjXOnkeAyOAGv
w5sAs9BgN3XXFD6f0gFzaGD3kYinDEKq7NiqCI55aIps24X4jPQP4OOB1ThIcAU+87np4DC7+CEY
L/4+BmdNVPh7npBwNpAZxd96ov5GblVGKlSZAiWjLGPI8D28otl2Oa/BuucxIOrRuRYoiy4nvK3a
VkAjA95+zjhb/DgoROo/GNs0lC75sd34aairL0sIl0i6jWD5DVaCTv25k5IkkYU/r4qyTE4qrBIy
YA9i6YwqytExGefzGyeOQUKyQMXMxZ842dXjRkH1VelTuIXOYe7zLtow8TDjTW9r3w7g0wl9ONvK
tsA/vbSWHI9yV+Co2sBqFuzeeypGi3Od9Iip0/qjpSELjLyRl59wv5uqeLkB3Dut39P8h18xnVHO
ISubZjQYhaX66edSACk1JVr4qC9D65DZtul88ZyLpZv5utDDe1AhEB/JJYhD0g51J0fm/XFaRUg1
mBpv6tPtnUBBNKOPDN4tFZg5XQeC6HnoMkFLqFwMonOw3zrIs7GQX7H/6Yy5SJajk38R7d14SNJU
JTp60nJgmO1HxF3Hfk1c2uLQ130FHDFXydPeW9O2wKfWzI2Dh+SuiyZLp8U2lpp8ErhLeV9uQ2zd
ixpBoi7IU9U4KO7jCCBoDmGm60EGUBVbBx138zxeDwgYZjePrKNfDE9u7ftNsxd+vFTTNkeVP8/v
qlqnI2l1ORVkLUBym/nQB3MQsv9L5BVQmLYmXWLLhcRdmnFrN4LVFibpX6J2ByhEXsSc5ojJ1U7X
15ToT3wvwlKjvZ83Pjvo2CqvdmVJ9RVsKP9nXpUkUkpjSSXlqTf/k2biQf1wkcEixXBqKtBu5Dxd
DN1edXk/VUzBzI+ndyURmp//FppIFyJi+OcLCPk4xM3fxC4grBXwdwY0qDHCPhnqswjsu14V/3em
SYHxHw9XPj0LM9tpMoj4SNYZeMRWFKWOo7CAG8Ch3kaauXPxcZ9OI6wy1A+QHQZyq/lSDZQqMBoA
BGmaJmsTtEpaktc1Itqs8rEZdOcRkKwxyUFsZUxwdkPCAuEv/Tupnzoj6Lrp3UMVv3JRVVr9gQc9
aR64YGAvqy1yU6PvJ5wyMq6pHbYo97ATO8GlUec9kfdiZU0ChCUPcmpbYefss1xyatRC+nODEdDP
oCzRWk13msOYg/CWqdJ7l54ma5VfKv1ACDHtJbxxIQgVOeiYQihZNPFjusXzjmG7MK/nj6pmygQv
QHVr0GtILqy0h9tdyRdgvc1Mim/RnWxBySFiYLk5hdDp9hj39+LNA74zCsOwCZkEwjBtaMgqTZ8n
PUHK/9UUwL1SiNpzEw6NaDXcsa1SbIGPhfJyE6rwlzaRYaZOn/zWoiUHLROfq2do0bIQWgqtGiwV
jfEN373OJC75bgG4MmOseUKvx6+zeBkkxiNFRDXkGD9R+BsevUisSwZvdu9wWU4XB5q4TfCNT2up
Zsjwzg+pwyuo3YwBILlWrxjhpn3HycC6uu1sr8yBZgZJr/RuJFMWnoVOXUGYSmnhUknd+i52p6G2
uCnlvPdrH1cQxTMkKwwFijRn0ua6xVRlvSuTaGhZHy4r+Qv/kkuQgpYpWRskoYKrYWgH1cIjyTDV
2+o4xVb9xA1nyTYDSI2tnZcBYUJD0jRERgc2dUt0187dfSfdjgFSJXFHSDF7s7HCQ4uCQ/8FKDsV
ujmtoaInGViJsYSQNuzO60MYRIAJHyZRVy62O3nNt444DTwBrUmbMGR1hxKbqTFA7FE9qkPL2oRz
VvX+E7jQHG2RBm4qom2TSXb2BeoEjbmazCPPkmlHzlVOeNOjOGKWrY9cJ36nujTZnunKwSbvgoiQ
1rowCkEvK6vfUhiLONFjCh61o5jmcrW2TLcml9bOEz0Ynv6pvOOPLGRuARAjz1UdWRxiuLUW1E8G
hnFytggDQ0aPE72dG3CrOYh8TnV8ZVz++oxmZj8jbw1Dg1wDWUJ3l3VLLEpyWtnQbyBEgBUm8Z48
qSoKgRj6YlRyiHrgloBTFs+sFrhlWt7IvIArzpGJF17cftW7LC+djs1i4KQE0sGcPW8LNQxthYrO
vtU/6D+YTxV9nH4UCjO/HgnxDQwSG61OMOYPUgy76JZZbcTLgYT5B1CDueq2WwzV2N6h3MNPzhn4
NspBRwZJeU5Ckk5Xw/zLvEIFu1oLQwbYL628638LJCOFQIswcDMFrP2aOd3mfgRUxQgQCJZSlOOi
XY+HexGAekhDdbr8vsxFZFY2nQ4reCqI3I3VLAic7TSnyNpnwvcNaDKsPmIoiH1mbiXF4Canpkgs
FYtSZlqouV7kqAaGYv2gcRG+O9ILI/ggjB3CNzNZBggfBolVcT5qBHHp7BFXhyUZJVoXld/W7HtK
iFUTRTJbKQUJEYKPR21BM6FVC43BtGO2A1kuWnArBPk2cVsZFJGZBVI0c0oojpBIFR5b0BW14ASX
K7mchtReRacnMlddBZk1xJBrGMv/2lQ9BM7h4wj/akFrzFzEZ2sVYz9+hdCcAWprs0KxxqEEVctA
Lub+/RcIlUSY+eWJQ8IMTiD+OKMRVCNPgnOTw2G3MM4gBnv3n4sRqiDNmkSW5vVXCnI/yWmwUTy4
CaoHUgLDSkYpCk/dacFdCt/RCXewoUGh2wadktc7qhavJR2NTdGBr0iYktA/oWShn7wG8gnNRsjK
OVtQPZ1ws1lgL/2HELygxxrliT8inVttm4PPvOFS+McXlvosClFkZtsF2I5XjU9GyNHdnhGBrzAO
+8Kblz8B/o2of+oa8xuTxwZLdpNsWXM0HWJLXZgb7gtdYVwme5Mr6ZmrAB6bq6wXM+OgSmNx94+0
KBR0rG+KOkGdCS0xhqp3pfjpW0TlFzbwMamuH5RhiHfVFY0i4AutnHj77HvsYdPti0Tx5qNesovk
p51y6dokyrY5smPUmhKRLqDiujHp0LXbUajCTnJtpKDr5y0MwBsHxeGSH5HykBnHFWuSdHLLsbhQ
6RD4IOAJxp1f++1e6LmlvFGw+rhU3WHe63IXdIjhs816baztm80nmRctcivP7k0EO5GRcs8uI1pZ
PTxDEfLzwcMTiJ9UOb67YxPvvTVsSMkFXPR7QUGc+Kq1q6M88fOPrN4RtUso8WF74+ZTfPpARaDM
kRYS0RQVTJx0K6QKFH8G+dto34Os7xThjwdiambnBD82Fn16PLt0jKIbaL8pNLvSMSX7M/VF5js4
6l/G0R1CO4TXKnrMiXxpWMnd0Egor0saZauRAfwCf5OjIZeMb9vPoy/W1p6Catb0CMckL1xDviMF
/nS07oisF740HM0sQM07NFV2OoAtC8sBcwPN9oj59hSXqiCqqII0K4Ao42mTsh08ngvxDpm4GcN3
4wnJbY2xisL8edOy0KNjDAOo030dYxKEc//qCQ3WWVxi42pQJCDuxyfrhgTlEr5KD7usfNavsczP
OU5+LHiHTOFKaGZDcGZFkqM4teAUYIeTGzK2CkM2EtDCibaw5txmFth161M7qUb7tJPd/Yyiv3kV
UbQ33dgFzqLqzrdDW0Xr0iMdtwCWYBTbuFiQKG8DGJgoEGwNCRZxjrDdEkqFuBHm18kZs6ZBq2sa
lz22UxpZ0WAN7+wvQTcZvdl3GaBh1rpnTV/mAgH1TjprBzYm+bQMSUeVnDKGvGyNH5aedhIAymaX
cotLGALlmbcZ02G6tUHI4qsLel60wytjXSPiy2rRmFc+pxh/F9llQwwfG5ojD/IQh0piCTQvZD28
FmTLbHLI1i9FCzKkJdDWbUUzYOY2N8lSX2EBVTHTl4pogC9Qcmve70EFH+uy7NQTBwgPFOiDcRVZ
0h4BaiPWWWKeeqboUCrFoQdBWnFe2L2C4UG1iSo8RVlQsFqfDN/q4FCjRp0KwFm7pNUaFuCytgtt
L0EIHeorO7KxrP8sHfCOcbO7NQRoodO/GXRyLD4SdnLkDhYA+1pNFiUxWHCqY98JfXAg+59xHN3j
5MH4uGzpILso4IqmbxWjnfZatJod9jDeuJFYtKt5BUkYcTcoVX03oRYBus21CophDzE5T3YDPVGU
tEJvKSiomZmc0Ps9X1mMG8WhhulvpxbMbSDQu4mQdnZYrdXb721CN4F9GZp9C5YNomUao2w4HS59
dzxXe9qnlLh3rL11Okw7GazQ4l78IOl6I3C+/N84C4gQpaS/HB2e5sEl6rOwaDmFMGSnie53LdJc
OWR2XfmTInxBUrwywPQTkp8MFeFGFiwAbuKDkCkxkJr9iNFNs6BxhQeJxKLqISpelg59vZwE1iHc
wahxYD/WPVwQZ9YcCEjORTb7wf8Sf+TRdPWJzi3ameM0+JeMrc7xRRzxW2xvBDEkEeA/kOlO4hJp
LCVY+iIIh+j1iDiGwvwMQHyQPrY2UvIH1yncngIQR8oUlj1t5PV5mkiynqTcARmwO3tVGLi1itZ/
0uuHOVG5x0v3wQAzkoNJFBUShnnwnVGeHuut4gx3/NsRcvVotyNvqCDkqdJRkUNayGc8DlfHFhYC
v1TZj62x8vekO/sA6tES9qxZGI5B3u+S8jn6Qz74AW3br+49FKaBXP/Hp92HukD03Mrg8Ow5RlWv
I8GSPR/Jhn+C40ANFG96HHWb+s4rzIHA+ms/qV739r8WDNLRTJcjGOTYCKqrG3nc9ZrJCdYptxOO
GDlP5Rqgo6n1tn2g0fO9lit2jzb5Zxa3Hnk6VOPV3eBO7wKDTYeiapdPmK1uGm7iUADwRsEf5bMO
U2IAJf+fI13OLpQNYl0k9AYG1pgm1Vi9XPRZpzrG0XhZR+Hllo0GgZiHOaCXFejb1nqLdu5BS4f/
YqGm663dsmXG2vxHAYuPRFrVArOxVVJc4FNiGQQEdngm5FBMedg8z0mwisx/6vyZrGL58g2jgNe4
M2D2s5kxfpwh2zM2tApvSBDRssVFXr0aADEuvzgthK4coLLEV0m6DgxNaUveibOB1kELE4WTSwxB
UPDUE28GUp306ytgtYZ0riJm/wuHYQuUvr8GAsdjv9Wy7VbkUDAXwYkMB9gysXQDZ8BvYN92v0ga
IZfugMFZtLzEsXOXTnJqL1J5kq6pXyGqUwdwtU7uhm3AInwhbeqOwquT7oHD98PXKTdDds+GoK5y
EONyOc0ahpzQOo9EobgHGpw08IDhmCqVTbQQwiaSZZFFeEuLTqNU0QLnlP2hUDK8SLbUinHlBvgB
bwvn4FCmFcVfwUgGd0yF1n31XIZrrRqavn8MJavJOQII08x8JWYeaRNOHaHp9b7NoZcQ+RlxkJnk
/P5yan8sW+9PVqdpOi6kVqLenHtQV1qbU5iU+p9xy1+h/0mNlCj0JSyaYfdcKhjofhbqMa02dclM
LuPBEOa/V1ehhkqokjDyOO4OPHlkRF2LKvvMTC4/5oLa/25w/R+4yPoJagNdoubP7jRXef+B5Slj
FIGBF7l2XCdATGx6/UjO9TmjGhQigYKBmP3grZG8MLIgcdKjjTI3F1C8uayJswgvEKXT1SVGWJV0
QgYbekx0ZlgJs5qmklE9O5dWNoI+CvQ6dO0XaGAQEM8QFwkAEBRZ8TNVfFFcA6X6l+Y8zEpBznUD
wB5AnPVf3+J4KYxADqOIJTJ8wPpZ1YXz8kaBwODbopW3kHo7kG3VI5pmAVDbZKktRUi5rTQ8TlI8
4uLZefkVhjJ0jku1AkH60G8gnJ01MuK52r7N/K377ZtNyIQ9OsOkLtXLKkXXFaRzr0X+9Qckqkhb
2/kuTJqFB1sjnUfhp2wgsv0MlgXFjp6eO00c32w5OK3fAvgoWojKzdnFDCVJkL2+CLcUCl3caa6h
lES4kcgwJEAZ9dLCUluSWH8ppONMJuCz44vc5M9Yg4lapGyxXXq9vk+gfBSJO9fFIMRlRXpm6Pqd
yE/iq+P9zduy5pyJAiBp7/FL+A0jy3EawAwkeFZZ5bl1XxK9aDOgBNW8k33qdpOlQu4Qc42xAIzp
nLZB7hY/Je7WQnUrLbyIvlFRbui3kGiBTIXZXf6J9LCvDHZfHNnUkeVUS/HGUJk1q16SjpKB30Zm
uNqvdacacR8cmkdMplFDljctRqSlYk5hcUObSGXF/e30tIjU+QsYPcxbzCMeRCk3ujcGtUOlDWom
FGuRJraPC75+ZrYD4TZScy+Jf4TKvpQgDWvUqq69aYmF7xMa/gRKKvXzvCDqyloSCGh9z0Aw1v5g
q9SRg0bpDfVMPojagFy7BlHyQZGcWZQybfyFXsz8e4PSR2MV+ZCvOsUUOezy31bdn19g9EOz6QWM
5Ubyqq1RtcjQPLc2mdE14Auil9YVcnW0M37GnVJUYCJpTct3CrOvetHid3m6gqSSQYlXa1dqtANR
7rpvOzsZE3ULcMBN8AMa+IQK+YrCDyweniJzirqmm+L00y9OT7EnpjK7REQQQrl8voKGMS5TjAN6
9uT15b+uoEBLxN0p2YRJzxgWpUzJaAmQ9DNv96oHLKnRHSIn+9v7b0F+fNv3FvfGrrYXJI6gBIoH
ekCdcgzQwdfunxdJflHzPp/4nVDsMhftXFlxSuIzUdmKMvkoJfR6DQ1/wpkBDOOIJRpd+l+0jUG9
WUPxz4ETJu2WPKFOfJytBhz9ClqjhxW3iOsxf3VIBuP2H8WknxHNdhrL1CxLLvAsWmTx0jJODlV5
s+2ZFzsttQyZdqgZsv7226s0wQ1Pxs4quVEwGTweJaLwkqLLKzALhmtw1xoz/0BJsJ8M30Gwj/Kr
WChwVoFx745LB9frC4e+wJ6i7C9Px4DCLmpWMtg0Ro/16/AKtTIiCvheDksZ66CoZegxQrDQLhYL
7zIId7UUn4avTbuRSa9N5dHSaQEN/q7Z8xK2g0Xv/3G2MOIAjyRPUt4jf+HNTRuT3ThjQFmo9r/j
ir1Y/hhhtJtc7xetebrmVHwb5ELnVc2Rtk3a6g4buvA4JAGivDynQJuoa0VIYtkIS4FuGX9n01IJ
fd2E7wgqK3Te0pc+sxeSe90iq1P8ps8RZXQmNw28U8tQQdOuI5Iu8S/oa+/fAzDM8+d4W6RAqWOz
BfnNAk1yBRLsXSEToWxPsiQLuZOiW9ut7O8bSIDQ12MnP31QijP9+Ep3mOd1UUV6WEAUNblVIlqe
8INpRMi0QermdB+Igm4o8kDBtAOSiAhD5Pg1vXSfLAx7kvJ75f6yTmx9vwrp1EWqH576pCzqt/5i
wVzoFWAAuu5Wgl0jbFK93sD2nXC9UN6/WDVqQ/7okgIjmp1X5Gbv3yoizOiYcyWARksNhExtDDXP
vCT5yEepJ0MUHC7Wr8936VG4+NAG2iDkfAXvmnUpYnB6VDBMChZq8xHSu73YMz6JscDyyebL6hZ0
akv/dvEonV66iPnwLl9tW0q4Fhp4InQTJ3SxQREL/gCU0EdWHMbCF6/ITgGqFeMmeqiFogEK9T9b
T4I4MRATPFs4uDBhKijGqjwAH5ONpYap8aWA+ncXlLdQdDsB8xpYvsfPATRPE6I8SQ48wykC51/B
MxK6YTQ5grnzVGE2jsVT/8RnpzRrIFgzaqR6o6a2W8Nwrr5IuaYMWVy6JdjmkohuekQWM3U0l30g
iKj/k1pZ0UjTMtEQ+UrceXcF+A+PhJbNrMAUQ+6bLAmhmap9G1Fchy276izFiZQSQfVK0j/zu5Qg
cvRFtwnyCHihgsRYqVNkK1DIlLeGF8OVLkwoukIT9CDrgBEAQyvFcZKv1cCBBXOjWub/DM/zGjOA
oGa08rt5nKv0ZA+arLbDLx+zRJ3/IEfmQVG72UILf+QD7K1WJzQlxf1kfoan8cFa/i4G9Au8rLEL
byAR6VjXmzZlIcY7SIhYZm8sPaO1wlWOSmQVtNQg3EVPU7iWjqfOI7EV9UTLw3SlqPfv9eOGQswJ
B52OQ66Vwx6FK2adpicfXajviJEIykcNDFfo6AuCXVFQ2SEkuLaJBDl27nHPt+uxhApCNzhV4D0z
8eB3K6NzYsM9QOrdHAeoXlA+l852bYNJOw00Hkr3x9Az0nCPw2Qs7m/t6JbGdTdjJtQXMFHyttvd
5arHO7KAWyajkWDzOhSXm/b5LqSe/2krHUeaThxf+Z98blQub0goqrRJpy+HJxKtx4WDGQcKErgI
wAhujwjYKmzkqY2X5Z2Fecz4yWjUhYAahqSJ30LcWdF+igNqNNhIfrJ2tHuOeiV7ajDRSdMll8yG
o8DTpwsaJwGMknHNYryAvUicXcNLR9Rhx7EFOzbCjskbPBn+ZXWc+zKuSuUED4qLQmEjrx1w4Itg
IgQlLuVwaYZtnepCEZT4+8+YLJiPm/NjQ/SarZ5ZeSvEffcmJKEvhbOeign3BKxv9kKhSv4QnTtg
sfA+IVCKcfTVzW4BCsK0VIXBNqzTMMW4zQQiTMB570WA98zZ9OERi1k9bXwpsGd7fhHLv39RkE9y
7iH/gO3rafOL2wEhWe67o3Aq73/JzKMuC28cSSxRcg3tAiLVqbqLKhufc4pTvG8/3Gg68HHOnv1D
GK5vwTG3ua6UyFQqra/actH2c54Qmi7I8cM79VIU1MuksauR4cnp/PDjs/XIVaDohKbEtTZi4t+p
1QiwaAhRX6xWbNQ1VEIRJuR9xV8vqPQW3tIoc2n4JwHvcsMMNX87qpaEbohq2N1vsT/uPV7xXGoQ
KcZJfBstv84idwK9AEDkNK/1lfsLHPIaFKDOPPmWH8RcCB5Qv6thsdMt+iD/MiKCh4/EA/uOHlOe
OQXqxukVypN0JAOYw23hqHqCiN2PMLYQkzX+dmTeKva/edO32e9O9DsbdKoxHJQTH6cYYMSxbl2M
McdCoxVrj6p1jyaM8/bJxUPOpAV7qBC2H14Mwj9qDXwZxLbEWuR4OorVubITUlJMgGnyrpc3IPbI
jStZa1iqaHky49aokofSOzHvFkjiH4Ig4v2fm9T5rGsU6e73EIJ3IpfpVIc3gC9MnDT+4z7nFwp1
pj+dcjLQ8ZCcnPQULeeZECT77Bjmp6vBSRloKu/UlkoDPhyeCKGVuxjWUpKJNuMeWMG95ITlthof
p6fJmyMJA1rTaIy4jNbzE5u9GPcZLJrR+nH9JZrLU8vVvtAITlmWZg/QD7TrxoAirWxo2ebfWCvQ
I2TVS6TM4XxGZUQ6qxfla4m3AmpSNCz4YY+UNq8jRc6gaS+8M4cYHwVl2+XNe6cbyIgTb1mdHtBo
ZzKc7zkGjjsfB10fu1cOQa78kKDmtHdjRQcmUJhHSfPobOwWZy9ss4lzqMtXi1FaPf9KllgSeIZ4
R+lFCTp23bC5LF//ml5wR0hJj3EycsQEwiCZssS9hyXG5BeDJjw3ynu/Yk7QFJP/srtqmVfK7/QJ
DLrbzCCJbRzCeWC8cHbnK3jCjc3aL2KM/mmG4swhwEh3QKPSZd7AOKXaGSh+hZG6gK5iGIQ3DmIY
H5PXiC5p95k1kwo9Jto0XoQHI3uRE9UCoKK6/CbXNTtgtfztLpzoMuvtSLrFJph0jf/gXvdL5qNy
itBMf1XZr9AHkhpf61VZpMCOsqgaEhlVpxKBT9/I0g2bGedOkJvmuN6Bu0QReZkQi3su3UdmvNya
yd5vNC5CweXWYdavj01f1Y2mDdxWYI/Ntl6zysf8Oy35T52Vm4ozFwncgJmKn4eR//5Ki/q/FjS2
ZZ9Vb3nRaW8Hpnm0w/JkhS+fi6H2yRFhkICNN8MxHglvIFbFxO7Q4QLSIlHOy6RwOIyFsDG90/SS
402TmCl0/4NzdvyLEnXPbo4lplhQttZNSTnombNeY/azt/euqlVSCwGLxL++5t5NAgXpGheRUM4Z
w/GIr2o4GS5QObjmtUrbQssXedNaSSi0Zi8NPl9+koufwzNOMA8o2c1a0Moed+MJv3yLrGZ2Cs4J
32igWyK1naYQoC9LCRBg9UrMTMWnjPbaHFm6utInBLskdtcoIiPNoLLNnM5QXGHkZs8lXtNlwR8c
7MnfMdINQJ+vXKDtVu2liD+bNaAEU2t2mFMVE+C1UHcONEZOAlGYT2ISZIXm6KK/ityBdQ9gnhk0
o6mYr3lNbgVEnj3EHAlrXMgZ7oKQ7Bm2ZKm7i/WRsf/3qJHfAgq8aW/pKzZuhFBjrUqY8jtgBfpA
gRpmYSo/Vx/9cq9eJ2oWxIEM7qeez9K/CRM09wwyw28z4rMXtglEGSstVh3V7mYSKlptev5fXyHd
E80wUhyfjweLyRCeJWGvr0xF31yEkPZA1wqxmTRJGGvTbABfYxsqaAyR7LqeifaD+ji9oIXDb0NR
Toyk9ShL+o12vC6RtY4X6Ikk50gNG8zQtxC1/SQYL4Oc3EqgObOAUM8TZ190S6JNViuFCFhUS5T2
PwoE5DP1yi8YVzf33i/sQ6ngAk5p352lqFI9nv2FeFoLxRUUv1OxknN044yTs4SAEEgSZBEYtF+I
nRJkk7J70+qZQiOkCPB4UuZoBG2usvKOWjCGMLuXoPDA+ckyj6O1XzW6NeDav7OuQR0/bdet8pdV
RMj3wQDt8sN0fvwxehLtYIT8Nel+1uzwrF3xbTrdP0+VdCHDysZlVU/ETAopaAmVaEBMz+ZlfjiG
fZ+kiykWt37cGi3lnQRAie3ZVVd07V6BR8Q2JPjrD4OdfALjIlB6fUg6VQWu9rYOQTFHFVf9pYQY
UwK2qJrN4m1/USV6XkzfSobnbY6pgOMHgG9qphCmIRal54Y3iriJHmjusUJhTMubwsEqosuAFoi0
g/6vAY2ZxXzgn2RTio8VudSLL6mcOoXLvlA2oUZHEdznaRMkwsKsAxSsvnyaoFXtxvJlpaT/8b88
MXv0rMKNeBCLJ++lxDUOmRRGyIwveI4JHR3mOUZW6V5XvBKf2n9R85U6JYzj0Y5XT3GiA9xI4zLD
P5fIQ6Vt3AZfeUKOooq6zr+hn5jfoAZmmGe8WPw17lKEbkn/Dl6l+yuTfdSIHuP2GTYP8cbt/Ryy
vShOF4Z0aa0CHekIhp1k5qxpt4UT8x+InhNbVMwDfi0gbnGZES+EotEMKE5/rZABXR7Hc1+yiK5m
v4BBGELrr/LgKy+RNbYMI1Ba0TSUdOvB1a4KtRzE1C+Sx+neKSCh8gSfpz7uYr58XBe+rBr9h0f/
9a4REQmBXOrjwOSe6sSQX4iULiVjWlF/+bML4HYd/vhLA7K9GKR14YdcIe2bmrGTfhGGFOERoIs1
UooawPDyJJQCnwAHRBxtnOokZeTdVkcr/mCAsveSybd2WZUEfa379MJz/uuZWBKgDhlRWJwMbZX9
BeGes9NdT4yB3VBxYv5yc+v3OigxOmEmZRiJ7VjcJsVoxNhDtD0UP7XzspEI5qG/omJ05Y5e5a4J
2J/RSK+AHBpOx9K8NpD4c6uyB5S2Idzetwox28IjMdRact2YMgKOGHfdFKjYGIODPk8ZxQ/dZlD5
7PWLEFiWcSc5Eg/bQVETV+d6Pw/Vq76406/tYi9Ad3KRhMIFg6O0xeQdIFdb2oOSOamzKvg8PG+a
kDKfANjmhmXPJ3Cl3PRHXOlSRuN9VVPhoA357SbianQiJAcyfvduRZjjsQPu9e9rg6ljdjf6NASz
t9u96gUh/KoAdd8SFQnmNZb7k3cboPXxO0gGvupz4CfrJ+Ei6zd3yjpx7lyK5/EQjAXoSDBDvo63
cG/jffny0RjXUClZge7cMyNuWkQ3al5dUZXtLDWCxwtn1i99zgR09T0m1xG+rfU5CvSnc6TlIP3N
tTIlR2STQ8eR6oXp6WQdxbpWgw7vhUhoP4rGyltYvM4ssJeBjP5mp0xofDwncQtnDg8Ez2dBeNUQ
81KDPmoU8v522BZuXOE/aPbG539qX48cmp+cIZxvYH4nmyg8ysu90/YClb+HV+UK4Vy0llcqr97C
dmTJuKSqdMS4W4XpRkmNODiw1Z/rZ+y1XU7Uj/zSE8UfmNCPn+RvaO4r5Pa3Ii/48kF4LKQuG1aK
Z/Kv0gQD6DSBQnlDjunQdKyxuLD0vg7rHszoJIJz6oYif9ngYvpmQR391FsvNt0BxFklTCfeC8Ot
kknpZVKQ9858ZhAcys5kFuRH5GNlOeiwrnCX4dtzZG+Ig9YTP42ky5iMS5LWmdaBzJARIpyibT64
t7bgsdsRxV7RG0id2Wi/Rq39odoJaFmZw6qjKaVhFHJslq/phvXeEB3NEACqTpsmUUj41QwZPRLF
YzX2eaQ3zQZGpD1Sv8IXAC2Yq3fKP+HwwzUnhaHzYJ6WfNjcSnSPXx8NOe/AmTnj9gRz3ebEzJX0
ehDHCqshwbLYygrw6ZC+p3V6gIzYVHJS+WNMiNBDJD+OWr3znqC9lMYUDYjj0473hCcIMhmTqUWo
ixZfCOgTmR/4dLc5HOhXhYpXHXX1CAwvqJg5OskZ7gCcDl1W6M73HNGbxhsd0ZEhM5Ayr0053o31
QuxjZ0goVP3nONQrjYSL3DlagoHA2DqBburtKsR0vK5mOUUiYmAnC6dpDASzBuhzfB/ECfv/xJpX
1GEaIBAuLeFYFDmxCVXC2Kv+kpDHbIm11uXBm4+GmcqOe/f87DyiaXI87Z1wO+pzj+8SwmwLTz/z
frL05uMlMdbKzI2ZvHkHXwbXzXAGvX9/zQJZIE1eq+2udG/Z7bwvJZzrTqf8W3Wj1XngBKofBh7y
lG5tzJsnwYnieAqsouZeRZgyewbGrgyuTr1R1RkMsiqvD+wV91f8LRdx8qd44N7yRqQ0syEAq8wj
YBInRjMgAEVqBxoPcvSX2x+lG38FxXQtLHxoyv19X/ObXy1p7Lkbqb472ZxdVQ4MtjVJ3+k+j9eG
OagZdVrTbjcKCSpfPx/sLsSAWpkxFg24URucSdiwBpgtO6fcBvEN7EWTyJB34i5TXNyxMmE+vYtI
nloOXimwj9r/WykIE0Jg2na/QOJkKFJtwTpn8cp0gFqtN1gPGLV/URLul9sTOB+uaAMlHUOQ/fzQ
UrYQmBxKGOkGZ5shw+ZsHkEMhrJATKd0WeNu1tjkHfphOyzVvTUpfBDgRjJwsqLcv68nfzECXoMz
bvXclG6UOvYQSBmmU42SWe/zfGnzjuPCzvUMgVNN6mAoG1YL08pS8Z3vkhxOzhQ4snvbMOL1cmUh
MeeOzTxj7Ci9iVfDqaPGCgCF01zz/uQSS88Hezs7NXYY9tU8ocsfgqRjd4cAcYhzbccuoYcIE0nZ
uvK6Ba4KG5s/VNpqDap8qlWSICVKzAEC1CxwX9CFou7lZGIYN0F+KA+U6UCMxKoigw+bpY6I6P91
3ha4bZf+9nuRcsiHhMVU7Sw5Pd4gI7OkojKC3PB9fD9rNO9RB30mGKgXWWRfd3mewQnpPb5pc3z5
v7xHLMoZe+BQGwqi2M61nPTWGc4QMuJ2bLCHj060dcgW5qzLQL2jBh7nvJl2XnztcRhGQzPzeFnL
28vAsiTOa8fMQ/TFN+WN5VKjcrutXfnVZ1tASlNkvJ5G0Nj8SagpY+G+guHqVU4tqzDbKliG/fNA
1XhJR2cryBkH+2xY6wMFphZcVZa3ItWEyT4zCMuQEMwDhMQe+rkiZSNJKWLmgWNwsNkgGjzzI/d/
+djUjfdkJgAvse4GTa0H+zTld7HTQRZzjDJtffFBGGRPacTlGdVVRYKLcuDn+NcfaCTfpfq6fL5v
RbK7i3qHGs4oTvPLB47nye8+LEPC4SjJQM+YEzajK00q6Ol9dhMassgWa8qxDhENtnUe8abIm8sl
pdZqgz3INkYY2aqiVW8tY1kmkgfAJFhYGRznybfdpW9GysY9d6shWM/N+oGhUwKAdlbDScQwdRvT
DQiXRosbSmK/KbNg4E/fniBFOZvDeR84aGai7USksTJt+lECM384Mzq0daS0c0u2KUuY3aWPkwDm
i7lvk1K9LFNj0uPie8r/HL/54yyMgvHnubbPzVlRYnkEScCVu7ykg4XXKdYjw3V14m4ReMboChFk
35B7Tcm0ZY+f5DhsLjzc6gWmcx6HBjqJs7JqvKWTW3zMrl5IpzmpbJnjhlqfPuPgNNogZQCjx4pw
/xElmJCGN7FWPrYEEZlKwaoUEkmxnKwkXvm+oe0I+Pjme3bJTPssiBmcmIIxFALQoytHFb+RU9gJ
DVqq9os9qNp5xXVtwdxAzr8PuypkgMt5fff2zMmEF3pKFa+Nl5HY7kcNKAGZCL0YlNTTuWrnBkD4
VptrI5urHNxZg3yvQIT7eecx2vMv74WhF8LwiLJ2oS5mF0DPybNIx3NKXR/EAblOeeTw8ezpF7Qp
c93c50aZjXMx56TQJnSm2GQ7nmxbmzBbpnObTv2kJ5C9QRfOKflqbZkPj1nkR8EEaT/9hlFVfRuH
TkuP6MRCf9ueJYbb1A5o4MykGfADbROBr5PugP9LI1qY58n5rA2K+Etokd4FY3Sd7qreCq33M4pt
vLaQ+KPWWYobll/f2gtNkYEYr1y6D/4dcXaV/2j3/EBvxAMHT8VvSwrdx9EVtTENkxQnDnMMa61c
L+YoNi85s94VZdSXTyQJnSYfswTDIguhCskF2R/FHCcIB2ZeqKIHk+uboeXy8PeVcwZGXYeUVD9U
5qKC9SHSC17HVol9YaFhg6bercHV8yOcm1RXlWYiZBxm5nAhO91kHuNB/Pfkgdle/+tRv3oAS8sf
NxAf9b5KwDyB/4fkOVOF71xcfa6fhm1jaEPhGomLOANob3rtTJYclb14rrfSyvRRn7Si+zYaLZzR
Rb+wiFY1awgFYNr1y7m+Q6FxokyszSNIrLBhRpeeibCxUx3qtnEortvhEClmrcroz1+zUpIByqka
iYhMg5tlKPn41xPnWZ8AWUaREgE/5k8NKnNhMYO5cHNfSOXUo5ITxf2jKUfXEdP0lf0eu2wKzHxS
zk++j+sOClnLCp6LsPPhkjKcMCe2LYyoQVDZUXN1JTwp3vSYk6Gs+WkJ/kodBHsF4wG7Gnc3ZX0y
PNdIoPZ9ZtrsKOOrbXeowisGZGsCZE3zce3u7musO9U6aCuPGvkgM42hvjVbAeIHbUWEgzljnJ67
QFJPqpC16+FjF/NaOja77OoPK+AwJKpBKRaUscZqpcKKiO8g6/F4j8VxfNCfr8dbJ0CjltKrDAro
vUoqqbDVd1zTXhbcvpxz8u8euKGmSacgl8F2KyXnjSPNvhZgw1Lhjaa2hter4ApYv9eFmK+wRpRZ
G8tArcU0SCZFnphUbGIMzBYjt63YRLJ3CnuEVCxJHs2pe/kP/2+JoTv/FBWiQS4auktIBezNalPp
jb3mD/061zraQoIIaah60+RH7WGCWT7CpV9ETk0+SkK25LKWARhqiAhp9VuqA6/mNeNQoWnEYzmh
a0P1XQgsdVIfgIrwpdWQkG3WybTPDaw19yfuVTnwk8AHajNsW27JbPnJn7mx3WsQ5jtYRUYW959A
GUrE7lY6TomQ8N0SFYabNsITFnYBW6+wYD6YjjEoB59rv3Ef9vLuuX2DDWnUJTbM6QpNv1YCov3a
KiPj8TmJVWhZlBNjjHjSIVQTa7CrKnkqoF/Tv6wiVkL7rZOHDZ6XBQ8q3cxg1Lz6QhehrnD89UCy
TKsEgbBDPyzuGltac2O4yd0OsuHl05IKeqvUGo+yQTiGzQyFthlAq2J+BdveJdIfqVTcQCb+dLUA
s3mzVkwQpUF6OXeBehRJNv1HTWXFniSVeX1NZkoiI8IkH4XaupPFhffwvPcOBeVYzk2f3HQXYjMZ
yPKADEBpnEJTflZLXU/NxhmjbgNAIO7U6NizQvdfXkudGmXPlIXs06OLvnSY02FqSVloNJG+TO6O
xueosJmwFxqMaiyxOAL8cGuYCxhyvQZ5wonMVLbmuEzTK2fulNozVdsaXfLd0977A2hxRucUiBqp
qYHK69n/72VuvNYUV4H1CELePpDp1uccuvUBP7b1zcF93FnF43zqjN98uBSb/iGHHFJNCaFPjDCb
/be/AubeURLWZaPQ6RjYAN4ozRCAukbL2mXT18ZW2StcxJYpxgOsN8SPnSCpil471huJxAIKtIQw
JJv4hJzzAFpnQwZDR1AbwY7CfELEof1IIM636TQBfPMW9mTYyc/652jX0l2ueEvf30Fqa7lhAsbS
kW24y6bmvKU38xj7WQqulShLuVyq0mhElT1g+FyTGEkTB7fD6li92kJGhWYfsPcoe7jRkTGEL96v
TqrlM+TDL0xUGkfrpGZ4LDlZFMrM3ZpGnxk0y4iIFyblq0zi1nap7U2zjKeTNUrDf683RHQBgOCR
6C5cYyLWzDPN7NhgpjeltiUi9SSRxVgZVZaT16NMV1SCtz+mkGriuYmt5Q5Px6T1hfijj7OzfYSb
wT1zqI6sEF1MCaVKJVcwqzAhbCTWmzIgqB13wzIJ0aqCoVls3BKNE4VdT7lQTvy+R9BiFvpOZHEC
EjmfbhJ4mf76UgQDgxGAh/7j877/D80Q7Yf0MTY0TBGfd5aVpnweor4bXKySOnYTwCXAfHvEo/ls
DesJlzoyHlWJe//R4soU8oG/kVvWpOh28sVKgsdGimNgypfmJsC7aP8MO3sQoajhr3ri5T0NL3UG
sCLJOd/M9BVZdDq4S/hdIeZht2jgIkIVQDHb7XroARYtR0RTAUkW62ycyXyrLVrEyKqPeJB6HjGM
KX1wCEGRIcVYzwNvM+TbE2zvWx4Q+pQ4+8bEnCH+xF9x+vHIOEDwCtQNnltn4uNwvxQ2mOBOep8b
4S6it52FwwTIw9VrL/S0ZYYpnkpzHLi8VVLu7/fsKcQFxscOdQAA4qnYCErn8KZVCloNyGdXDVWA
wudlI2pFDbJ35dFn200uHs5oyESut38LRk6O2LvycocNuizWencgz2Lz932Vm1Kh4RY0OydL61BR
nzj/kN55QRF0IUd9MoZW0bJmy++6om5QNh1qRYD8xNEw7ANsZ01p+Gh5nu2U726nJs7y2T9CrzSE
vMOkaZ/JwWsr6Z0VumpPWJxqXYZ6TShbOOhKEqpFtkudhwJKvnwR71egPeqaXKPg4CmWDLCe/4yz
Rs4ga4a/19pP3CcnXB6/IP/6kb9reoRoFVOcXqrcnsBdWw80XomuJ+0msL9xdtml1rSSFI0zfQWh
J63bG7EDj5VmFBP7IujR13pY9y3N3wuiBW3CNTa1IAs6gtPvdvmSdm2tunCh9sBpIhsmR8c2eI1b
bPABy5HF6Tbe6bphy2Czgxn9hNBH0EAro73dtVu3cw8KNmeWxq4WANqNRuVa6geVxId8q7wQDe+e
eq5g5HkGVDnEJL5FALl9AfxQoG2EQlzvZK5T8Ko2TIOBtpFVgkg4lyidgsO8eaOGg0w+c3H0yzCP
aaX2iDIqrQFGJVOGGlp23z1KF3EXb8MhvtCizefNoGgzqrG1EPvRMpkFZvT0awQIhcEzCiN8r1fs
7N7kuSidBqyQIEXTBtCqf8BzfnDdJyy6jB/9b16ykS2TAlK1ON1gu5JOqwRxwWPlVFqijhELCP+G
oqlZkyKhgryyXlv/2Op+x+ZdvRl14CMYWjqS9hBOYIFFowLo8uC5Ln9zn/BwwLsGa0vNUUEJSUtr
OElJhbuHiO0iiHVPA7UToQdo+6DXkyqV+hyci9XR9bbjAQr/v5SS2K6c2zpGi/NN8IK5o9uZTLub
4eRwKizYDi7Hq542gV0DJio8NPuWE2z1S3glexI4WQ/F7s+ZPw3XanPQBxBrQSZ83iSwRjKujurk
1VQUUnl7M3VTQGdC3i6X/JETKPMkXiuBcfRaPVnyZh04Xu7FHEu7j+KXTMf13nImZNjdDPehWrxJ
OuhybbZ5oWXO2qT1PK/G6/jFyhG+qzInGfvfYCh1zWKikuJl2hdZtC1DWO6YGI/c0W7zJDftM94v
E5oloZVJInSizBxjxqKjTF7scT49BpkJhFG7knb7Oqx+0noBlrzSigtiNsoVB4jkzuDcJ9JrGyNR
OgHPtwEFCGNlv/KuNzIAA0jxJImlOeh4MOQY7uyhvQ/wQ0SjLmGX7afoWRJyONkb0jTpW6XrZ6BS
vQbUC+9oqfqp+hr/wS1/BIWVw1a6qsLPk7riRAFqIIAItWPpp+Cnq3qMs1PFPk/TjqXVoy5fZyaS
91FiwyfrH55cXOd4fEuB4yLG/pBUYZx3lioT8yiwhvNDtZBOo4XkWlGvPurfatqDhTurgcrgsGXy
QvvxDsP4SX7/5M/WhR0BP+kkI0fV9NkXAijULbomOErsO3ftbxSFZOuffGJg6x1eXpds+3zvyMBt
xahozRrDvR1iZIMcWxsJlHx4FuFDMyxcAq+ck4PnXLLjL8fb8ti/oRvLOJQ1JNjGgB9EnsCDoQKa
uxECHQNlIGXtIBR3NoKO3s9lnpTmGdwTfpdxCe6DHq56KBfKpv6Lwo3TA/ovtWnZAhDDqYJ+2pH1
DlZXcIKqYKdj6LfISRLbA9RXjDs9eHn2KIz/zzWJ3D+NwfBlhc49vYx14tLf+Lj2TqiMQTh0xHrL
FuL3680QQsuLHi/bslShD+Ev6HDuNUY4X+XdCfYCwZWuQxMSmFx57PiYB2C3d4dzEGccuZ+RbFsp
ShqFdt7amUgKtAlsvLl1wSNjs5RdKbQrmTOTqG1PE1gyXSE/4NBp+CPgbl6Lh62yUeJjccdK4NIs
PEG5qPn1334vpbc1E/yEuTvheHRRplH2sUnEfkHkFL1pS1pRRF/cJyNMVk3XWmP19se4i0Cy7pDh
mHz7C7DN8KOORwLVR+4UVVIIg46pJ9J55HA87SYOgpS9oXhLTMjSHx5kRr3fG4iWzgPmfrGDGStj
wP07HCPJ0G/6vdzfU2/qzBUM/Kus9xve6LZs4s9ZdHDo91mBjOZX8lcGXJ2F0Q2wIV9mFHAcxYEb
jEgG1rJCvkOUpkjBQ9DY6bXwM98j13e28rKDW5oCBPBjyFbeEUs/KXbIHfYN7mBK4aOZDfrSxJCH
lUxbrZi/Lb+YYzs50y69t0jAEb40YUq/l/dLuBr0b5GbVNfsHRpATzes4LGawO0A81Ne/szdZ3KJ
C/U9/Sy9TP0+rF/0LKltpVjvmuqTbCnu5QhITAIfuyba/bgzpEh2n3QGOx9xIe5oxt9YbEOXrFzj
1uwpfKNpnlmKHywTqMERwNcUYu/hBr7ePl5QJ7DXpsKZEbpxCN7Grh7cZGk5CtaPb4oqaa229NSk
tkRWvxj/5qSA4q2NtwWA46fWdVXQOMyCQU9R4lvhZOAvxJKWfGYw96Ht0kFKhEdnq9KjIfehqKPg
so3fm+j8teAgPy14+ZBc6ZFjvCB5YB//6TiRmEJi04Xzf66F315G3X5z0tkqDUjcCTd/dTHAF/wl
872t7ivizfykcZa+gvhfRlQiVIQeED5YAMBAWMYQtvgH/5lqnu0aKSH2uWJSjnRjf+aGXzzBNo5f
oPNabOdMqD6+ZWPQhBdBINdPraGqpl8Vx2zI+D/EGDaq0+3y3q8GdxT/1Itu8/snm3+6yRY9IPuO
fev1PQ71r+yBjs1FTP/lf6Ld5oP7vvo6XKygtjLH3Tr9vVh9jwJp94plhK683goN786+ZtZAj+CJ
WMbh5WN/ybOEe61umtpLxqGFcXJxJBAcN+i6aaGbukV5pqSW2oIar4hKYTyJrMkSIW/EcKt4JJ3f
3wVwLNUvmu3FP+MRnbG9mNZtdF1CK5G4VyLDZCGYX73cRpRPox75y/RvsyO63GrwucnaUvx45qaE
8X9l6B4Ike5JYJAc36SkfC6Qe609WgeHbV4cKALZwHD3i2+K9/RMLxWZE7s2RzNKaNxgunEXWk5H
AoaKUK7ipIy0wE8sjXZZeKQseokoOvrX82GarbD9zL4NJfMUTj5VFXoojcr+qn/+AtykPla1fbTK
Oea56OWiFYbJxe2i1SQCGBljserxQSitORJ2fF9zOxcboyG0zXH+YcKUtbEKSi6xDW7ly/rmRhE1
APLPn4rQ1Po6Q34QyOUJWdRRFSmzgq9lpBOQBxcCDbCuSnvPJOr2HMVgj0T24M6ZPPAVVaq4HSO8
WttdX/VBso3/0pFFrI+JS2ETkhYJQeHHonMZNLv4joLlPFi7VbH0RQofmuDSOL0mqyOqgxIVt+cr
EsaVpWGtc6c88IxH4s3q5rWYWQxukgJD5yu0HlzcFmeqDAP/43cYxp6TbL//88XNx92ZND+88HQa
P2EUL8M0pyR/4Ki0kQx1NEHbYaLqlibgZRTacyc1E22LpET3F0GtetZG/SGW+BmpfwWT+smqJ0ZU
id9fljEp3ZCQed0GWFKWqq3VQ3kfCHVuSyPDZOYgU5YmuC4ejxDOry5/cWO70i0JZfPb7afTSlej
lIELV9MnYVx3Rr5jhdDSDA/YksTx6TbwQRwQJaTonQjbdxWTAb4g7//eldSo+Zy1gHZVna3O/W+g
K2dl15IsKuJYgSD+xxrylU7Can+7t/VjjOl8J5l13XbcXUSCQWVuK16EAfChHu48X8aSJT+9XG6D
v4bWu/e+t5CIXz526E2scEnTd7apvU/toUoWTD5JCH+NZDRDEme8Yj5msZHFb9s8sOz5m4UmW8ty
BLQBiWvAgs9amcnHOqMzdEFW0DBUeL0pXuqYjbOYx2rxXhl5O11r3NEi4KLpseKVjgebiHXB1Ajx
7Bohh8V4FbYP/cVcipf7K2KmtmFA87DGHWrMpimWXAljYlcXeS3OzshH3ZgBiNHbJH/yw7/g/712
0f8qzINMm/9F3hYNDeHotj7FeJjJcESCkBSGcJL38paVmNLTOSvV7vNhiiC9J6KczdA73rB9pSD/
T+DoVZ1A9YTIBohMppAJWGl8fkcEgTNsFEsNK5P/t21JcbsjAzoo5KCzXRplVQnZI10eA3yGKOEO
3jCbIbVEaiW8RV8jQU5e2cvlH0NLZ0Mu9/+4zVDejm2g1A8RAMeIUOLlqP894IKCimvkS+fDHWlU
eP0h2s3RnLUk3vIdUUDRi1UVhrqb9+SvzOkHrUySIwK2yd43HwhhjEhCtMww83rjnLE4VrBI8czy
HJRd6WCebacT7kmTZu07z6Yz8PSsO49vqDQ4kq2ttD/h9NhhU1mvyBe4r0W5GXwpgCI6VnlmDc1a
D/NS3LhY8oKMt8rOX79I62ao6PMrOuxV/FCnHwLr+6IfXQG8G3PEFv8lJaIN9GFXkMN1OQF6Jg6b
tVeUOP/S9H1x+U9YoV0ldFs75Kig7ooC40pavSBQgYHIW08D2gQfd3LCsjILLhFq9TPTXa6md1Xv
UurdDtY9uGkYxgeM/WdUdf3eoJakgTQEkc8sx0sPSok/mTgABlD6/ygtJUdel/WDA2CjZxEkEuc/
uj1DP0WvLBEQbyVqeq1W/Rjns379NKRUBFAJUdx3OZoExfIjJ5t3tgdHkjcIGN2BypxuNQoMkxvw
9sxyugpVxENjoIUL9aTkV5WkOGJ3RqcFiOqDxEYRckXeCfFLxX+kPZFZmTiKKhi1ccPo3a2lKctP
4p2bFL8s9L/szYeKoYK4aDJBtdFk05gGOxlUCI5hiwRDC+SVvqdR+4qEg1MyDQhdLx/Gmoqcy55w
oqWdEtUqs8ioBLJHz80aNSqpf3fH6KPVCb1HH8XNs33BUUTgARScjIxvcnMIPHvOFCq1F3S5w0C1
QanSRtbgfD5bgpl3TQxwZjfYEzTA9blV4kBYST8S0mQwISQZxFhVxhtserOMbZoBnMIoxOnkHXrS
WdfenSh4xThCfFEkoYnxXB+TNfAiG6i3W5Ff70yaajiCnzK0huHSLEKz6C1PK2UHfpp3RJkRTb9B
JjLwt4+2ljJVKIyuma/zyDGD39A/BPVYW2TzPKR3L0DSscUNa1cet5oF5mHAW7s4QpPZzpI6oyvX
rnJMISdxAXV3J9mY71n8etMLbX/VQiaVqApjh4JoCbE3fYFMP7JXpf5xws72kj1rIg21z5kFv+K7
icKwCrLyxWrIjdff8FlnuP+XdhKG3YjHgpjDe48iqUbmGhOn0Uy0ViBCNAZRIAB0e/wO4ssJdVh8
KH3kDpEbY64dOA+Mg8D6mAguQ/8YQbifaHKP1VcyuyUCN62pkBAz52RqzdgMrS5M4lvPQj3uhNXi
NFylZWrTYEnUH7pwLyTd1uTCqPKSaI+DBvUvOyTDZ0weYbpQ6419dSXznG3xNT2DoVDzE09lDP1M
+hIit2m+e8QVh47UtuxSy7fmaIz/EzUizuAEZgpdeGwF2DD+LcWgJfpxjh12s41DoM/k+K76KvIR
NgGCIQ60Esyoqdn6yzbLiNcPmx8Z6PW8e+AhZvkASIWXhrs1/TB1BSZC+yWMgy0FF0oozftyh6c+
x9gS8Hm8HXjJNb9f2qtXaO3UGmBg0nZ594GhbTaTl8WxWgzLej3SDYBmlavrSKD13oOf0DKWfjVI
7W7Ykwx/HhsageR4iZj5Yjvs03k5kYyCDYFpowYsc7+qIW5N0ToJBWy/5G31f9gZjMqH0gnRE8mp
idlsXAZrWER+M45DF9rfu9ZhOCyqdutUG+BhnY6q/WTA7ORJmM0EucZ17TEwZjDR1Fb5qkdUuWYI
A4ZL6lm+34E5sAo9RZyXK6wrU3pdDaC0esN05jWe3IkgnYXdNHudwb8fFP8GENLDWPj2cI6CIabA
QiigF03Z8tpRrfIEv3Sjj1rddP3yk6gMjgzeFQIotiq3SjN7PFB1/3gK8fLwkDcQhPN6kHch/Pyw
ZpN+YiWJOrQPzDn+7kz8kA0It2ebSC+fOpaY9JRN4OKo47Ku/JWzkvWguIYSiICDY5LPo0qwvmuY
Z+78ccZsJrB0d1DCzZSZ9+Q2fqq++a38lw3FZ0yR2KStYFEMxxFj30Gxi7QSBVtrX/zmbZ8LN862
pzjQXGUOGkE01WQFA4nRwKRD34fvxqM0qjoOjnQCJQV5uZrW/Uf1HAtD6yf0x/ZJFT5WZ/Nnpm9f
THEe/kS/oVrP1i5hyCfcI/kq/x/buhft3EdRfZCSmGTShD8LKKCuAugSJ+S37N1QCZWVBKQm0V3y
mITYo3zdvjbuYSbdB/BYDXE29m0oPKCnCKCOrCfF0SCpwyOdOwL1PGM6BZNTS0RPPdlwVqXvryWu
+gRtELSIXknxixsABlL56BwQ6Xk394Bysx9BaO04QL8ixz6jI2A35v/EytkW7hNb2QPb6k2/qRnR
mm76B8eW4kuOrmWwrG8zU7UdLSCU+AMYo6KCrSQbs52l+OcundOqvS/mSPtsoPk/k81NshIyIM6u
FMOij2I/VE1Rmr5XUJJJjVnR8L7N2+zakD9SI7Q7J3QoaYWXfXURPn1kDDurA0+O9S1d+pTWSlm9
djYRPlHoGRW+yhzgj/uwsLGtu6XrZmvgLP4peUvs98Bj5xs+2Jeo6/RymG+p+tz+pIljgp3fc1ap
/zX5Sn29UEsPa2hznYiGUSvXOjXbd0GyTs0iTS1+oF3hf3gMUsOoLB2NqGi7upkWik6lfGpuoQMm
UgQe7EHG4/sa+bTySCcmoXB7VeHrwy4UqHsRNtVZEM/bh6IkKTJJ8cH+Eqh6k4MF1z+5Rsl3K6j+
ohV2hYVKE9iHOx89ZdEhpbyi5C3juKoAIG5Oxbf/7um/F4wiOKKojopzCiF5hB2ueeaPtxJLUwGV
idsF56GqIuLb+pXFiQ5IeQMCCjRcc0pEHqXs964fu2sVSGnUuJBt05cunfhzfxhbdt88fCNDSIRc
9asdQOQf3lAZoSbfpPV4Eqko4r9w6LEA1OehitXbrkSqRityv2hYqPzPhbMd9xYy6g6SKsLuymc8
e2EWS+Q8W4SxnJejDFqKPNG5vsLwZputGCBmp2Ed+fgnZEd1IHYVy1fT4P99laaF/2sHOvFORxjj
McDBpXolbermT4QbPBVxb3H/8ZELth84/yzx/PvDM14ME1m73E47TC4IeqEVl245Gt6ZX46csfwc
rZU3XdNe5iRnvgeopjlgfW63C97nHmeMhco1cInMbkGfQo4CA/r/Q0AaPo5QqTnLybRNYtOpyBH2
OLP7RWIEvLsYmcZbd8Xqge7136ZBISeuBchbPSI3kw+ECnRcpSDexupUv6bO2eX9IpRVzFuhdl/U
d+xR5BNfrf8qR9BEXdetSOgBp6FW/Ah+A3ocaucIX1b6Iu5yxcs3Xsp36mIBfVPmPI1mxXYYLfaU
99lpFKR3JfihAldPzF3n+XQkwX7NZBUv0lJFGl/94yo22Nqe77ojSoqmTeS8RPSW2j7Ek+Yjk+sE
HKB5xOG6NfhnOHKD67ZKo0me93gcX1saQU2JQhwvNs+GumFvXAnORLWOGxcviW8HrTYVV3I7GDD/
D/lg7asHXXJTBJ+ccjq6ixFpEEXYb/lzSg/MsxJrjmr/p38fw8QLwPYxLTYKlTMxo+MkIWgGLQIv
lyAyX4NldTtp3/yJhDU5t//X/usJBrsLzCV3+DvT41O6hUPj8yAivNGZyDeq+mkP96lYrgkyuSMf
lSt7Bj6ImwhPKiOxzUWYyIEzbZSAC6dYM9DL/6xc5xYokvWDEqls8CL30/uWbj5Elgo2KlbydydC
/PSazaTBq3p7BCdSlDsafbhzfNEH0aEuJL2zCdr5xPozxjeaNbs/3Z0WJ9qWs+56lsfWCApmKrpD
MyxK66VPVB/hS1KOJaz4YymGtCoOtOUR6uyvgAUI9JuMxqgX1RXI48OvFtQM/17TT2u1kyA5EQt5
tpeJGN2A+0Q1NK87+L98l8UeNyMztd4o1t7JbvFQL4m53CGrmF39WW8obAULukUVS+ALVMmHAsCq
C7oobf6Xw089ubzKSBOlKGAT4jw4wsboRptjLnVqxEViBW7R3tgCtXbfaS9ToWGg3Tn5/z6pXAUA
MMb+Uns/DWAbgCFi5xnph2DyeWWsbhOzjcIo7mgVzB5EcwrR/4IU+QD1LeVgGJl3+TztHvSgW/Sq
CEMoHX1LHLZ5pvVK6nZm3VFIPMg/jvpplysmr8aJe/a5FobYVpQagDgSdj64J7VEzc8cqpinOfyj
3eFBJbXgyfD9tCRZ5DTBbz63nLaueruElgC0jL375yo2BsnKaiTvhEC5aXSc0a/rCNmosc18Emiv
j47rRkJBhbEKODHukAGu2T1/zZT9HV5vcgSkz3rdxqj8vVcKLpbn2F9zFoEQQYVcYEsv2MDOx2/M
wrqjx7nZI2f2NOgLRB4/2vYN9yzmjBHdzbAV+d6e0NlovUtzZA57rBRV5RLFSqmkudH1kckW1rp1
g/DRUYSMkmc/uqw3As3HAkW9NJdxXYzDIrMm1GtI3TetAnMU3Ls145eymLuWHbz5yxVu4ReD21NF
QFDr8XHGbZONNdWWIrzmZ/jnjUpds+/2F9DqglPNUt4VjoZCGl19qGTqkjuEWRQun77ASdlMOJ3h
kFiXxZg87srSYj6wX/jo4tBkEGtBXt7qamZjZFsKoh4l/jT1bBJdE+JfJnE/WW1uqS+wi/LG/DQI
/jxneeuH47wWStRVJZUgDS13tkV6o8uK9L1pd+ZIy7+pOaUIcJLkQFQhVl8SfGioYO2jWNEDrWQz
XojL1ZiziG4gxlWa0jyDPSDWTz5D09UWHzk4nmQ0B+aX0S5r4EtQFqTFWWzt8PFUAiV2dOV4+VXu
0i+w9OyZZa2lFR/GaRfDava/lOo8tdCU1mJV17E0VGZjFIpNG6UDM0NbiFH2YAaMk2bpB/rYQktv
TfEZtbji7aqhrLV+XIjSK8nAa7nUvG6wRcR9fGeNLfbUKBzvzpj1ik6GiDW780iX3aSeTj8mclXT
C+lSM4chclbXDwfZs3Twp2YRKupKIR3wo//ZjOq+zhuOJHFTkc39BmFY1Fvdyi/YsvQbIPlaYtwr
8uzgXGC+NYUe9xBknH+yHMjGCzr2R68YqzrnJUBftd9nnzkPmHSQBNaZLpdDOqpyWNf8hav0ElDw
b5uPQfqxA/tABLWOVAi4/Pppt1xO7nCVoNcGljSqAdUH003M3m69PlNKrHiUIg56QBDG8BNFgNAP
bLsjyR4QoWeAPKTGqq0wQ31+v61jVBRXDCLrIKSWJ8WUsarleFkejXRyYYcoimG7PWmqku4+8dCX
m13QsPluPaZrlfgMLumHKSxMgNUmW+OsgWgGQKaRv/oFA4p4KdW4kct/IyR4O7OVBoSLyuZph0xn
rMgWTzxfikMzmf4BQH+gg7qmE0hmdmoUFgKljORGsbGudJoIPj5cENyjnRDOV7SsoI0PYuE/JfQh
9rLCkRSeED1Hu8zqE8i76M2TdT5ky+khFwpkgIR9Y9pkoy4GxrmAan/X9W/thK9NgKCiNdEWRp7v
PWE7YAq9NOFESwAKQtby1UU4EmR9amM9mPM1dGvjdIsp+Z5Oio5rrO2tcPpOc76kQXlBkT/Vrh2O
hCTHOtz9jBPmSvHJMufbqqvCG/sS6AaeXEgDLJbDMgFU42k0gUTjnPektr35moIbx3Qhu+2N4Y1H
4m2oF/VhxdOCIQ3BgdvgSSmzBj5+UPglDwdQRFDmp/cKmMi5X/frTOUtu0gbZjtcRZnvGnW9G//R
5b+idzfni4DbWAIohC3gimIN7Fseanc41X2ThziFNRZMneFoycyxiunu1ulxxNYLQWSi/+3b2ck1
/CYdMcYBnLkZD6/EJ5NH+67VYpGg4KtcBho8gsLQputfbMu5+wv7os12bNk1C4Avo09+kJYcWH5I
OvCNDK49qvNpj/N1hp8fllhcj5zSLq16Pey5RYwMf2Ywp8RK13ja+DDq9SG2nyB7wru/0y+Jk4WH
MVGA4RGdmtT3dF6e2u3+RqtF4J9ezpgHDjuQxsd75Z5taK301wYFY0NTD1lnIU/DcpmivGlK7beb
dTVedkM8A4cEKIDQ5TKuIb8viOeoENGDXpElI873VRN2Srw0NC+HW98Nd/MpFTh0x0w1DP08cwAs
92GMWK4yCFM/36tnwnsAhAZdrlABmB6m+hbdzE7sCJ2VXwZtMPgs7BdB00oOycEyA3zuR7Q2PSFn
9bQ/biGLrbV0Z//fO+HAViDj1Ai8FjfnAzQQZVFD/8Y60ojNR3J262oB0o9GoR5X/xHmjRjy68o6
wVT51yF/KFco90rvZmfxS2E7G86uBKeMpdW6z8tpCTPH3lg9HKxx9VVMMkZGGHNqq9ahweukJmSx
i9CGTv5VzC2awU88cjedjpXUItF6JhOsdQuatYNcew2vgPZv+w5EI/P8nTtK9S5u372IWJBHNrrU
Ai2J8FsGwVUKsv9DrOE04xCU9z1SbGKdP91fsMzKXKn3i6rZvFhCyUJ0/1ERma7Y0R/w9rxms94z
AAd/rafGFTQBVxsltSFJFhEw2UTn3G7OTdOK5BeIfQ1or3huBFafv5LZD1+b5qgT4dLAgVG5jLOp
DhQVmXYXdTGzG/P7xq8eNjC3UVUXsxWqdjF8aRWuL07pjgXB8D+Wuym9WCo4DjjvUJ67qqAr+Sbj
NxWaFkJV8fHf5Ce1eUfNAvWOi7SSueRjF2COHsBGMoUJ/qm0ssxhpGAB6UpcqA+JRttJ2qSffRob
1vVZxCeFwOZIlJU4qMtvD0NLkfFN23KEM1/xfqsLcJi4TaZRvbnEl61A5rjmw9rCX7jbQIaHdwad
xrT2OUBaHA3yvb6Eqti+2113JN3hK+0N+ePRC4dEHhMPLUW2tFw722KJe2F45CJoae57xz3n2lxz
pqzhyMmkXywyq46bjaCTKV8XV3xkXvcbhJOaQH3GGKKudUubdaS/bc0XO4CxT+t7TtISpoLkFHSV
5vlmavZOjXysyEGeYyc9yUy5++c6zM0nrD4hu0wQSLYQIXGM/D5Mc34434gOzAyFUh6F8igHNvMs
Vx2l/5FV7K/h3sv/Oc3u11qVCl/GSvkmUFLPX8tbFlpL2NYrIcDfyc/AORaJeTpnQdB3S73/gCdL
peoJphw+WrbtY3Edd5Ky0MeGQwm5vjN8qeGsFiqguSPavXGxjmuBzcvIEZgM2fhAOqEnxBxUssvR
O1fmuXErZagO1E+hwDvgXwJrSgYJBKDjwRyifz3e9A88d8Gh/KenemIMynFdomYJO5JWmXk5HKSU
jJqgKlcAib6aeORqj7oUck2mF/g+EHLcl5kk+P6HJHV0MtGlAGDfbO2UwoA7GT+guscZM8/6d92s
kqlRNqJvKgPmvnoFhgWVULb02e2S7ftMQoWaIXzP9hOgi67eCIdl9CB9qp2pny7ktPKK9KVRwpnJ
EbPKz9HG1LXFiMyKnh4dnfh1AhH8iEICrEhgeOtOuVYmMUj89QRujfDFRkoZ1als2fKFitdUZ3hm
8ZY302Eil7nFSNIqTPvkyIhTcLutTxUnor7jcJsfsOkwmhwgcOIntKTPS3gRsKwHugCAS+PT30Da
3hD4Y0n1SVRQ1ibH1JXFTlqwB5rFeV0Gs4yLIlieSA3yayiVLlL/UKKnyZXETZYxx0wDK+5KkFFz
QP5F5MBPHquUm5nRP17gaxsPgym9P3VS6ANf8X7bn9HQyT96cSJisYWgUwlWX3NwMXCnMp5mxnK4
zLW13ZJsrdFravl3bAGtXmS0nZHDEGG5mwrLEKBkvLYi17WPRP7QSoZkQ7Q2bpayIHvhyWPkeaB0
Lk3Q1SSNnRbWN2NiF/ieSRR/mlxx3JXvWf43x11zfvou8knwpswweu8WzX+ePWR5h7cWhytw0Qin
NUvl+gCpVMthhQPI4jOXFeTyOX/QeFG1mgLkOBRdLTrzwWakBMjedVTTJzfA9f3kVJSw2aAFbJ0p
kEzs5n/SwDT9FcoQFGpmn7oR2q/cQBCCsADrJ5e3fnmgcgyBeTQQiBKP+lKAz1sl2zICF8QdxG03
UrIJA/WW31TiNyrBd+4AnU/JXggs/FNQgDYJp5mNu4EaptH1YQB/P9//0D5zAufORlV20urCSqoP
Gh1X+2pdQ1A7uHQdxOUhtw626bBAF1InwhY3OoW/7CMYDDoUd9/bDLbtCBR1rP+RGz8avdoxzBbY
oU3BHwJ1aqhVOuzHIh8oYgRef2U+cSSu0pdJ+L2JQGMRacCbJtn2cRtDoAk18Io4ZOwdXZtc4Jhc
WEB+8wKVlazPCB0WhbSbcC0SaDoDaxdJxI/P7VY7+oojMdJ7ILNYjyhtf+jcnXG/4L+hKBq1C9+r
PjgCqbYaLJL0IhYAoRvjuIBelVwJl+D4XtzOb3TuRhbopmDODJ/sjd/n6Np8eeCdiczIf90jjV2r
qk1OQy7L7HrTJ0Wjex2YhQi7QXPnpBv7rjfuydv/YV1VvNCx16WMBLu34X7JZyTnl0a+d4cw0Nb4
nkY2rMs7BuvrwisKxe0y9kBfQUgv4iXgPZnTOeRb8NNJ+ruVZHVfuFoWJDEEq5uUq9rFD2HJOQYE
Gka0EnethtC2TkJ8ls2PSNBa0ughB+B+dLxxa8HxfotpCnOhgnv/ovXOhRVZFUAvEvt3IEiTVpUD
weQzVw1fBTI+G54DZg1iSN+nJiqgvWwknSlVI4ndtzX5puCoo5E66lf9t8C6brV2AXsDrUHESXCA
HkaPr+tEtstoIzEIusQz+o+fSeWyA/Nm9vxT9HJ0/BS5eaNpVn+e4nCelztF0vwOdgM7iN7R7HOT
rXrogAg97zRmu08PY7cqtZYkKmgn9UGDiInpau96asLcFVHD0poQhtA8BrvTZyUtHmKEfqq6Ns+/
NbIZu3smhV5rI1+O++UvMBs2AV8YFhiuQDkU+xKlyiYbAlnTk1xkDJBq+yJgV1MTyU7/7wkxcFg+
XEFE1IW2+yfmA6A0WZyi1KVZscuUyWPqnRLQnxnvnUUj9fk+T29uhk3bpxnaSfWTUcOmyRhrL/F5
eNpf5DxiwAyOJHsOiPZ43FzTId+858y6SSBejAOg5xcC//bEoU8iazWHCxWc3TFtcnNXDmkzQQyi
OHsGcDBI9EeAshnbjC3ROLjcYHGhC9Zqc7q+hbVa2nnzhOEOjRQ+1xtnpydSDi3DXjcsuLk+sO1u
gQstEYconM2jfMvFuP4Tv3I7COYAQB0GGQLSzxpkJgusJ5cB3hj8Wx9Q6Vgumc0k6bZ6UIHR5q5U
DHw+Ixt+LneV+QOaWYs7O2YIMejhfyrdtk7S0lQEezduP52M76o1M66hhg+2CT7kpEC+JPwD+I70
jc5g9VsgK8Wr0N6rMSgUD2EdE7d3RCafXGwAChbK12otnXRgpjCHVjtZBcEttihspOVyXI6WxDnU
dY1F+3hSJMVjueeWnXtw0+LFAd5LsJlxRAqTz9QwjLzIUA4KtMSG0oBVtAehwSGi+2+InXZXbvwS
HpAOHhxwbL5jGokyO1G43iTxhm7PlyCtkpT1TH9UpTv4cyJRgUFqsdfT/iuz0e5nlAUGmMkZCW6p
l3PTciL81u6au/LPgDSOhUJY1pWrQYWnITw9d6Um/4l7lKUkI18NOUOxc/FdmTUp0woZ7wtOC45W
QcEsFVuJNN5GQ/RYjt+yep6NIrvAxrWyfdiuT1Ed2KzzGh4wOzXWSl65baT612jbI8FBXC2cMPz1
7KeVoFUQZ9ZdrC+5XPfr2vpL+qJYeznc4QAEqZOF3PTnxbWMKXkOfyVy35qpy7GIZ0BygGILsFNm
hIjEKMj4V460aSWj8BPop2UteCJZWCenj7rJkXqXRxUhgmhKAxECbebeKsloPO78fnkH32HS9GQ5
8ZYx/KunWaich4dGJuEtchz2eTvhTdtEWNQz4OwPjEdsESzH9alFGIiQF+JOxDzAisIgOx7hB7XE
q+zGdAQfRiIcU0LCfQpD6RhE9qA6QPbzIw6V5EJP/n5rhBUR+AfO1tBN0s3Rs8Pl/6bwIHvFp1x0
nKDCKqo1u+VdE9VmdJWeBtbjSzKbXfWtsFliBm4q0JQU50HHJt7EFqvUFZxQrH1mDTLpBCL1wa03
Bu4hZH3kUytU6+uz0XMCeQsAVXjpMxxymW5DJNU89HGKVh4EKi7spLg5R9D/UGKfsQzOhm+1ktKy
0Zu3cwz5hxJQH583+0w7jle9tirN/oeRGQ9HcYwBrPSwSqZkmKeR5i/X9bSW2e69CbWuocF8jiy+
5CDlaSOB6KmRz+dFCABRpoxCl59wjQZwLUpkOxioVL5vF2BVMOew9IW9xdxRc4tPmxig7LtvBMvY
uwTiuVnFkpJvkLlMU2ERMIPCXlo2mu/ve5leAS1c2DuIkqeDmDNRHC+qHAfajc5A39f7tRjZHzCC
UHJIzt6Kp3knv9ZaP/tnvj9SpLboGftfEoropEFVLGtEGByZtj/zQzRScmX5T1u+7Hnc284v+oQN
3M1qYn5iaufoA9f3UdB+xFFIxKomNpvshUWHEbm65DGaumP8PeKJ1F8kaKXnkwYGTG0u4BuYKmSn
WIaJbnXtcp/PdqBCWXOhEs9Ozh9K2TrYx9/2m3YpUL0FeeJBFzElVTYVy16T6qLrwuN1vbIV5PLA
fmWlqYDiOpgkT34x0EuPe/SrfIELdoSOSFLeXKqaqKbbbmcX08vLICpPOvdieDjJTV8mEggHa7CR
X7AgPtBr2mrKFDf96rNBRIuybFqyXZE+Pj8zVP1dJSx9X34SsEVDlYVcuuVnVxUNpZPJbxFSt0Yg
i50Xdxr7cKBu1bD0Vi8Z8sZFxI57H4w8bvFnhM5pmkAIQTIFjZXW2rfs+ixQMrmxvVftOk9Iv/Sk
hHwQvI7kUPzXVfa4clDJNOtcJQvbJ8UXop4TASFWD+qv5/qxFyVfKjzkGhkG5BUup5IRnoJK0HG7
wXDw3HiZOB46cmgSHFDOtGamyRnybj2G1UMe5tyOTZQ6wCNNX7SHuFP7tycAxKyYMbFItj2M0CFd
GnS5WiA8prG30ZJFe5WD3K1OskwF1KfUVJ9mkdAsIla9/xwpDsEv63bqv0P1C+UbpxuKJXalN76G
uZ+iv4+rPMKbuJIjSjKR4u1nuqBOQJXWm/9virkFov8nBCydREgSy9lkA11TuJwmxwo2k0mum7ya
d3YeN6f+MVSRMxFXRrisgufWnGWU2sEStxKnKA2L39xR4d0sbRXwuc9lieKEreZqaGTulID/+QCL
CongoFJoPqa0yXKZ1MlrtYM1chZmN1lyXZj6GwmDNQq60MeTJ1KfAsQk1qwAOVzV81BQsWRD+6n5
99EcaN4/tqVV8YKc3a3vNycTP2zdkMSVdQPxLMlvnD0TZbjkgNa8II5/ryeCQOgN5y2du56QMqYu
8demlEe4DDtr8zfmrBs3dBbcNIgtlbc4PKwz3gQxapfjYZRymyH+Y6CNEsHWl8cTVYv0NcgtKJxo
l+oRQiMQDc8ZRwbv7bDmR/ZoNLe6MgkjNAzbVpMdQ6ZHQG8vP/C3mxSubcUC1hQRcEs6kZeZ0jC/
mdK7GTd18KumYIvB15RHxqCJFCxzSBLSHYzuUda3DUPwo1LZVk7x3Yc+5ZLTwzHTVYIKlgmLJsw0
xfE+ky7ud1fnMXDxgw3pDpoFic5nehXx0XPXz6Sy32cVQ03qVQrOZlO847UQnSmenbF+DoyyF3VR
scXfeDwSwGl1FmIxuIaMi300bc0W38P9NeMgyjKTjpye9zfJGgq9KtctsOSK2cGCQ4TCqiOWpjpZ
Usa0/7Z4JM/vnA36mbDOMY5WndWgjwxF3NanZQevlBgngFcUfkv6fnw8A+WNiDDDcKNn+4p0maUa
GwarhlRgCnlURjFXIyvcGdYqJEcGBOcR2qGEMwzYfMtR0dwC/4vsnv/ySicfFJVrf0Zk8uXPN2lc
zj05P6s+EaB70m7AeYhFEk42njObCXZvqefLwgO5lF+hWWYAB98AAmynM6vqw4MqNSY3DLEb6GLT
yE+GVxRRLVHduICvVbWCozcFHrK2sRON3E6Aqxh1hlfG8h7DiuL4SaN0ghS0K1EYTQDcLvFQwK6K
Q4QYnfBce7d9ZC9AZiXz3B1YE7l4Gat5VJzMhkTNED7fMTKf/e6O8DLg8ttdBdaZvV5QtRm+8yrB
GwQuMyJunPXlU5Xm4YpS8lxyO0xMC4Em+yF3AdrEIfsMAquhv3HTuCcQ9tHPqoii44oQgUrtb2rt
b/3DVBii295+NfhjzsydYcHY1yopfp5qnz7fbJnmIr+429rYutH2txlhBk4W8KzvlmnlRZ6To1jV
+niNWB/iwk5mFtbq7+mgTjWBZT+yWgirV6Ar5gcQpFzquvf/IQ9LbvQyVVrfDbZm4IXRX00F57dP
MJ8uovaYUViBbnxS5X/xsB7+CdgaRMGv0P+tNII4xTh1gTGzF1NOeTLmTSUrMrQka+ZH8nxGOqN5
u1KpQ6hlzmQBQCkwlyHLWwbiRAvhC7tj/HQ5UDSCRb5Dyj2Vh6Ku566FmRYnLPs/x34p2FSxpCuM
kES6krdOyZJt4IEEHigijPz4nj3aEaw0xRxCBf6JCGbDTZ5+WpAmLZy508CJlnQmHkPadeUBTQw9
gCZtgpmKVJHIYPpG9Gos22nQ7/3+NwVn+S+It4RT3McHdYEgDg9DPF3dcZW1B4aX87zCuPrFsLtz
G08cksFsoVX1MHa+gr8Wm0YrzjDiyhvX1xL9qqdokd9m+lwQN+hd2YivZccsArWJ8vs6yhl9ZedE
Wc181YJBL8ZKFV4afgBcoP+/PI4faloO+xnO4g7Sm3IW3Fwuxsx5IVcy692nEgSjBWTQTfAk2G/8
D/f8Nh1IYq9UBI5bzXmhQ/9CtICiqSYPf2V7/NmcrbcwUM5w3XbKy4DiJoKWBQPCcRrtTiUY8S6+
Iha38Hb1WGZBQXHW0+UCkHXVqLucWZgMzwTFWpg+vZce2pnnqo7OBWfBZDI3ZlFDSRdZRdxgTcWd
wcJCzQLlv/p34oxcSY/uUBZZw1LYOrF2kC7U8fI9uCqI6qvNUVWm1mSgoiimRzwhbOMjSwyp4n+c
S4+X0O166hRNgng+dGdOu7mhuViqIYsVJZdjEN/ADQMmCpRVM0LGKkoq3kthuI2RKvwDcMeIPJ6P
v/Z5zvVq8KzdCFyJ5NedJdrTUHxCpXGTRiWfx/5VsXDSAoeMIoSvWaVaT29Ac5BoHK+t6JT2QgVO
GTqqdSkS6um6d+ELqf5DIAxNwcuQra2+0hCaHfeBp57fHmrDRQ65XBuATuClJzcwYQeK1n9QQBSX
yoAWLmg190J40+w+i7zhypUHieg4oEc2ayfvmbtagSIX7bi7AOAZMEXIMlQrSukypoDbG9t4ZrHP
sCN96UY36C9sN0dmCwxnpvNiTMzexp6FHIYgz7Veh2y0YiF/Rd07rZVaHfWUf5RDOLkiVsbo+ki5
yL/BLurQ+PTBG3GZD2YHnP1zBetlcClVswEFI/dG8+FKDTUchm8yf5eL1Q+CjVLdq0iQHD0jWNxJ
4DwrzOBmR62u+VglvvrCmKOFAJ2OzG66IioIAeTmEq8WwlYvmS7J8UCvCDxpljebHGHzTcstfTDv
A7I5IZyFCDVdag+fueL9eaNBpQ8PAT9ZxZJ/yBbxqzxD9apVcwnC0L93Ow4YqnLBDO9NTmGKFEhi
qBWtQtZGFjGml/gKnYVi1Qwow8pwb2HoZSHRjkgC2YMctsgeNw0uMcIM/Htl7qlAyouWeVv+woY1
ZJR32odzJ4lpDGLtiID1jbJnLu3vapKgYnrEjHglpZYJ0z7nJfCeYqsN5dD7k4VJxjPb1a+2tkUP
1ak/6WHkBkwLzkL7fw3Z2x1rSz5nSpDnBvS33I9MvDjR3O5wZ7wpJ4SV7G+gYKmggEt5CmZXambC
C/Bts7Ls3ZN7gVNUSwBqe5AIlR1xr6JOmNbTaToc4WTYVXJ9qb3Bas9Yfwr9Me654jA3+CohRtFa
/Or2UWWJt9sIKxVlKuB3MkMRWHd7GITvTOyZrVPxMeVJFFHOBhrhDqGtH+gKsSq+1hJ+mAyL1m88
eu2AZehIyLuEAghYwXc8xbDePyHyWfBv7pTTjIpAJk30+P5T6ityueDrBbQ4OdwmA/w3Oyv3sBbe
E6AMkZm8dr/ywOxbx4YTNH+wi9IbVcFkekfS9hB3m/n3KkvgtgII4yi6ppMbw4MSuWN3fDFSykLF
eAAiBEHAbu4JX5KPsDoLpJz6mYKxm5HvoINS1ZmNtDJf2TgW768SB9KE2wQmvJXEUd1MnLDPnt5O
vbQSwBOmXyJdZ0RLhzrMCHqWDPA2illujYafUVXWGKMhxnofdExzX3y2svmJ0YIuTQyEgrHFHTj/
wLQmni72hEMZvdRmM/diWUwl18vRP/KVqEzqNv8EYPUY4DzCyBBDpq2YCg4LAqxY35fBUv6Rc5Z6
vV8jX1ukZhLCzVleJRGeu4SUEu8pr6xNWvRV87p9I+J8l6AjFsF0qDKTraXSiDz7D0OZW8ekvDLR
1ijVjjsfqLmSwCxjeWLHkV+YiWMUt1K2fz+d8vdxwk3eOVcyVCZ/49h+/u0g3zZEL9WXE/Nv9Y6D
HPKqHp0onnZAcvh/sc7ang1PnBjUGne63nJuDqhbXQDFuevSH7fZrzM02SZ6o5jQRKG+XSvjhFmS
GhejvKbV1VvCc5Ka2QnmGFmufCNJFQMo3S94qQvX3Qk0qA7fVItYQ5RHOVimfS5PWgKG9OGbSrPa
pf9Do5CX9pz6OxCaCS2k62YCbGxZcaOFJKRhBlJHkRvNh0E4JMsW6OAm4eMm4+kFs2o1HzC4plqF
cBvVMk5mzJfCsQmMu2iIMRfhjDfY6O22kldqDzfGzNn3LcegHLnRdEwksmT4HyphK/xCvLGlXL2d
JL5PrJgk/X4WfQNh57HJTEWh/VqdZjLihlwq7OQF5aI8Tks3Xhgj2AvUpsRgxGfeJNG/atxEdzog
3NNQ3s/GnTdwEFbIsL4SziBe65iabw+k49Q1h2oqLILKNEgzyoU+ywIGQiH0B2AyarptUMey8L6p
mcbpiYSjT/PdHzDIIqeVY+LhxNDI2hkpW34m+GyBOfkJGV+z8FL+xuNQxNlB/S2R0KJxQyB994RT
jbDby/fQhRdrdU87Q/N9mMqomyCIefNu1sKiEPo7kfrSF2w7YRmGhJRgaQ8vTS5SS9rZfieLNO/c
Hqs/1XZECBmrD42rzav3A57Wi9pDu7V/gChvDI7avCAhhhkalNw6gSryqp+yQmWSYpewJ3ZkpI+W
Sd/VN7BNXM1cKqCGQFX6lpXDuWo1soD9XJPQCN69DA9NnG1Tlp8sAYwadb1fNXzUcrQYK8fbx7pu
cA2rJQ7pbHRFPlADP8mGVg0RN63nh7dwayPKc9BCX7mJ9A5yLNjmgYohqjz42baJnWnSIStJ3tgv
rOfjZwaQtUXmiqx7TmB8G+z7TMlGR6veOs8M3MU1hIvGKwv6scpnSyRNoM+2bguPlAdC+kNS/sh4
Nhj0ES8/pn98IOfl7xv8CG0zYY6KaZjePsfN9YZkYuDM2FrJd8KneggdNNLpd3ZPDVnuC1Il4ffp
o9NXoGjL5RkqZwv1ZkHYeKgP4+wQp8fYueZPUQKfvFP7ZdVCOdoPT/BkD0djD7jQcV078o1QQkKK
D5SvKeuEV56MD5cKKet7nBrlId7rJvED9h3sCFHblpIQy2mHCanRaKi+IJFH84/1bQ0WPE78CRRR
RFIBhnnj+3YJwi2tiSwbVDew1Krq6tYXIVh0kECx37CpZ2sVy48MymYF5mmkAzBHmrzdx5j1CuyO
p4I3nehJKkmwFcMHrDmirifPp7yo9JuWixQ/WHT3VWotj3M5K+BlNMopSVOT/gtiq1GJFr+M93Xy
KgKc0HMFH6Yl3/1zoWAKDW7Q1hO9yh5GBdvYOX4vTLhPNdftb3RLVcholvJDjb6418X/AnOQXdvD
r0G9wwwFwGmwpEU6cCWbyTBR7NmiGAR0nMbD4mmpvyye1lrypiacFqxIBzQZi8HC0YWVfkvXSxKM
+QCxuEGJRnePsSGzKt/aSOBSmW/5eCh2ZlNs4EOqnh916vFvX59WIK/hO4yB/ZLvAxvtt2yjb2iE
Mf2RXCQQAR/j9SYj54RQn6T3svXzSKbkYRP38482re/bzvqXyc8EJ+GIhH4m/lf9gTmoRy/zPy0F
7PLnnRtfEpuPy6j5hl7xE1qSLJW4wGXSb+y8vCISJ4mKBFvZNWEl9TsmDwhzCD0xmgSWlyK+7w/f
kEaE2/Pu+JuC5LNeP/Z5VDEeH89z0smqfQdOzPgf//zpWuitTxMABnA4yZQx9X2R05Ojh7wZ0Raa
SURkNMETlkK3KpBUfxzwbQYLJflGz94I2T7x2vS1U5f33223YMFm2deMUPdJEcWPl4swr3vxZ988
248jWj51kR8c3+Wshv72h60+S5opYLVLG6HPP/iepIGeS2haSw3BMeoWWBcGmRdhOSJ7VyC0R4PJ
K7BnVEwSXjY8A5o5pVjtgqoLAJ54KhBnPtEnvXK5woprRhzt/Uwf7O4OFz3GIjCzjv/mAq9VGbUm
l1HFuagucgWrLFSJgKC0UiDIGEvnf3K9Pc+sZB4EKqoyQLzkKmxCe/EfTf6QewVPPNBqTI/9b5u9
G8c6NABLHFYtumremO+cLeWCZx4HtFlAJZ2Ne22hjr988mgF/b1yrUx6vHxYHXyH+mL6/te46zJF
Tjw0jwKC4tN9vPnJwrMM6RrgxyXF94arCElMsd7Zyt4FvDDbJZXbsByovjD86etxoCN1VXc+odEL
n9skvHU0nd2pDReV1fbaHyDi5kEWrYGZX8IKFYFoQma7bOR+3glazNgc2DWp2a/fr0NA++2au6hY
ji2CYu2gI6L3OcZJ9k6yyuQgCR4KZWC4A72xP57on+2DWlCxPj+zzpqwhKBcSLy8UZmwlnThn+Gn
5fTQaQs8mlbPlPFl0As3JUaTSQVDV8vHM+7LUy2hwMeSF2Mtl92yX31zY3+20S/ce6viGhQKNWVu
A2OAF1M6MdizagzP9aYjl1uL9pxoD1gWyoqooTqGRpVhuuq68HWKaavpp4hMgh3i1vBPlorlTv4w
scJ7e484u3BRmMycYlZz1LUrwoJ2TxGO9HIceiz47VL8YzDySCptoI8oe+5jTPm4asFaK4nUw7d0
hQjrPXCF1L0xSgVPDEwf0LUdT6yQDauoXiGl0kKRiVLt2kEzsYO/+eB+j9gXOhy27+bfLFxum4na
ife/+JICfczzi90E1hTxkbFTAQ3QfLReAcDenFvJezSWSH0hHf3hbFkjFAaOE563VF+0r06l3AMT
qCaov+RPbRi/ND6cvVKBnmP51mu1gd9BLOVMyseT3NIbQw7NX3UgM+LR4/ZwKChfHF/jxRBSMtKY
Mw0TrKQSvPECCqFOciCxfcWB3eqVUw50iu2Vq232UKtK6hHFs7ixMbnQzok3/2lcYLF3DkAAx0pd
Jl/XKinY++YCxSr7W/K2kwUC3a1sjCMXu6bExR/Xi6wCQDnpbLmXgRQVz02om4W9BBjm52g9busp
Bw4LsWe82ZA4qhOUEviN2H/Q8fc31Cr4BfMW+gOLg2ULy83ftYp3pFKVNVZSMAQv2Yu+l3Jo/Bi7
PjVzqpN/82QyWLX7yj/iXd9IXSn13KXSL7vsXerGnvj2KRJE9Uy6JkPh6uwa0TeItcoLCFKODnrf
MOWv47QD229voiPwLeYBQXCRfCd4Cy4tgDUmcHOOJO0dZzYQlsn2g3v6a+uAch+1ssjqrLmraABm
iBH5cVapBB37BiHj+nCJCxra8zDuiQnKMOtjBFEAn4sPIoh8duTwR7/hQ4ao+3SE4BFvqrddlKkQ
yLz2ZhtwKWbanygSnpv5j5OcFTXx0AQgKZ/OGXy7GuIBrRG59mbsUiquXk1iGefiug3NzlbKV3xt
T/eMzZ5nEiGWBRgv41Kw9Mf5s572qDdRyUtQAA1UDbTJCpD/cKGdMhVptqRlwTI9G8askDiERMCe
PcbMDBANBAstMJ3EF0OkZvZ3o3d7Y5rJDfL0A5eXGywprT/T1MkWcIgwGMOfr8ID/9YrGbP8ylEW
tEFa3Xhe9It/sSuiWO1f0kTUkIB0nAXYAnshIIhNuM4auCVrQHmdRhy3Xv9fHwp/W5X76znnz52y
AYGdUUsnM0tJHRm5yHvqphjYjbM+YD7QWl2lt+cC02Nhbv+vXMSn12HLjATL6arr0lr0Blc8WOxs
djRwinfrHoN8IcA1TT/CoU3uEHXRrofPo69a2+xEUmKQICM6EYPDTYXDx8U3iY+aGTpL2mVuvatI
CSkz24xGwAJgVgJcVZH8ymrPZwlbKbGIGzCKs4SOde4maHV6oXL+ne6VgPqPOwFFyL7QqwVPBcn0
8FY3g4cL7Th5C1ZN1+vy25TG5JHu5hXFa7qQoFkuLm6XOYRfuEX+gZKrUR9O26d1jyx30O2QfRbX
JabA8Fltw75v2mrAs83lA03hWckh/lPTlcYyM+IClf+YNlg/u7qvjjZG+utZlL0E6gix3Ttg5rek
9tr7xxABsFnQnvh+LqK20D6pLU9G+Lp/0lxEXrSNyj0RSdVsTczulnbfdSh8txPUSsTWmZFa/J8c
7FegFtWcxTqtkK6A/MCCLZ8t0BcmrFy1ggfkLvVxZITrpteoq0C58+uVTZnt2OxxbOq8DMlZW1fJ
YUo11/P1SuePzQB/HxEwaMvw+ff6JzdlbLBDqBpWqMSkyswV5gd8fgrkrJEgKE67STyOrFzka+de
DtbTRlCz/i3eZUvenHwXqJly4tUX7+or004rxSUBSCCo2qlyciypWs3hKRMAkyuU9yCRJP1Se7Kq
1nfMlg10J4pqmwfClZtg+becmV4+iCf9s5/H/CIea9P5QqISG829UvrbC4QI4AwCDp0YLuT8A83c
gcYn5B+rpEwsMAIDWbF8RKK/xcTFjZdYnUlqdMVKB7cesUF8s/CHwdTQB4q6PsgalnyeF6PA6ewY
bUkLrlMKVR6FJn2tCdKw/UmoR8Xcp5rdghyZQabQiaj3Du8nIy/mwSzxDJbM8SsRQnvt4fiNnq7X
UcshE8AG9wfIPI1aTNsB7dc/xWjK+HAvh8xmurEWtU9GWCR/3lJoHlreiPgzovJu8hLSocN1JKuu
yQAyGMArO4R1Wjeof7XR1jG7Y8xw8oj4sVvJjRylAOUsG7n4lAhmIHfPqnnLPvqY0RvQER9aZKRR
gBlNUlIxDuNSV/wMjTlJWaX3IvDBgFUSc0cmEW8MRoxNf6dAcU1AhPut7/EUBjhHrSIRMMBMw+Xl
jCEkH335Z7iZe1Kt7Fa8/dYXEg7q4KYIWrGDdHko7akPsEMMeVrXuI9dhNc6mK1q8/iZ6z0/PQEn
8R+zltpfcABUFn6CmZvOvApjrHx4wXJ9+In3Frpx9wWzbulor57zPsASLdkwQHjtoG0KEZ87LiNj
vap5oXzVv0pXU6F80S7N5k2L/4lao3QvLBdnpkafozm70Stk9uBqWquy1XslCtJ3VMFP+y6DINyN
35oIUVtOrw9ceBEIKaIFZD92e2L+R3MC41EshvIeVhZTKMPs/cCiBa9mpwhFo1Dn5G2lGtoN8jId
wPF0od9JTejPoS6GXd1Ypge0bcgDOYhwLTRoqoR4FCIavOWIsrTDrg3XRuK6kxjcE9QvgnCY86bZ
BvhLJDOkvue609ZeN2cgh0c4Bc2dHgWiVmJOR5/dvhXqiav3LDnrBU3YzNdBJ8OeUaxVy5Jbz1K4
HvYjE1/2af9d79n4LgANxFKq/mpSjQFPELVztHxPHgstVwtqH1ctkyvxUGYXlrVrr4ZvTXYwXaAs
1SifW+ii+13GaYoJY9E02HFkczQg15fIsTORGWgXy04G+Ca874pfGjsfc3lGV5WNCQUIVWIthvAy
Ct8WHoYBGAv4l3xU8tqfvaa3TAaJO3c3+CcD3nKNHKpGWAyt7FsbBF1lqCwZQ5uN6ElZLnIlgZnz
4bGoJOnKdwv+ojiWclOyLHvO4ql49YyyFnY06MwDA7qe2r2d+8ZSdY8eMuoio0pFoHxhZSfqGygi
vsG6wgSVMFYyVrZTmAuO1CPbADloWbFwXxC5NvE/p1IErNX9dDk/ZMYxll0yPw92kwYoWcjNQdO3
IYgiCqWuy8koLPDHpSkt3RFqwIfUnjFTt8tMKDTQTG0wZ6SwvLOn0SFuUtmqkYmsDuEZnSwVD22q
zkcyiRFZn5QrGl6DkPeSILvP6OxiMkTRQOIqzyGe+PUJ6mzSpkwGb0NbIWL0Q/oHDi4KivPP0JD/
5VFWy1ngC7SOEq/d+JDNMKwuP+jLv8nixXjAkNOHR8q1AAGAGq5LGJAQzROKxwnOAqNoqldo4gBN
0KhuqFiikljw0VXOsX0NulQmB0ZA/mc4A1ks1DjlXyUjmQXDbAuySDC3DB09IuOxWdPe6osqT/bD
1we8IXZKoHdDQ0MkMZZkbhU8qt0zatV23lKCLwScZ9BRNhMgpVqoBMUjat8HIwXOhsr0F+B0gzuE
sMQ6xzuFynW7PTWUweahI+ZDfM0y0LI46HzdWtI+cE/bTXFU6GS0Tw9fLoRacORCqY6oOu/gr0ln
lUAP7xyiFpXSOmLYdmbYn/JI1wD5tw7ND+12upMQgyXLm+0bWV37DYNil97oFIl3XDdNhb+gjJu5
piCk8x03Y3y6Ye/GJTTLSa544AvsBHrHA2Ssxu+y0GXMusGpc6jdc78+xO1rNTlyKWaA+QD+wSyr
gNYa5uMxNo9JsD04oYqwzbYBBOvXMOQp1dy1p/htw/nJxrBG6TMdWAiA2L+RTZegOv1hky0fa5Rt
Bb63JQti3gdoltsgD8+3vHj0oyw1ROOMAgRQbeDCW0odIMik24ctW15jeljzUqsI5O0eeJXRpaWS
lv2se/8FcjXlSgUsFQsYkE4OPICKF6lfo0cNha+Axa9yVonEtwqJ7qlhqnNri57buSgco/DYJ99u
miGqtwnfxR+UYb7TtCVPDy1L0IW+rblL4NYqSsCIROM4VKVQi5c9cbEi4Thl0wdUAqSfsGlZ2N5B
11yIuND6pKWFbRszmuUgjQ3mE8VLGXrm3746CMDeiW7FUUuAQfiiPsYSd2k3AeVis86QGhRwMFFs
43FTCPNsK+HFSeZ7H0u1GmISTAtg2hG2xaiHM5UNbNV7rMlp600kxdfzSj/9Lt6HcJ6nXFmVChaW
qdB2HxHAcOHz65h3AUJZQeoD/ZHKIyI53pQXM/9f7WmA4RVx4NwqLsEZuf4wqzoYeyMI74ne3HsB
lfbv3JgkP9MGW6pJj7BgALDTPNSjqEwO9P2ZsaoOjLP2/56CpdtmuPTuUo3yZh8LdPTrd461vynm
ve6ggZHRvjlhvVlQ1W28jRIpvZwMpSk9naMACZ+9+6NWUxiubt1KKBEk6Rj5TopoXV3zRPpSm9Mn
p8l64S2S7gwl/dso6SEaIUTAs/Eda5bxQ10+pDpo34uTHEI+yDEA+TonKYYUxknm80ARC0JJO3Su
j20lV2UOW8VPoQ91MKm2eZ5+g3CtcZT0Alph6Py4L3osmRuE0Lz4deyMjk1lKKt8SG2XlIVpFiES
qlwo8rhVlq3MMJI4g2d3+0CnJUAUBe4HEA+IqKMVw+IBG3KpxCm6fEQCghlEH838/tjVJyq7xNpd
iHEm0tVK5pU5HVl0kUDrpYej9rYCSJO40/AW18JkLYNiL/hDJJ6ivrCGo+E0c2kEGKFhYVvmLLcL
E1Xne9tsN43CdB6rYgMgSg9lX/H3R/E7RLbQUq5ivsBkqlaqyiceK2qxN726B6qjNs/Yi9nqSZXg
vR+91stiZBpy/5nQka92W7lIZdbHewFfdFU+noBdma5Xc0wTd4FYOvpQsb0m7/jKccdN/wLjswxU
gzl+Y/sAwtlH6eO+649TsZ7IOtdX44iHv5Ems5Qoc+UIjkcz/sNNPwrlP9X8R2cwb61CmFbuN3Ck
JoCBXw9XQ4bEX7gV5WBRvFfJIpe2Z3BvmMapnTL4t4l2Qbf9ihmaUbrmUSkkD9IjBO6L+K1n+VDd
mQ4RWIbWaVzgrL7BaeBzqY2oVJs9XcUHeNgJw4ajajK/3yGh8CGEHN7C0pJbXGhaUbNX1zffyCuq
03Z3pEHQBDfBX2d4OCpv9dH2ytIxWYaTQGVoHPsSGdloLIZ5TFk/5QE9yoOEZkPCvlRJ1ecLYSw5
lJ4NHQTxPB7BYL/UIfzaaxng4r1EDL3p4iRVymVIH1IqxXqK+b/8IDlt4BOVY+nvdcp5G8etXSr5
GHI+zYU9v50LmOSY1/kR//cVvSlOwosieUJpfTzdPWn3K3nDMyqs6MTWErO4qMksqsZM7Tb24xEz
sBgZdP9UGAhu4zjXxzpFpQ3RqgrKnJL0gJk1gcb7ELXW9IlVgOFCObi95EWDZgrFNBFMnLP3SviX
F5JBDlkaK1olUo28e+W1DttkTbTecR4ulU7aBrYQiZ7sGJ8UX0pm1nHe9zrFLHX//L/EOZ4RwQb2
HzxgycVQL7MUF0ch2brxdAKetTGL3BCSanwjaMgdSTrIbNCMVl9+NpMLgLqd4SNqitqk2D63y88j
AL8qD4sJoJQlVDDjTNSPkN+mWNg3MTmseqqmaFoc90zslOuQKjP/99obdTHaikkc+ppdngAo5WUD
6DjxuVCnZCXfCmg5YJrv3zpJ6lMdFJzazaWOafadske2UacAlNTO8db8PpGeCy02js8AtqtzXvdj
eEZ+240m+aiB/kXZlL5BDCHrVScC2gfgxUBIk3UU+VOvCl3q6TtWyG9PpjlXtb5EDfDvvrcSZKVm
jhrmTIHCAkZH76yDj9eE53nP6JG+Ik1Yd10qHQ3GUpybQ865l0s4baGX93ymbae/Xg2RFTliAO5Y
ohPR9pcnWgoqu6w6Dnkb3E12/ZwQqE9Vu8HJH44hJ3b/mjYVAcZCZhZjjLJZbaxZ6Ty7X8HXl1qC
tIOIqhCREblH/LduxAOkxBgCg0ikA+CwEbs3GNjir9suVwL+SSB8/m+OJdGaNm9ohndIsGAh8eaA
qUwzPqg6d0s4a5VNFtjHQmM86oE0YUzD8diGkU0+TQ8+TNSWBJZ2Wgdj0cIS9l1rnd7tINcy7QS6
B1lMWdnOexmbtQdmWKUAbRzLCLj8UH6Ye1Swg9Z52B4/+PqqgULm2o7ZgIzLqRDE4DDe85oOIn5b
BxFqnoM5c92d/gMilra2hlNKkO09+qyIzvrsfQiAdB+dwX+l8fSemGLcrenLsZJN0nrXgpFRmaeJ
iTE8InjQEwPmQ1y1WFlriKEbLapv04BZHPXqucHRTd1GT9UWfoczGjaZUIEwiCMtgKg+eMnfw7P1
HGjbv24A6kp3EaVv6CB5IWwjkSh8GvwSEPB4/fW1iUBRN4TBhK0xPSNJJ839XHsHTZgRJVJ4G8CG
A4ynBAYEt+adLi5H5okIfjgtC2c0z98VGuCE5AWVBIEjfpoMEXqFq38CPSZXHVd7x82xOlvCbskW
4pcE9aM7OBqNoEWUJ4MH9C3dIqQrj9x12uhC2M5fKg/Z4zLMdVWuPzdbSzeuKMtS3e5dJi4bFc4S
G7E+yFo3HFOsJ6WLL528PVa/Fy0FZUASyONGAFlkfbxSZ2CC4rBaQJZLi/B2ayMsTXfalpbwEv+b
MJz3y58FCFEhaLRkg4nChKJSx+PbJPhM2cGJO+ffZ7BUKMU/9g4lvB2YZKgF2sGz1gIKF4AqKG6P
zjpBa8UJ8Aws7SkuchMIv+UCMeSbkR+AM7Z3vXSifFEVgeX9MUfgpu+8JIUmsnXcFVjoLEShnTtO
f/ljjTlN3gCkA7zww6l3my7wyNhTcYN6+aOLAvNARt832QQwEq4EnvYi2iTVdhPwKPQmshIde9sk
J0mjgc4bqcbidWb9zBU1oHlfYk1TZo6YofRqTVryDSgmOmX91C7/yP/NwqXe3c1GNyxmvnKqnh1D
Op8RPHiCSPgDgY5G2D87rWq0H5cgj7R3lLhBfq/OsBDKftywrdcLZ4vJbl0GTbVCiM3+vMP23SDD
rJevJkf1iFVuQYxwB3LNttiyLVKb3toZYSIt5f5lhdzx6kRLTYUqqr/svLpsqRI+//eJ2nDATVbG
R8Zxs6+Tkm4nsmmCbuQHMMAn4uYnh/T0fmngaxykKh0dR02Shu9FECGMHhLIA03i0d34pyzFk9KS
0sJ/EtXH7VPzMzGhRjKV0YqcWhStt6Z4OTWtO9MDk2HXhg+EQ7I/bKiM/PwpDEbXlKYc0Vo8GpUN
c6aJhMafn/5mak3+2JkeC7vPX1b3lduJQpQ1nsPf1I372hwjop6cZrWyHtL3IFySMka88nXbSX0p
z/Fze/UXcwPPkLe5scsZrJooYu6W1FLNWmjD2TEAVvDPEOxmYWimTG7FVlnpf/7E61aWH+XKImX8
1KeJUlUJIS+mriMbaTRRreouAH3fcR//Wu67XkSPIDLrIpRXKIKLeXvcKCKx9n4Jx/IFZaihAWoj
z7kLP87oJbLzxkU9TaH6z+Hc/HKUGU+mL5uHJiXgjGAJOC3GNJDPf4ruFZLZnGvFeIopbFKJXzP1
+EduUZpYblzchw6jy34ySdKSYFL44TjXVzTJF+ghCY1NbuVOqOhHKWY4Xqll+SLPq7FPVma6NMiT
qfg9znW6s8b2skYRJwcMw0NbOPl1uZQprahWRmiIOgOkKOE8giCab2dqYOt+505tEDXtHTmENU2u
TOX6g4AU60Sf8o7vUHcy8sC3m1Q9pX7JcSuo7AEPpDDc9yrMcdWpnkrGOf4UXxF/HVY3D7YgY+Gb
sOvYt9Dhh4jroRNh6VdfOoy33mAAEs9vMtz+dyhCKMgKWawYfkbtV+2ghvQF6zrL5TgX5L0PY7YM
bXZt94hNqHXVJfqL4bBxywAYv7YQ99HUxzsXxMydlVmP9K5RE4G1WeSglKqbPGlBR1cj0E6tYUCR
3zFWnD8fhvR4oa169pZbs+/Mbzr+CQ0UhGqtORoDcRcuH0rLyUyiHSeLTBH/w7mkgAD5oR6HIxU0
xjQ7mfiQPCHf5vjKcpWHW4tiva/hfEiP5x3ndpbSAXl8SCoG7payN28NxTkX2ax+Y07xOgyHYVua
WDbEQTo9Tn5ECFOR6/o4Cpd/4EiDPs0RHZqeN7Yuuoe/nPBzUJrBbId0V7MXZVsvFMm1nLnSYjOt
1u1S0O1+DlpTbBZ6Ss1GuCXwxmOIPqH2xFAwkNL2qJfjABCXbCxSmwgPuqWBGyrsnfA5/XX8x1Lm
YYoVT5x2BVEhnxsZ+EivKVgFAwviBnOgjAu1AYeNM0EjAxR/QLRlg5fetVktjxLB1tEDNA9F/tAt
/JdfVH6ViStCvPjPibYeVhhO5KkvkDUHcRtjjAu1mtqV/kt69uLmItw3tv9eyMUUvsvPd2QtDUJS
z/z9N2ywaWxm0BL7BHK0edgyhmKSSlz+jKnjk8NSeEN8aHUnqaA9SDMN/tIGMy/vJPYv3t1curqX
9TtVQkaavTKfmrOlNviLwI1j1f3jrPkLF9W5466/89QflWr4WxYhEjN0HAoK/vAG6YoRTsReqNDv
kiIaqzC1fIsem6yFt617Vy3v6WcdgrrPD16cRATiafQ7Vz7C0e6sSZevnkXboliGvuPm4qgsfXGo
ctvpI3ClETJaVYGgQYFZ8ckIhHkp/v4sMnYF3iMgKFo8Gpvq8+y46JTUbqCSjCeWXukHo+jVh1Pb
6Ne/ZGAYGQQ925B5+qYXANnajG9/mjQC9vdz+6vMmQjycAZh7sqwNLD7smI2le3Vy8+MyuVMgAtL
SHIft9yPUkAthkTu8ZKMq6wtPyPyKwv/lOVXahVXTApaZiKIwVLX/7rFkAehULDa/XPZITECnmqK
y/LYbCmE1l0F9WXTdYyVwKYBMrOoRZzhA6ZKmAHF1fdEODDQccj5JjlRt22IJJfrQaXzpWS6T2vb
lptAh+SebBt4IxG9EUungDld4YI8TqQsSJq+Qp4cZ80Ti6a21Omjpikw6q2ttyuAwItrYQVrWmN4
16Ama2tgOy5urd4/iXm5/e0KBc7YNJeunYeBtD5XyFfWgQ2u6VoKLkqGozZxEkt+AIHCXYQ/wjsE
CVwdiWhjHR4C1uYpEq89u3qFoVwS1lttTSCAncm46NHc2wqcnGShChxAs/sX1mw7iaoJYMnclGrd
x5Gb6nrrr+Mx1lcEa3vbfq8XmqdFcqWYGEn5P3kiBFmX9KO5HBrvfLsrXnrUKy0vNw3l0QpVXgxv
FFq8iy9EjlO0w9N5Qf7WGLUVftsSIv0qSxcUtO59nOierZsFJTouGfOhoS+r3atGQg9SQizVwws+
QR3zOFqHNUj2ULkQ0Ml0PlN0bYQYtRU6ZJMA2DgMq2ZR6wBm1VtMPbHtLQNreD9KcaHFIPH9lom/
+584yuxTidt7fc5UUnDK9TPifv6M0o6oLYwiuvuHspfJoyUhiqsCny/WfdAVcHiqkYlmEyvDvSY+
TVctlfmQcyVjYsnpflb2D1oAyBKjJSr9tE6MfDbVYj8SyGzONXKx+0N2+F52NH9E9js8Mqw4OBWT
aGy3PoWMMaD24uRhxKcjlg2sZdN9/8yXIBPnNS3fJyPPLVoaBjTjZQv+BN7kZ6U9CannTj64/edr
rz8/funB34bqTD0k/Mk5X+0IlCuj7D4Uw7JUjGFgq5zt7syaquM+LQJaGPMKkiLj8sthK/14wloU
RV0uRLHAWOO6GSLaKdarCZ2Q4COXKAd9DR80S0yBxP8sbTeZ1ins77wxri5DzWPML+6ZCoP9f/5N
X6CUgbrcMqftzNKBLrEtnSE+/Cc0aIvC9cZZpiuU1uyk+0wPQBX9GxKdPWnM6r4vUwpr4ZZhpC0S
KaPEh4fooOfza8fYY29zE+IAiSxniEH+5huLnKtiq5DisLmMg+iBu/AC8RDFgsSRoGKQJiYqvvAl
8Ey0xTn0Aeiql0S7ScsvPphpmHqgtNQUYxC032hsEP8IjbljhxdMIUKcYCKNe4hACTmOa7CYg3Z/
OPHTbYB/UvRfuSOOv5sokXbKcuOhpS63DBwpg8vP7lMpq+JD7XqVdyJfihnz64Hc1TvwBzF6PwRQ
YCCArqGJgeL08XRgmUsbKPpihq8DhQU7sHblwLEDBmLiuFaCV0SGjGOvwcSHUjINsZX0HEGDSA5I
HhL+PYG9+LrUMNy/IuoilVfqyCCJ8fiE7CuUYaGULpQAWVEzNetZHNpwqx1RwZ5AOif84XxK8EXs
SwJaIemzzzXtneKzcU/7gHGVcWv8khkSVm+RyG9gKXogKdjXXYI15s8C/Kc7U6guLBaBFFPK6C1n
zwievEpOnjmFzE0zWpc4myR+/XFo38OvECebR65R6YplssbU1lJQBLoOtMiFzhcFciNa6KAqmc7E
SbRu//Xrkz2OAcCtKoZ+8grTtJajoUoxNWqDMaGSH9LMi8q4862J99czkRq65IbEYbWOKjPD5k/F
cei5UZpipM2h/eSGDGOt0mI4uI5Dj0MyLofl3+8dNj941IE64eCIOkUBJt+a7fy61KZRdjHagxz5
rpiYz2ngzIaN1pdHznzzoojJfC+LghPTUNlAcawXjIjgQLKT3ZCWmgYKZWcCAGuydTJLb/hYIPiA
DLthi5aP3EENZ0Lyq2/Ey9Sd0TTdQo7mS22t+7A97sQUOmnRJQzH2BLSVQRAO2Z2L3K/GZg14IJx
+c/Gm1am2muikP5vCNCeyCCj89tNi/4MAfVZ0p9OPWVwGAtlHcHMUnRYdel1N0FNNksP/ZQKc7Fe
btdzWlCUgcgHATzper/vk/qGJY3gYW7RkM1DoSC9QfOHwLfntHFhVbH4DASIY2AfO2NvztkijOsa
bY+6gMe8q8rnJRhhXtV6xdM8cV3JfbexoRiwVtZ4gOKAV4gK3bfWZeBRuxB84LRGJ+ZDzkoUTRFZ
VKZuGnOgTb5LVjnpal4t6G4t7sVE7jVzPNw4+E3Q2OOsWM1mCWKWVjljZrkLoI7rvhzP4AvKd8pu
KPBHvlKTyqXJLoMpIkxNA+Vf8LafEFlQ+3otyKM8a86HALrwXV5wnqMG0gAi0JBzrb1NZIgT+foR
J40477E7iBv+8t1b+nop+U/YKRUahRQ0RcvRKc1YbnsVMRsz2g1xgIw7Uj7GFYQnH1OkjoSZu2xM
Az2YRFYZdUfinnzYmoHKDt5hHKYCxw2nO/QCKgYNu2hoVOt4au3RjIDn4UKQEITTTZ3E2qAeM3yO
WDJ06scJuJ1wCBI/VAzUpGILtlVAOmhXxvjX+wME2USj/j+i6+ySrvis6iIUukF1m9iBYIr5K4Sy
OuvCM5NamKlm8xgKfGPkmibBywQxlRh5uhkpZESQWGBn294H8W88K1Rm+tpSBsr86Asdk7a/OPSZ
T0cDL3NP9tEemxXH3Ip4buKs9jvmpXY61RN/lmvr3cJPgp17tDvArXaviv74zz2XvapmBoSf9ux4
cDt8nQ8DLyAPO+w5fcPV6t1gCsxpXvetcHM7vjQg2Sm1J6o8CL6UluV+P+wdVYJXVMg2gA+xbapZ
n6rQjq4dKpmthNLHI//leUt4zt78zBMD6hdBgTi7BHkwCRmABnGVzH4xhuPLUpCNJvBWrVaaEfPL
af88JHkZKr0O/45aj2XkLMtRnJ0RgLEkYw9V5y5dm8hG2XMEGonvsd+7F95V4A/N4/qpsQIFjfsY
+XzVMtw27QRVGQ7EJ54k8rPxFUlkOKqxc4KNG8DT2CcJQBtntmkyHgyBXQf7+izmLTkiTKemkePY
6LQ/RNSbtCfi1fzTUiuM+N1kRDjRIyMpe2Siq04oEEItqACpoxX+JYdz1MufqUA8+BmPVzhLJ9o8
D3AmRetLQKmq9NWoDo/wswZCrlkxYPXE6lPAv0Vt4E09fRfuVBsCeNuBDgCFEBlylOvmtnfkz3cp
Eo9O6e1PkpL5WJXJuU95BTgUrzciTjIiBJ69kgj3k9vQW8cmS7he0yqEbmMtrkvkzlfEhjfNgdTX
BUfBYts6QYyCVNyF++9Wflmz7O8PQCIVhtTolaflGTvPAasCgmpTj7uXC4iBo1vFVUZ0G5pTsFEu
UcLOUooz5KJltH2YSz3qTQITV5lBUD5UcHGuBKANiRmJZwoBy3PL7FClJXSP5QFYATLnGN1OftJs
iZhE+3wWUjX9S60hzBYyuyWYAraXxPaS51vFnEnnpaCf71N9hgAJ1JvK5hH8Gbc+xUNseELaK+T7
iWqvNYVwi56GEsEQPRo8EMDNfwsD4erXGBN+j7lg/4AeDPLrih1BMy+QTiF+rk0SPtTgbou7i3yB
hrL26QsqFnO7BtVTMAqfr2p0IqtyBHVIiMUMHA1xmmbD8YeIcbCVjnExLTynKlowoliOQdWopQPK
/3ImJVeVp+snK7eZ7VDeY8b2yzQnYtmoCWHPeUwJcSGc8eWH7F/2K8xCsxF5Aq+LVEt5hpNcNbYp
kWDKdapT/fqdXTsd5alvb6uuWtrKAqfA4RrACNbkxaIMmcjyixX5vF1YJ7PQybSipA/kaUnFhmZK
FT2MmZH2tiKBRXU68X+ffTGHU315LYZlG07iUnog1WWimc+JyMyWKxyeer2pulKietqHcjJNY67o
ctawFFu61Zx45rnuzp04qESjjRH1oNy8ixaf7coosdgeSatwPmwSTQ93TLgJHv+Qqof24g1SfOtg
yGO6bfafqEhkMbMtTvknB/TjtfivgFuaV1d0xsI279RB64QEbP610pJiErC9ymlPa2Co88cTqcvv
iBVlqdoC25hGxT1ajhX5Gwik2MecggTFGZ5PwPDCsboDmVWLXYU7j2elDawu7Hk8tX8r1+kL5nPv
Bc8sN6YHZrZjtlM6/fy5XlkuwQO+a+d2meve1+ECpK/XmUX9D8N3EvXTIya33sGg4nHmQz6fcvDb
LIxd99p9GWT880aP6BiIwTz3pEs4RV8z25HqUkAkxUoSEamn1ONzuyXu0QrUUpSP6uaB6wzBJ0jw
A9AHBCA04hWTO6lxfa9RJHUeGIp40pAsHMMbIGAUfdpdj9hhvmsGI/iT6yCjBpKfe4eC7HVBaj6z
V0KoBo4MpTLLWIqgHTbj4LVWVGW0RanHSzuwJtwvcBgtGKr/OmRG0B9bklos3fsPEokimA+B22Bu
W2jkjoqM3tzPio8kbaEOBrtpRjkHl9whbY29E8l2uKIhQ96BfGKIM2TvF/MZcWgRTsI+AePPzLe5
YhiAlPfQh1K60oFz3usYpGdVqlnEo561JUQE3icOGudesqYVuKpAdeZJNmKDkfhNImFofnc52VSG
xXEPMol89R1igbNSBbv93Fd9QlhTfr68SF12IQh7sC44qyha+xa+aThscTIUXa/kBIBs3ULfs5LH
dpPlq1ZCNeCp6jcr+RtBKW23DbWEgd/iMkwl2jsfZSHTAOLVWS1/R7KwApLxMhIdvbmenMRggBf8
B6nsjh3L3GWOpcIwGiO4Es0a/BssaY1wt9kqf2YdPFfkteAXB7Z469TOLqQO777XKx36Kmq+Kis8
/yFgg7dQzj4KW+HFx3G005QXWc/KSgxygU9xOaqYd7iwPWmxSM9YImxCt1C1iZe7Xy4f4z03h8rw
qzkRQf2VDMQ4KLy6m4XHTjLna44yaeSBaSP/mUIeoSnJCMVVWrUqnux6I+HFCLLTNJhPE2V0G95r
kF4nxC/gxuoiJ0Ni/rAp8rUSCkdWYtEbaaMkYBq1bK5IJNUI22YjUalsNxhQ9G/ophMqFCbXiHvj
cuGm1QqbKHra6VX2GvRh5Gj/i4EXJZbkwRrZZkvn4RBSLhEZwwM6gQsamJgPuAnPTAnTJeR0lFkj
ySd76oy1Ya7VSkVj10EVY7kV86DsllP280+c08kbOIwABUTvh177JRzfO0wEMhynRwMABZQX/was
WPnThrHM8/sqZFk2f05YqonN1wwtuin5OsbJUsB6B53hINXMWJvIZjPsOEPNrXx/pLzZ4b1BBkIs
3RqeKwjC7vE1psSwSnwzHmtQnVou8zyYJvo5ZN0LHzCudXxnanz5oR/b+3PtN3xCZ5W6XHeIrxHK
7DxhlIgV43o0DF+iwSzkQFYIr0orsyuxODStRD1eBG1HqsjIdOmwjbyp8slV2ijbfSwZSFzxojCs
6cJwKZB3GZ9TjNEJtzWbwglZNEXa2HwFZqi47OPdxXLsVF0xbgVzGXnUHi/OBuhLPsa9k/rUMKOh
SCspoT6mV5YSgJlUjsxTLq1ArZmJAWmjAFmN3ck3iuV3wbE61vpPzKT6LljXGA51F6gl7lC8yaWO
ErmBMX9dBMMF5ua0zxGC47ydAGU08yq23nZlUMahSFsM9FPMzAwMR8QogLipDSC2hHDn0jcHFVDw
xyOX4Ypkh0v0x8pX6qZ9FvypCIITpHcYAuhdpIfAKqdjPnyDTrESZCNyL1xb/6Z3AQXjpC2wy7gP
SwPcPK1gxe4/adMF8zjJnc4EIxYHtLgjHlH4ZRCCQiKsifRuHDHcQfxMeYfPBbhge3L/muVfmhog
9UOYdh6FLndYb40hFlC5ebQAi1HCBLv3b9Yk9228d7bBDwAg3X/nGNcevAWVEsVgS536grQ4sYrf
6LTQaeUg/7TP0cXDAMrI7dFU3k6nm6M1SqE18eSvKr9MtyzD4x1sYZvfkmwWOTITk7eL6jxizxSo
jMirutn01N5IRSEIdAI/xt3aMaoJRR/OrjSleNsZ4FLMK5sAaOjIoG3oEq6bv+bb2HcF9/w2eKJq
HJVIgIftE4+kx9Ie01ksz0JHQLICYjikbo1chJxT/Fky37HYWgdgronAIl90E92UnEyI2Oh5B9+s
MDItmj7lqyRk6A5jtCAD3L6tsqr9yZPwJSu4xgOsRshiGMJWJwAsXlFYVdrQqB9eGYP8lWLOHGHY
3YV6I8UHyJaG1FZ5ObLC0mS/8jP2K7tPXm9GWpt6pOe6c7+QFVL72DwKmv2PYgGSwn6TA0U3UuZ3
UCAcbDCBW1vrEE2PrYxpGj1/ZOLHYFPohJ2ylm2DkMGiYs0l1cwi3dc5P5Gf7astcC2qyU+gHk62
PunWXxYwCaSoP5b4q0QkbnTdwE3fxTe/s4QAyhbC5ierGRKRT927NWeR88KF2yGjL6qp7ZyNdCdE
hplc7AgApU8YMEuuL5LguWrzRneHdj29INbRj8AeKcuwpFsuuljSHrVcyumxkOzpz/gMo+yXLBhm
rgsAjr2ygskuCrWcXSlHhQNihRvdY9KIa0sK7woSWSBJUGQq3qq5xqg768PWKRtIPYekdO0xbNbV
7jlA5VC/veEzzHjJacFhCysFK8Gk+pX5aSrBZUVmiJretLP9t8tWepXeMfkUFzG9tYlt8S+WQtDQ
w7m49dHbYdDSJRq96yd+vfASh44m4bBFLsp+T4/a78O8pR2k+0mViwdSebLsexfSVaGWTofwoly2
xDa+wUVAulMpT+MN1Q6xfBm0bjAHtbSbkqbgUxftoIYric/yq4YFz7v3Z8Am8Ugwq1TOPCOaey0t
boR1c/idpZnIo6LaMlkfxIPsnImNCwvnBbjhlQ1wKVqWm/MFG2u2ny9OJi+QQwvE5L3pZdW7zavs
tZowmR6f13Radd2iF1G3REx3omnP/TxoBEnHloYWte0jsDTWza4k0N2wkXJ55rASjAgMY8CSsxbv
bC4pCdGV2h0Gn7+HGAKArYe3aw7kWyQHTlJcz7fi5ImojIuQc7LkxeZ7B0DnSQLkrN2F29YL7CJX
5DQeJ7ST//wI5Soqwrm+lvUsV/KBGVlm7BJ9EAeXZrQ//KKfA+HtUxJkxOFE9XPlxVJ0YgRHBJuF
PZSZkmrFO+kONj70Fwrsf/xTYn+xQ9eDoHOj+8AXASKzOwOYOdKeaU70Fujgoxo/JEQQ/hiuCcz4
ub8iOAnvt6S1YS8EHPbQH9/R8FN/uykpzOMlG1orlxLvTyC/rMynS4AhKCHS6eLqwnV+bke1wBN7
kDM27WW2lR0Djc6D4UFqBhIfHsO+InAIlMsi7cdBF7/Hta96qQbhCOy97PdKZ0Q9m5NgoYEy+Fkr
SVKjftpCm+RKUKBdoTSSfhpd0YDQNRVmjgGeYn2osYsOa6fjcppGIYSpbYDhJbQjUJKiNeQ6I41z
QDfneaqNqwoQfD8/tmULzgjFcTC1vCeDiZ+tClMB9FVUtAHPC64F7IKVMxDtzQV3WNguzaVq/823
HasTOX4tk5f+9CnFisKY+A+t+98dLa5QMtq+SDhx9uLMhiNIeCBhoX4quBN2Fjes8QeQ730Tqllm
PUVDw5gs0NubTGXMiw6kUf1YETIQcWs5nsaLZ4IJiKxMUuU8lTBqt/eHJNXjJyjmrLvu2olD8Eqt
PgZXMmux512u4tqfsOhKrVoPebjbzgwH3TZVHhbMAhg/BaJfOaSHz7MgMtl+d7TWVOsAFWLmCyLy
Vrpz5G6GjMnBtNDR7FXPqU2rKnNuC4NUS8BdKJgkCItr0fJA9W83YvJ25v2WuE1BqkPPNYj3gb6j
7muwsyUi6XEyzrhpJwZSOCRZGd5wwslvksVexRtOEjofib/udQ05IwlU4gJPO/+/Sjt5g3Bn9ItE
Kye/EtgB53D9NSq0aOrj1V9EmiOMW1ryDkdmJZLRCb+SUZaxRJ4e6Znp/YkOYAYrAgeIXXLktsqN
JhZF0RwA7cxU4jfwX6PULtmMNtPndTMd5QPJ+unBEMBcEGbHHlO3MeIxbHgHDhOUoFSB+2TPbgTv
23tmTa5nPvRjmABQ+RmVjNdSvXGr5v+cw/v+tpZtXfiLT31SOx4devpG7xduUbva3m8jMCZqFurq
szZfu7Dx65HOAnvIO3pO/mCbogkr4JiNQDka790AOsDARTRCqrFsXLXDyEp8hCu7/8ZYox7f//u3
ghsWK6ZacaAhYsQJ8ITwEAx+Wb3ZdhUyF7hPNGJQjFX+lnTkX2/iZutmEv6PTTX8AV4WEu2QfGtC
6QxZAMG2uvwtddGnGZzerS25BEzTAbKJ5nCeVnVplEKqGzDzNxvH6zOjuDT5ekSVLsZEQoQ+gq1b
V+/uZeIwTUiCeuVgiDhZbgg5G6rINFhlilVypjNCmPs6VFiF9U7qyeYXVRoSZKNxm3r+HlTv3AoO
qdOBH/JnBAwqJ1swRS7LE0i0irkBNXQG0zoRsgzCnp0+p0mxqRuHq9VfGFbtV1Wh3zLM3fvPS70a
SI5992ngKHOPwbPZrajI0oO3ELOaGcJAv4o9tkUo6wVQigRM3V66bvGFyGmP9MB0cXmOj6eqZ1tr
moJNBrw2biM+0WH0WsnBmLkjTY/FgxAz8AAnes3HRIFvZPv/NeC6wGKpkZUIttIdGX68T4NOKBgg
BQsR7yj2WRUa5Ip1Vi9zBy/h2cpagXW4XZxbn+TK0GMZJhePh5pY3DjqW3NHqyKO/k+Akkn5hSEK
w429omKUlTJrEfIwYaBCc3cQd+IOAgGQog+Gd5JR2iB5sJjfW4hJxBbCOARBINym98v3rLr5/iIc
uEoGZcSAtl1T6Xzq8stnuoLZEQygPQLzDNtgfX4bwZWj/EvHfL+I77xGTsznCPpJWfiCpMYWHdRQ
6wUdUKG1tsbq06wd4KBRdNotYV46t7vwpl54Jdy4vvXxQzvyJs+dVJbQCkv7ji7VGp3klPLUzSCq
KIYNGu1RIc8aj/0HXO8z4tM4AWRFThQDPnh4wawoqB10Qbc8FtzKvpIOvZug2tWqAx/ahfn1LHQz
12czk2ffqFSGrAAnhvqyQ6fg4HZWXn+KseEwT5NnxRRa4+XYvhDqSejmJ0TqJ4nInANIkmoT3/it
h0siD6EmgsxR0UeXGqgm+nhO/JxExrec6ofAsqbI+uKyJKg64JtAfilv/6+ilstW/FDbIpNQ6jr+
2Ognm0J0oWuziDmy7TIeenfKgaof9KCeudqoMj4891zM4c5nZibYmILHS9yXWe/HtRd6VzmyRVqt
E5Vn3aouw+NT8Dcl0H7PUHC/u3Zr6BSfh3uhMNivGAZ8Pb/EoDl5CCry+jWW/dALRQYnCsXVzsaH
wnM1FE7Fnm1EceU1hPTmps44g0Z9dbvWblBCRHi207/X7CWJyspJa/PV+Z5UR1uDgJROhQEq8AR4
St9f0OzvoVc5i+6DojLvhAAYxHgwMMhY87dqMc5FyRP7UPoajer7lISsK39D2YM4tLtfu0ppHOie
mjaKixhCRgqtCpyHwRBoF5kl8pxK1DnNePM3RUnQkzzlh5t4Tn3KLvTnsrTrqB/Tsrd5UkvmNU+A
N3CU7gZhiTtM1oRpXZbdTzxGA6niQcAtdRf2yKRjPPl6tM8mCOXeum0LlbiCkyxXbXI7LjDWGaVM
+ZlNwPsRYbXso7IMuLkZC2A4ccfVzouTCoJM+AiIMu+2pMltnbQ0D/Mki+7trZePGn2m42kNQDeK
LyiRcBg7w3cFZ61XyMmxkAwOJ2UgIs7QEzfeMziyRuGoOfkhQa6KuRqoOrvYA0/lJxj5bnZjpzj5
uGvqQWk1C8SLqce0Uhwat1hZjlRCGQ0sxmo01W/XMwF8qDnGpdDkEqI+txsPR7zAlbQxuyzDySi2
AfxILIcHrMIvVzzWdy/z+qe2V4cDpqs1rX0lASogdhA2Tc7svy+iuTbTWou830aBkbS3qCRIVZjB
MMYFNEQzD9Fq6gUCF8ogMyZ70kl4XWZ0oq1F0I5U1KIOJNB4AN0oTLV1cqvBNvO2fCPd/ozstxY2
7ooY3kiR52r02QvOfbcO/ceadmYdYQmW8RZe1clTiXJlKfID5FOTCrP3/xcWD+9ZEydUc7/9ehx9
iIRiSgy7TWhHr2zyviInQpf5gkgTM8lYuijBnBlShm0EjrmyFSHdKNQsTu4MvFJuY8UXWZpfh3vs
IDGXsEPdyab1HSSWp6Nf+U+pmjCBMdPB3/42IaJfYIrOZO0O8teO1Tlea1P3NxD8qxnsaGBV2XJ5
QHBXRwmfls+xyWmF1E3B/Lqjk+AJwqCFbvG69PPL/58bIbfrLWrJH6dGnYsOEXvr2YClvrrgBv2L
HOuapqXKj6EgKvUG9aNzwKMWQXwcpZW4BXhwdVDYHp8H8d+Vrtqc03HrJmsGo1YNl43xpW/R1iok
YGilFRb6LnIzuyxTdRZbKIOVoxgTvtxwuMVpYwyA9qEcLDxOoAjTabyHMd93PVePMUie0iOHliv5
VC/Ruhc7/U6hAMNoF6siXg12nOmWu3mGowDQ9eP5azejL3vsDMSke1H4i12Vs43qrw+k/VyLXOEa
7QeFzFi/EUsa2Y1atpp2WMq2G5KvEPYHeoFnHp/PD2J9YgdboyUCcryO20uNwyCIcuHLhhq37Eiy
2Hln7jQPncZoi4Z5gr0MLjye9pRUY1vBUzb/PZS945ba3DfTO1xsZ0dqN7diEIb3LKHx+QbHmQig
pumf9wMNJeu1sTxtdQyJUsIma7gL+BkFWfM+hTkJZTtgE2KgEUtOvnCr7HdbeqV43IkTkBtXt/li
H2efQ52xRTg8Z4jVzyvEy5DLI7Plw2fkTPtjTFtykoMQJkG9OK/ErS/WLQcLKWnpJzY1y44hDbo4
ijvJubeISMkAFqBKF6cE05tSRjTv0QILUxB0bZGrkPBQDFSXgxtdsml5+8uNsMI1nHo38nFH5b9d
qV6kFKx4eBZt6T6I6aq4zDuZ7o/9a/Ye9Xvq2pSwqOY94mQqlVp1lAgspeUsEiLwhtJwBgvhaA0Q
icBGA5+3kz/nxoI5HtRHkChrSTwWHzovmD9YvRxTKeE9r1yWj6BW+jafp8SMNHhBFA97lv7LdjBq
6NYDbk3eVKqDk9BYDsKzkjVBPQ/K67kGKIBLNBucfYl65enSwpBmEJ5f2khTPIMplxJWL3TPTens
hCg67eKzd4me2z/z/ha2N/JWHuIeYC5xvCGVSp9/UlG7MuvUR8Y0IHMCWer+IwT27+R99X0Q3YQd
DaBRoTbNxim4OEvNi2F0cvOlgS0ygvattzpyHD/3XpmPDPLtK3gooJVJptRIN/4odx9p12mPjAqq
MyHBEzn4VqizCLgwyJWN/DbSI1SCtp+CWrnkMlj6uRwGctRuB3Nu28rSeW05DUVCYUDuoVdQqykx
x0YuiWynnFKiAYkZM4grOkDTz913ZcZFIf6QRGBnMBxKQPCZQDydes5l67OUeyoOdVA+aUmOcL47
9C62AiWoVq3TuBfMm9OUL6REvZA1IjhiuHnENqnLVMYU/2iG8deBml9OLOCb38/FMUAdztB8oIH3
G5JIK6nukk/sGpm0QXgq3TPlH2IAfXXqDBH/ixA6kanicmGYJVeJKDgsDVr6QHXW/UoFXzDsiMIp
GrV8KSqVQzi2cMavPik2nWRb/0Jz4Teb11uERf49IZjlonZqsZYZRifmW6wuULRJ24JNvaGZsqUQ
QWHQDmllqnv8bRCB/GQqyndYx7FZmuOgsxanLqF6MJbWavvkCcAwgm7QmhmwA5QWKqATeQ4SPsRn
vUBN23dHGVSWAk/K8EQBKQQhkfVwbMeLaQG3SdUyc9ebJZGkLId+bBsUS5hiR2WJzuAm73wTfuVp
M5Wl1EXKVLtivzMPCigQki+jNYAuvIM4QU/kZjTZ92pvmIhSRxRu9NvXB58DOniK7LI30XQNKyzb
jhcTF9O2610vcAXllXLdjm0EExo5MEm63MjFiT4wNk0Wor66vyUfELrVJjIrATPkPv/0zVJcfD/a
NHFRPOExjhiax6GK3AkZx+S8mURe6JaLbJaO78DVKOEicJcNLu55SYVa1u/eqWm6hko79bWjjKM9
aNbvoAFbrujghfub2LDzszS7G3+g0PgUre7AMkW3znYik+/eyo+BAOVjyeTCmzg/0l8GOd2XE7M+
2c6U9JwVGfCFbLAUOn25WhOIODv48ZPtrJTthsk5WiWIKTjl9HXHte5AX3fr+tCNN5JXyGPFTFSB
OPM1uj9HD8QZNGb98ArW3+RxcbP920ZZe5Xk8+zNsOS1774Bqln5TlbDsnNIuvEF10CjpPdK3fcD
vr66llNpYFH2W0KYSW9EXd1CIc1xEC5SfdnzMBtNq/6q+lh7eeJNXseLDD+1Hg/x6a1k26ISjnvU
ltbg+NjIbambJHXctLih5mlXBgJ2Wk+xP0wjawmZDtk3JQ/JoapXoOiFmo+cHJ749z7AWraspw+F
uPsv4EOfPNkDS6Mp5GA7WL1sPJgSZJBYGs+Mx+I0oXBQofd3y59Yuxi+NBu1i+BRp+JUbVa8vtx4
H9R3ZC/FyUdT1WcdCF+huDePZnUJvUZbb7hHaGZpUcxBTlFUiGXG9mls7DbM4wZFMOhZITs5prU5
yCO0Imk/N3bLGf9PidP13no2Ow7BZsA2MsYxs1unspa9FFWtglVdacuopq7CAJdP8g9kSIzDP7eL
IO4e0AtokT31Oxto4K7jTc9FmYIB/DFsBxEiAULuEKBojkPlYJuppCcak76xUNCRtfLaoNZSVifm
EGpdjVJVW6qc5yoa3O6BYWvJnBGcvylHx+Bzk8Kw+5WCMq1eFKQEsAZm4j8hrTqUWHMM5GcgvPJs
lWMe0pdjSLpxXI+1eiiHIWe9iFFnK786DRXLhq1JjajXOBD0BukzvqlssXriDq5G/41xOpF/kmHv
Ua3X4rQhtGiOrg/BwWIxzcCItGD7KJx7Vm/mYevJrZHjFPYUNdFUqmCwel0v/1gUkDMkUqL+Q7cp
52t3GZWQu915+C3umydBNvAUsJqyDpYU54xeizzM0QPSiTtXgUMqVmBGmszINVhbh72qOvjfNBf9
KReJsI8DSAzQa5YhynNuCsKUdK+iAStp6+/Y1kzQDBUDLsa3eNkh9DEUSQokg0yw24lFYMLyjyHU
LYV3yH5VZ8yhbVMP/hm70AxVlQCGNvroQVYqdgUXaped9JDI3pGIaSWGEyeq3peoVXvpUa8t+ksx
lAiaWVbNrXoXff2Op2T39+pDSUkHMfrJKjGNGH9GZJm7tZssPCZ82830Nk+xHyJ7NuEyy2IgRSfK
t5JczKQbe/+XQYOWQvrTbBc31ISluY4O+im8mRRSYLnLoM5klANBz2f5Q9gktJp9V1S6pmUhjApL
UVP6eAMf8e9sgGzqDl2Pv+QB1U+lixaKhat3SywSTioEGwYFEDfq5oenDecA/w8mBei9D3BnAxk5
9YMt0JzTCxDEoyVE1FPQC/r570Ic0q+HMmU1t3fovmTm6yk2wVdYfn6sbKKZFDT2EEkEGN1+LUIe
ZQEKQKgxywIO9c5YoQX+RxgnRGEhPA6iQGHPGEaAKIcmF8t62DWVfRWc3Mr72ugmgU84/p82wZbk
bmPQFumY/+A/myoTJOHzSdogHV47aeS+X1x5FQmhcr9SE69HXH4w1762VxW4yIq9hxvcdzGOTvGN
jxeDKvph6symo/KLdkMY0LOU2B7XP26MfE6nUhzv1AHYWU34rWeh8N3zqyckYzWq8zSeLqYcKutG
rQdEhm2QiyDG54O52yyyElfE7MiWVIVJF9lq1DTWQAM73maEQmrWYBCvD6PVV+n9cxv22/pjf3ss
xHcwZ7lO+ybeQ8Vrc28gI3uEI4nmko3T53cT//IHRfm0ashV0MZ0/lzr33n5hLvNDAqkDHH5muUy
YLccTCNQ2zKcs4v4utxG4ydgEeaFoD14sJD1j0srBILGOCXdZdHvgUkvxewFQ8hkt9tBgbaWLBFv
B6B0PD6DNifvUuB8uNJkEmbct2lFJfjPNmgUmcOG/MZQHftjSXMuj+AsNPDzs1u/n0GKXirmd+tX
lKgLOCfPPRbsZuBar0Y4pEFmc/0WKjq5op+9ex5X6jsRzap5bnKexKtn2gkwjHVHeH+rFTpQpZG7
kT7NQxr/sXEWaHGzrCvnPm7gPlwsbp0j4Bc3bbtLjc/+Puz0kwy0J7oYyaGEqDm19Bk9HbIfUPGa
25ia0fXMB1piM8kQjqTtAlM4JxEFSLBZtJ+3bk4FvRSXWN30vw/WdpL8T/UrmCjxVuntrZwSVzCE
hleRoh85Ltf0j/WRV7uY5u+zYOrTe+kEGZWKdAME+Ysa9qnQadKnxuNl6/RUvNXH1xMz7JMnNxHg
eL2pn+QDm1/kbjj8qncYiu/EPM55u56mrfZf8rJVh4wxP/lF/VlQ9CAhXrqTbcL274h3saxkU9t9
dVRLr8rOC527a/19Mczar0Fo7X3YRM5fXHuL6xwMt6c28w/6c/x9+qppmnlXBiIGqs4fCn6UShDj
yzdgYAVefQRPa2yyoS0fUeWhbFHE3A30kgRcCMpvlGmQvWGr06Q7iNvKnMjQhPZgBG+jw47QNHLz
Oh2fDawVNq7XL5xAFZnGEq0y70Dsc2NsZLJ+WBA5rfcNded91AgjGv/SPtNWL8dID1D+DXm0kLP1
asxG5RDjO8k4CyIhqIVIf2ntnhc0AbL+XwYCadBTcDnTHaqcmxLZ0l9G59rrydzRwkOnlZ7+QJez
ULvTm9R1wB/QNitota5hgKDQoMtqnDdzAKLh7IDSL5RXUZNVg6j5j8/xA8V+JCurrn5FTlwC0QYX
HKk4sOvXVBw+UPfqUMPW3yOdMY4I6t1jWQbF1RtQapBMaCz4RpjKUd5pAH/6idFGnPlMgnTWQ638
75qAm9oa5NWk4WFhtRUJKaG8ghl1FnXOP9gELD/M6U2buMMZue/GyvM+5Pcz/vsp3EHg6Q5WJ7gX
9SjcpdYEw64G9VUECRTIxEMK4N5LdzYOFATN99sPFdXkkIW1zz9SgFPRxPRXxeD5baDDhGksWzKR
YQzNNNddxJIOofByZY3M5J9Y2HD1GoKuy10wW9lTELLHJN5tUcFLbjxl/Rw6xOk6mVUJaS9OBsD+
8a0JTuPBFa6IxxE8clBDGQSObpNBqICVhk6bDalC4JTmdRcPsIp29x8jbVsUK1j3GgHWN6eMlikc
jEeeLc8y7NXO31lIrc1nYEIC4dLmSPJicu3kQbz3cRFCecC7SHvobUDL6cS3JLiHrYovs9e4gcGF
q3DUHBE4diAvX32XamlgOq+qDKSCYVWlA6yZ2iiMGjUnoYWJ0WNrmHxzr45x/YnYhb1HNdOmPIIk
vS//aQQtj0PRgpbHD9V4zpadGh06y9rNDuGpIc7p7jHN21iovzbQQ44siYr9k03gv5/dRt+OEBcY
yB8NZiAJfDJMpRAo+/TfUKqrhYDLTYQ4Pf2A/y/t2CvjTvaSZ2X1Bh+4IblErs+emL11n47kHItI
R+sy8V3yaMwWAhQ74popcV7Yy8AOIEcXGyRxcb8QM3vulCxtS7qRFxa722Ry7FpKyZFNpgmKtyY0
TpFOjapGl3swvr/BcMhYgJ2ijqbQmdDZAwBT8R16gnG8OFffH3MS5jMAYcQrAmvRJJE0TgEbuu1d
kUNyAPqRQMZa30U+O5lhFBkoTYx9FwFgDj2ZaERiNhiZTWMdrdqRZiv0MA6Mb/nq8vGrpb9Zy0p7
yZZCj1HGjLYmElkY9Dg6FbkdnOiVAXfeVh9r7ME1y7mv9O4Mu2WFLqgQ5J78+7l0lOe9oTOxNct7
jaXevD4+CGf9OWc3Nx56YR8pmtdYOfKuW2Hb596Iy44gBL6HE3p8yLN7DrbU1PI+Gq0069f6YXnq
0jEoXWN/1RkSk5FKu9+0ZvghbCehgQHX74IPxcY5IyIjXKnLMHpoJtDxqkLByiRn+mItxOw9TAkY
fXBVGrNwoFMl8cv/wrrUjRTKWV3x2lppOhWhxSrTjIRP2TJGzxGF2AfUYtmQPG3LlTXEB4plxyUK
WOXBIMbY+iXxStLpsiJLahT2CQ5VbG08dXNA2A6e1sEJ9FGbf5hd1S4ISal7nBURfok/winBFgTi
+DHoOCGgMVzL2qqfdvzw3vLQsOEXcYDzXKOYXO+EMUaj1pEXJgi9tRz7vzp6ZWJcsuLk1mXTHoNN
+y1TZey3LYo0MsrdqZVeoeCXtiE1/WJgXQNTgYx8yq6Z4Vcm1ovmaxcrcy9/dQ7Oc7Wl/c+z5mwo
avpSRbUGkrmCE2bAl5TFawj47jUZd8G/JPelkkan32vt4laBK+YMAqiUEAzB48I1xGtXcuUMqyQ8
WHg//ke+RHrl45Dq6U57a85LobPddkRdMq13oNk15LXn9Yls2yR/h/T2ZkO9b4FSWdxcH28c7a92
ejztx279Pwio5EoHU8UjSnkT72dAQsxOmDGEoj1QkxxBh0t1r50JYPr0igSR38gJpE11fpaKN0Q4
sCzSncWGR3N/TUCOIYCadwtdkLXUnHmLiNOfYGdsJpvN9K4Rutu5MbpYBCHD2x1khi5LWltc4QfP
aBoeoCd8MpvA5G0B+SyArQI9Le/x3l9fHOTinE9q2iYcF1XTxVgenylddrtgSoSiu8PvwO8bHzdZ
mhpg5MAQ2Gs0sVg3UCDTPxDcMDvUGVcvIyxm5AozP/z+xQkygcyvKg3aMyJoNokXtd0EQ21CiBS6
roxYZjZoTB7iQdXyXJlqm2atzItPG+7fi2R0Y8747V8rHABzirwHUnRrutDmftu6CdMiW1F7m8ij
yn3BroA5+regd62pVFwK52D4rrQyPHlBBTR6P6PPJvKPWpm3tWNZAw8oJZiNWZVwLys70mLMZr4c
sZCBVeGiK1Wqi5KvyMTKZ3/NeBHzii6GoGp/YkApyArulMoqzq6qyG+4tu3GIKbHD3OXDP7LciWY
SBaB9JGETmhnEZFYCmxm9e7cOyNrEISqlauDTGxvT99nlpw3a2L0jWhZ7fKbk6Zj4vnKbeW1mws1
ikKHmC1XAMeNBo8Chd8nqBdy+PhLs9JemHUbcu5KF98z8JR1wij6/Q5GivaePnlBvkouKzRy/TDX
hHSLwMHI44W+2gUjethikcLjSosK28fl5O5uaV4RdjtoZvcZUsM1C1tgdjfOPU+pnNxnFcltbgda
6CUJ3brkGx+Cqj6no0WrB9653Qg/J7f450Rz9ehWgUOsIFXJmgS21zvcXqZ27iGblOXKBrrs7ohp
XhIapiTXXrdXW2JHGUT4XOEnXM7LKhfm6Q925RN3nvxG0jnR2jNsARyVVH6G9CXV2lbtmjrelyi0
Ewrted8VW6LgwFl373Z4qO0OJAd/GjIpapLg2seNKGqomby8U8G+tvjr2rFsTuxyNP6PCsodyUxy
9aZbf6WF07UW4yiMlV3HUtr8Y6FSCkZS4bjVp8BgP/WeNxONedIcdBpsIIV3KEa28Vok4kYrKIaI
6MLfWTrp2oQsZ+SqQP6M6ZohGgg4OXAtgiFEQK0a13hqERDqR/47sp8eq2ZYMKCACwfnx227cwOI
CzDimsuK/zfIW499ahKD8BxbLqOGo4Vwz+LfaSgnmvIFv8vtoqqe8dXB9i1FZuGYvYwDiptwUzNm
Yb3XqphhQueQh2BZKgAy9kieTXh6xfnn4885LWkr22j9NeGNA6DA4xpN/1jdHLgx9y/y3MIhTa1l
34wTiZfYi+Mh5i1+3zR/WqfI6alQQq1yDu0mI01d+EdmW2xFFcoHCRsX8VD6Q8Xhc53Y/a1PBNnR
5MhRd4kZ66uGLu5BbiDqMXa0eQOrlfoAnqfr9tNn2dMqmwUUxjU2eZxeHGHhe4Mn2fN7HB8EqIBr
ytrTCjIusnHCw1XQOtBN4ziBlOM936n+zBNoPnDWQPDGTaUMBTuWriChP8/BU5PQW+0n0VQSXjrY
bhPoS6A22Lrab7yjmstkGY7vNFSO9MKkUQqioWy3Slq8AYWyurm7/xyzObUFrLkwqQOl655g17zT
O8qr2me6rjQkYkJqCBvE4eNAdrTloJ0qphO+Vvi9a5W2WYGiefxXg8kGzhv1+TSu8tGf3L6fJiyD
oY+nJxjoX4yri87tNvwh0ZMpKRfoTqc7jtcSw0YF32lYxKSAFUu/CkrGMsNuc+l163APxEKiynZh
MkDPUeGu7ZGEcR8dS80Paj7qgpNtYakaKzDoCDehC2n6TOdNQlg6vv6U5w4BeA1qPoka4w6/h8pF
oeFmC6YdlMyuW874KDyaJQqjjis5VFD06E1xgSRDF/d0DBbR4EaYqyFP/0fcH5uMLIKZgtYf//yq
vjINwx7umiFO8Ey/XB4d8DMfLNpwQYD5PAMM4G015mVNj1ezFtBS71xoti2M9Cjywxf7wPAGOexg
b/xxtLnp7XSk7fYJ8Ky7FmecziJKsyaMirbarChobWmsUbg6fFmMDWG3qT3d7rzw1p0TBmt6VsqI
uudFNnISe+noFfr86zbDb8qNgicDQWXhA0GKYzZtfAD657NBdJ4Ou1z18P+NJuLwTK/SNniU9GMt
rGgNxzVGUrOkC5Hlpb11kHRERlYNMj1V7Bl9MpG30bDNdbk0xRwdmVcDn+XYHKm3NE2ZJaIGTEAL
nkCu0GS3QxPGLha3q7QNF09pEHKbRFxSoYG5JM/iR/AZdu24zxSxvwtqerSxQbBUFJ8HoXsOlyVP
kJxdxuOzkEb/h9EOVOVo5r/rO/CFqnOAizL6gq/TQrc5hSXkbTeqm4BUimrzYX6SRix8rwjkCDjR
FrvWrdmJT2f1liVqTn+a/EZQs3Zyu0GwFGlbERG/WQ4qH2IZZJXtjdRN/Kx4PskPfAQHIT1t6z52
A1fiemK9+JrFqvpQ7aUDWiMcKDfVUNDzvvsTPwa7guTFWDKEsll9TAv5Ddv4/NIF0XsMUO3gYmcG
wj+4oiZoonCDtV1JIyTDbn7o3zWBBRsVNlPqet0zfOWSVb0YZHLmlKZa8XH7e/nL0yYs6LUa5I7Z
wAiKfn7TXS5qyD2n5jiX//N4opyQvDqdJbJXFQoi2ISP6j1CfPVM91BjVBw1p1rmlX5wpHn2DE5q
eKIUwvqLp2G1XSdqAhssFmU4/ducuHgTTBOZJOzLZDMM3CCQVElKVGt6sLpUx+oLEHT8pgPLMACo
yvhYs25gT9QjdGtvg/sEcIaMVRcUOmidCQRe0u+B21iEFfCmUVu2flkX3Vn9U8XhntySHQxHIzU1
tSbKO1HvWULRuiWlTJIQs0EEviM2+FeJH1O2O79hH/0n1zYjMNK5gXZnZdR0LMp78isKwLDjC0+5
u4oE555VM4T6CwkCgjV/wg5HzthBTKzgfoNvHae/4ol8MYD3CuXvSINJziMU0Yak4F+iNzsZJQFR
mka/7nVbiYzqOmPDkXFgFZ5fJ9vVMJvmSXlTlPcxYHkUaBFEPaRcXouo89Ydjh61vK7EIyjKNpRe
x1sN1UDgaYA8akTjKmrAlJgv4rmfLQWibKau9P5x/08UgbZgp0lwsslu7gOaCgtsPu4pNnP4dz39
JpqwK3LN2TSKBH1omQlFAyS1u9qPcQOt5nj6e+A0gyBymjGjtGBtjsg9Zi7l0pdoRYsoPGoLh2fb
vycdq76vM+lfqEWPbzHhVuZMABGVuHQqhNPjFQsLL3YeALDh+VYINnKzH2yMrnhyUiLZO4rUZ8Le
r+K5vQCJHwHn+X/ZDC2d7tzyZuGu5aCW4qDCPEDTu1oaTM1kxx/e9AdcCL2uNNMVTCgNN4WEVPOX
v/Fny9xCg3bjWxHqzU8FIixZIURF7a50DsmSjwDuRtmVfiC6mrrzAZyQ27u8xIi+dZSXOVsBTBwj
PJsUXn06xqrHWymFgiCJ1FjCe54JQMTyRJGy+YzO7h61X9BCq7EbhswgQ14PE//GRZYRXyWEdqqP
ZjI66VbSFdvrPPK4PxC/35My6Fn6EjlHya8o2sJLxWtbjQciJP1n3KQaQaJ5hGDZHn5lQMw9ficj
k9Q8UD0j3GxltZTf9ojWEUsH3pjlXoRgsoGM1PjaOyzPQvfN398AxyJ+4FRYJHpZAzDDxtBii0aW
SMWR5cz9THoPVZRUXCuyBYG0SL+fQDmYztkLodbYw7UT1Vu6kwk3S+/0U942usMUIUsk6dRGZTKP
H7drXusbaba5qySzF2hSPirqVOA24JuYclXb3etjMvkjkqTpYAAqd227t2WmVRzIbTrBeyu3Srtg
dShYZ7rCfKvYZFikcP1dmH7/dwwhKIk/R/FMSy3IRMbKtVLf25CFjBhb2WGiQfi7m/uCvi7qoXRU
bMuTYRavy9uho7l2il4jzMid7/2cPheSAGja2l7YwK/MuUQYJnIo54vqoqV5tec+kIb+L6Xl2D0q
GResyvXAH7+ICeMko0CIqMp2InX8VOVv2F4EO1mhMG9bwLFHa9cTeHXvfVaei/LqZKLI6ALeKDlA
IHFFgPJYBExOhli/hPe0S1WP7BfMBAUOegq637zUQrpHJilcdEaDlcgj2+jMFNHH294xIZ4WJdTC
TxkWNiY0uFrI8nVrVujD0s3Yjr9uAxepbCv/BfSJIHoYGEk0GDPnEu5q7IPUNxSBJBbXm3VJ696g
4qc/8ZWJb5OdIzE2O9exB3FuXtmT72jmSK7WcPOdtbsQmg6jHtVZFfmXv0fEoQuzP599uqwWebjY
DATvhpJihfMz2AFu0P8TVzERR8pRBm7ZKqMHXEsy9GWxoGWTUcu2Bobrl5ND1JZyuS6gwvZXjil1
1ECq0Yk+Dqh1l1wdB/Ud9OGzqL3uKxpDwGmldP7BfugyBJBJ/kskVlr2o0CCjDwOSVcbO1alJASC
7Xy6eHDZayY9AyoDdcD4IAWux9f/pSllaIphlNYtyujluWqzswc62LIKGGnlBPtwttRJj0+85HjB
Xkd8cKl3m6sICJTX7Zgh4f57Kz0W315oWhUq3ZrD3KURWeh1GwGR9JBDIFUBwwlZxlIvuZ5/hAup
uV2tZ+XFu0/krdOCh2nT5Jkxai6/wDV9VO2xVZUAvYKO2AUR+EeB4NI07x2msTxoMskUbhxOkRhR
sR2gxfc1wnTyADT8hsWblLnhqsEdZFsrm/Z7eW+7ZKcuxOCcTp8Q6/HceSI0Y1WaTUCzGeAQfX7C
L1be9WFtgnvAx4mW/YutnmkzJ4bMyBaF04Rk74tMzWafK8B56P9qwx6raxFe7fz1AaeBR7N8x8zc
RBwTqyCgKpU1P3UbRyLg6tmdc/SgBhJB63nYiquC/zJVKBzed+R6t8F4zeIXyZPNJcmEI9fPMWMo
2JIWnBaWAv+FgUeSLG5XSy2Ji71u3Y2MI6fb36W6jQiPYIdDPNBU00cwVjV14U4CXbHpA+eApGLH
pQNM60Dz6iznMqDVdBYzMOcL9KZMz6nSDV+1AtFyVswu5qWERGGxWc1SayZ1Yn30etJFgpy5RLTQ
lPyUBGkZb6z0UKG257bGXIfTHTPfA+XoDO0O2cFptAaO0d8nOEZnITV2X5BvkepzFaihRfO2DwIC
IEpJ+PGtGDM+jlI/XPqYvVZdq6UdMCCGM1pvSdYjgRRVr7nasrhh7VSmgsZCAGjarbyCXauksvgT
GzHWIC8irSU/3BITDnItTKYnKW96SYurvTNJn18LUlvUamczSLlF/Z6qOq/nsJ7xJC8p+dK/i1vD
bXMyIJCFfeSvcVE0QQWMcZnGeknJLYJKV8HONZOj7Ra4px6aoRHSfDPTdgA7icfyGzYRc2iRNu7o
AGIzxl0cl4FYDz8leu6TaalVjay7lLQ44kwQ7LEBPjCY4eWdhJybyuKtEMaIVWuaRS7ulwNNYg0L
vExUQXuR4yfGiJhkRuW68/fdEyFzEruHLhoz4RnpSj+EenQ1m1Gd6H1M11zUdAndMDbN5jSx+8/w
1AAKXCJEGV3tagwMaDX6+jkW4FjmvvLQAjzYVVnnzoA6nmS6NKPJ+zghDlD6Mt8onG6oUKQZhXsU
6HzAMGvD5QeGcwpws4g5YaFIXhso8eVwOhmJpArvFSLeRM66fGKrKn/vSnPFTLIVa18NFfcnbcxU
y5axbvwufsWs03V6qaIDUnLt1cnh2YaxfsKsT+JRdObEyCKu1xyxlsqpOiKTVcG6hRlajeYKc+2U
xAleGQhdsoMw1fWP7sXLqxyRPBXEEAzUNovbuEkREawoMTt6cwWE0bIa+BoY0Q9fLjSwa7H44V7K
PzGAPElCA7EIo7uz06oqkERCg+X1+sqAbZtiqOxxNSjNPuVvSWvWDNLpcLq6Ow8cw+jSfoSi+22j
A99yXvkYDVa3TI7dw2l1qHw8rji0G4SI6hlsHY/m6Msl6PYi6HQ7d7iyF6+HAlvsA+3aOSW4Q3aU
xd+rQXP6lq922b7xMODKq0osQXN41NZQT19VPXApqv6WVtN8H4AalgyoAbh6CFZ1MtbvEdNKPZIw
7y3/j+iAenq25/qHPiLu74hlQQirpRadTJnmGqbwMSRFL0CmN0u4kwxXc0VSsfnRKLa7fBzrZskb
lSgFliDYdXx2HzdtAdNg13t48zeJi5ngJWlqwV3BTDI8zckVINnzeIL5fgmI9WP9aHnwl3iDFzdv
z/QzMks96Ju0yrKiCc1arwVZGexfuNp2cECd9qcnyOYSHBOrSnm23RFM/KB7ol85r3GvDQ7d8jZz
zr19pUpItU+mQSQv0yIg2gAjp7IASjVCJNF4psCqrlsAb/GWeTJzO4JFRC35kCoUKwbQ6MO7MP0o
Qe5cvFp5CJ6H94nYW5U+z3ETS+0wJaw0XtT3q7i4BM2NDz6hGWRz/mnJU5OIseW9s/ZtBPBXcseF
UpBYssilL8v0YKNIsVi4gIP2mz6ues6KpzgYSIZyRF4qHHT2eXSU8TSpKjUcGDei1AzU9Onx0y07
/+TSOPv6cQWKEa1jNSUxwK7LpcIviqpt541rsl+yesYVeiY7hPO2h1QEfc98dh8JALWyS9X6+U0s
VanYV8M6wtHtzRVRoLR7IcLZ9Da73TkzQ49DSmY9TSn1PKbZGYCDYK6jTkyzqBjZnBbYWGECzFFx
M3z/xw55fvRoXgh/2h7XJ4kdocJi14JespjiW9x0zwbm+PnZNM/ktzqdbL0kEs9ewT/DQN5FxDlV
r+zenFBVVLw8dqLdiBcVAj8eL/8LzCickRupwhMt8/M6hBeaI/B4E72iSpXVIVPqAI34zsFSoS+s
u0X+vf34KzGbXEblm6baf5/PXGddIYaxvBuUaaAz2uI3TNFuh4PF9VEBf7jDwyChPbvX60nJvHQA
QDEljsH1igFJaHa+RnNzrhNHvGIjNG8LnO4EW7NlRTiA9D0Oqe02TWvXJU6Y11Aga0H4VzrsM+8z
RCuF+G7Y9+m3/ZFwfKHVjYqT+sGrfGzaRLZrJzXtcbDdguCbqjwmlKqsdhBy8WK97sf+y9pnOIpW
/eC7JZQUK/84/OAiuTRbqu0UPlFhA5ltPpDzlEIgbY/syV0dWLTspztyM+vayMliks/Ulci09N+w
OQ4aJSbhfUphNQqF9V9I4My7QVqOImEoxBlr/ycga3Hf/BjeajLrhwuO9vqkcNvxK0nVwttJgzHQ
9a9edL0hKSP5cL7QMcuWigAFWiOJ4FSI6tH/8nhHsDrEBFuOrhRFypToQxuhla/gGo6oGDMOpCni
/KkAoplPFd7DYICyl5my80zI0GsJYdYwC8PdEeYLcwz/l9qyWXe4/9uyFLzqqGQYCLTduXnn6LVk
YulRtqdQWskwOBayM4Ko9rU4jTkKexAdaG887hh9gQ3984LnupBYZ0wUD1/IYU/Sl6AwJ4ZZK05P
KoVipSFlJ+z6UAtHcoZynRKqeIlTuluwgpRSlvoUgj7qgt+DaMyK6KYUSKU8OVEobHLPmtb+0Cuj
h7w6a+K0QGOL7K3mz6Sqt9TAaLtP0bNbeeBnWRR6GZ7yUgJu8kUjksn+CwvRXt3rNsHgbBp8MsS3
PMLripwVDJbQWmLLR6dC4pv8Z1As3AW7PkRrPo3yUwAzDKdiGLXSysHc2AgiZ/zNQseH4yyBUwDi
StJmArBNLBTFkmnKs0cog/R0rK88SD7FHMHV5iB+CfnA7mf1DNi4GlIgrdMiv4aOPZ4MSsCC/YGG
dUuHjfc3RxIbRGttoDrYvqCAUZL8UyhhRfWvPS+m9dTjBW6YQ7Z2dC24fIjzEf6JHe8c/sj4rUXo
VtHDeHFWtWbqUcJAOuiTE9M4t+3whKR5Hk0Iz6VywFQe6B/SpF/CpUUTE1tkDtbHHuKxbYommvbd
FH5qiCi+suZXCaBRL/r6cZ3PKcbOCf7pocAhRcBDoGXcfY6NCB6+x5EkvRXHcARgxYhwEGI2gpD8
ZDg/TOxajf1wyqx5+NM8GpxBExX15ZHlfoUp4VWZeq4s4wKpW/3j9zRE0O3knewv3iyPOm0VKIMz
VLy37VQonEcqjaQKW5YJuo9jvMxDvG8vrRf5LLPjx7vhISAaLlN0giUOp+ZfBST8sp1XeguhZ3se
mdml688ZBM7yZH3UOCtgzq8FF4doYujmRh3Cyu8wziSGPbO6CaJUa9s8VQ0OiylFn+1QEmVM7W4z
/TJp+dSC/Hez0cio7H4sgSk3k36lMdiTBMGaY5DPPIQnOiw6iyNuzcwzHjm41HXi4qLA7zBmLLyr
no3bAT9VnLdowIwHG51qWRR6vQ9TLXkV21H4kyFadWHREKyV6MTQaAZz1rruAgJbv41I+x7cHq89
puNurNjzTO3IEHwoiYSZF7GucpH7kTJNcmGrMdGAjD1OoE7cVwKTJcsaxDTy3bpd++QZrhVFOhQA
RQkgeFlu+cP1z9pGcgO+ku2aGQPGkSqYBkKaMp3dJlMqOgx8PwQzkcFo4A7dCR3Rj1oANNB9LQG4
e78wMA2G2rrBed33YkDfnWktrv7VAV6NoPBPObzAGunbea/dPxLpQwvWqisT8yLjfY+AhRgz83VV
yFu+IK1q/RgwRnolhsWtlvXi2+K0kLNdTa2GXPW+KEwq/HkNfYqArkgHtnrXJya9PRCe142+tKN5
V7erVnVbGeAAcEHFM5iev7m2dD+omzK+wa8AfvcrRafJFXwaSV6McJnDLczSWu1QU3I6RkFNW/1I
2l2ca069i9afbg8X1/BxhncyI7sO0GUYwtEkqZC88ajojei1FgAYGNGoiICFpr1b2JPj0PjHDlTi
DlaS78ynrpUsWGHKUWpCRZUxvnR9Xay21pDv0P6Yuqcwyveda0ThS4UqYfgJEAs8R/lxNC3LYKtl
7JFdd8SNFvomovi8RREwSVNOfIAUWNQ9VbZVctCx9+a46TNYO1BoRBACYzZbh322Wd1W5JcSfVqN
9oJzrcGVtryCG/ehGR88ZXNflxadU1RBrxJ0BlhiBNrcaVa1tqZ/VEZ7NqxOiFzUNhU5Z5oqBVfJ
RAW+tHkCv97yciTH4oAx1VaJLd6jv/GLM/EfLCHmtv2touirR55TCzDocGORc0ZhoNw6CHb/IYhR
EN1WhSZ9XehMZlrdDZLiyoMKeotA9lvUNLDwGH4e3MY7OhlcNOaHp7BFJQlZ3CS85fQY2IwY4lAX
6xH/gQ7YCM/m59FGaD8oPoW8q7eXFyi/CrI3Xag/YNHqc36bFBcCDmBqhIziepZWHF5LqGGe5eBJ
wJD28o2KVkMAKo7ZG9Yc9DKGdHCd7JW/5V7yafxt5FaQVB3vUshSxNsBDzaxYMvjU2A/WkS+xS2z
OPSOb5f4cEWHT4C0dJ4dID9yCwBPjbH0rX6i+nY57+GWeShDoepL4TIUKNf6LOBt21LwWncVjPbf
NqRqBP6vn2rfZkbwgO9J2WlQTcfSfNX2NHZ86r0Mrv3/TYvQDFPOa+a89+rMTqxmq/Jjb6w8G45v
pX3Cv1x7UDyWRDJFoEvdcWLFLHUo7AK9eWyOx73YZ1PFvLAIUDLt6mSBIagy5bgCuCxSBAen38J+
c1cUwLW6+f1IGwFiPPrk1NTd8ABT13pB3NGYS+pQ4Gskc/C5JEqCUFBnqM6wxEk38btjKSoqWRgm
pCvibs7qHwLQR1Vsd0nDPDH/Xr2u2bQhaUsy6eXgGNFmdk7Te5dXSMdLunmtnwqCng13Os3MpM94
43XV+Az7LwhQlEzQy0xu0l5JoQPS4TwMjPUwZfj2yr3nREPNeilXYNWyCYXXYN6/uMnS9CJV9Xte
tuajU5vJoIrjnIe0xiOsShXbvpN58fCQJZX3QXNXGD5eIab+miYZv30vwcduePA4J+TPPOViJ1na
FzgavefZ04rkwVVXzoPDWnxF3OH8ZCLOEYq5Ms356UQ1MIsGg/0SXoxyY76AIurwwY9kUykNxAhn
AuiJxZJEjXpOjunbfkoVL7Py8qPtwCMzaJIci8GzcSN3HS1AKOLoj63aXe4V8tcE5XjNjTcJQImm
etadPGHSOyeSUjccizvjloYWAw+AVbfWLLR9sN7PrGjWO5Qg4iy8pQ4+OV9RWU1Sh0lrK1+0mmWo
e6nW5iog1m+OuUDBvrd83wXVbJuo2tP8RHpUHUcnl5GoTpO+1fRKpX8Bq3MsLZ6NzC+wg85qpIdh
ljTXuJkvAhzPn/cdQOxppkKonZQGTf9C8QEhmk3u0Y6Vw+t9QDB6tJoC11NgEWxhv+WTwpc8ToCW
55tuypd5AewaKD2dJmdVCj5jq1NbXfa/v1EXbjwqiFXCXzvOuJAT0qUnSArfTxlocOkC9V4gIu3K
BYWGz1nj/cuE2E81ZAgOakSKcpY/IizytA0OcEnSrSuf1yARIy/9PGvU5lU93npLaTr0FNVVs9zS
Nz/4O/1zJIhBwr1enfNu9axbp8Moqncqtjn6m41TVe3IE8ZiMKhcynaTL+d7miut8GrZY8QL89vq
0W3lrSSH76PIFKsEo1ztckbS3AKlRqwfvQhLDULq3oVQU7ilefkfsN7LBHBOWAFcxB2rw0nw9U/B
cr1YYwQ1GBR7e+jELrERBCmc8fM+LezSY5sVhiBfc0eHgjPIDU7Xjtyfnm1wh2xQPZcyShoQDiy2
quZOs3qJZROFwMYkMHZn+vowjCFi3WAvIPciuRGLW1tew8WuHo6x99j0Efg+2HgioCFExjLiNeqh
dkezD884uXEJlMke7rmHJIJ/4mg+IsUxW6sLxyq9LyhFwcl2tT+958X+yNsxR3fCxbk51ULkqKeP
/5MGsq3rlMQzbs2UJhakuPAjm2DNWJecZg36iZdY0NPcGiKrh9nwUDPMbg14JN81vA6268qSXsi7
O+d9j0WbVFs4Xy4Pz7oRLTeYhvAHINuPTRsuAChG5xdPYBfuci192X+v4ojrTY69WOEb9cdqprQO
2+GeUqbGs7Knv0CAqdGTdlFEeMBS3EvNMvRUaQg0i5aR8m+tXjbRJ3EytD0sLkFhkbva6MEpOWjt
sHuuD9LY+7EtoM47RAUGhZXQFclNqzIn4Ec5lK80Igqp8Pk6QcIftInOXJb0SEgnFsm3KMhMEUkZ
wAm2hjdGLa0FM90hjZRW9YbzPgYpkDp0bqnl3ao/w1sMhiHSJFPCCXm7XZJCTEBQPSboD6ByE5jX
V0dByLCJ9eDgjO9Ddwb2Dr5hbOmb262EBZPx7gP3I2U7qlwTYkITZurYE2DCGb2RtuRyd4T9E/Hc
5olVNF3uOdJv4OurVxvhai5JF7KdyLMHkeqeEH91X3TsBmsYXZfNh0tsDBRLAaW/wpGTC1M51Pnm
HtGhx+ViRHWkBWquyQS3ZSgf172vauLPemaXQHMUwFBxEYiSXBA2cY5mll7CGfEHw5hAY4fRMPr/
N1jE//6ey4D0WdCTDFFXEE31y5MhD62QWU9WtAnKzjcDII5NUedBfa6LT/YjmtkY+txAQ/Unr0AM
0VpegfNc4pW262qCZP3bnCYQeICPdxLe0YkDWDofu5/7eK6Kp2yifQrOD4i38zj060UzWIWjEX3/
SwqfPvThb7v2k7uuNroXINpiuSqm8PqTEKXI6iPcvvxVGZ8Ok77GhebAcQyEM50mm/Dmmno+QE7D
0neAWfpuDBYn6/U4MGVkFgle2MgkGfVukUutoVxaBpVp3rxZf5gbAvCB4VNiuLtFsqCiRbu+2x1Z
zrotIsj2tsvhN/F7oGydykFJabyy56Ms8nyquh19CqXyKoXRtK76Cn+dyxh4HypKoWTJTDZA2it2
w4AGp62s1hTh4mNwJ5sA+t5scIcMef4ng/6+sJ6IurlpA2WnGohFYmiPuCBCTwndhJ8nRIFpS95j
WKs3dsOkF5MmnidbxDbu0KbFKAzw9s205hE97PiOEihfF+rlkLm4aytlz5/EnEsjqOeCgzD1/9DR
iwDBrap8F1Gqbddra8BTtboY/gk2uEZq8tqnpoKrhEdLUrm5N79t0vEzUBiTTL9jz/39PYp0iSn5
eTzx818J5r0RIDMZFZ0E8QuUzMxMhmQIW8eRX5HlMGulkULG80hwjoJmXtU5xn3JnHeDG00Q/tvC
hROixUgNpZmhstwehA5Erl2KZYMWt+H6Zo04CkLapaKgyNXEVxcj/VahQ0Mm1zlHyceqo/IuzeVk
DfeRcczaqCTypviONUKLUjNSPyOVgIyIBW4FluOC90er8Ue3CruToIeekDeEZW7jZWpqVUt7uHfV
xZvtB7KeJWQt/xU8J8y0noSvzDd1DBR2jwiv1vMAdnDi8df0C/2HGjSl0SWb4kJeFheBk5AqsJ5i
rRNN9IZQchyfMuCl458AbigcbwjEVFotxCHklhBEaDNcXrL3XdgPnldG2pnik7PjCZUt+nW+yzSw
9LsHf//jORCdaHaG1SAAkoXNyjkkVA14BTLFPYcj8dd64ltaiAxTyPap+KaQvYcEMjNBTsJYF0SK
+TVfSXJtrv4HuoPe0rfTHz9Qblj+ANSYkVW9gEmBn8rpiw4J8dGsM9iav02snxNQWett+qB2iIiB
nXp6X0oImNPUEMRfkoOxmDXRR7tOTMW229GMtLhQBOzWNAIAYverXWHznVKb/4VNCJcCM0vHLD8X
bik90YiRg5HGQ59akSheZv+OzRzKz/1YEsifhB0SrMtGz2S2ukmurBPurvK0A7cla77ckzrGpmVf
DxbUpFnYE4LcREk5gSR/fBSw3o9OR7x6UV9D5C+T+W0st0ecnP8lXiz0/Cyr3WppKK6mT+RJk0c/
O1/1+Q2tDCGU8NlHsAwJZut1nCkmPdZ/Sug8zuqtmVBD0VYIAeVJoau2ikh9D0mq29jLBuORztQo
dFa/Lid4LCfGN/6AV/R4XOsV72qwj1mbUIqX/QS1ctrQNBCh2Oy/3FIioMzdArFysptu+HFtrNq0
bWkzMEJlEZGb7H+jKIC16SAO9U94B51UgJNiyqKCgZBGetuhCkcEuX32coo9CGTk60dWQLZSskIk
v0kiSiQPdQ4oxqwqsssVJqT1floH23sbaisjNlLaVFHUZHHvmx77ABz173B+91hXzPJ2fbFU/Cup
MUHr3sR/LeuMiLVl2Ey0w8NPtzFU7SAbrh8fpwqg+7Ihyrn4TmLn3TVSjLKvWJk9K+zO0HZHB6q1
VWT+/WoNTWTY8D8oi+std7LqQ1R73KFRTtUEYPeo74YHn6SdFjbCRQSBtQWxSRtf7bnrCiog/0ke
QLGSyaUPn2bwBKO4spGVKtUCpFisLRApc3Gb7oPvn6Re7evKn2gTUh/nXak9kLNhw9/Ptl9bCqSz
hQkwO80Y6aW5OxldYEcSdGw7vloWBTD4FwcGh401jgTu1SXoqlLCFts+ztnZ4ocFkfWTNbmKPtjv
0Nb4hLqY/5UT3/VnxlOO+zR6VSrprBVEkOVxhmookQuIHnE+hxfb0CgBU/hBzPhomlWXAkHKbpDl
8hyEUywffsZKgh0S9PpnvCmwcg5YQ0X7H1+C0TehknazTc9TybuGlNnGn0NSV20Xj9RZNqWi97Iu
hoVXecHNhDSGv6rTS5qKJIU3vxcyw0bnPUECIyS8X8FMrKif37l/Fsi0ZW3SQwJyUt+8FHj8PSa1
xG71MRLdH3BmX+WRkyQn1GrHOdSmpxgc1zMRAQS+5AIcRDgL6KuF64057LpZazhp3Lj5t3exN85W
KwcEflaT+FWBjXLjwjzSTU7xN5dROipTH4dYg3bItUpBT18QSY71Lgl0v6Fj5JnL8o6HKZ1hGKMw
qDSJuCXCSq+r70WlLo8+pz0TOQRND8A0A9HaoaW97gcWHUhn1mvXiGcUTu7OqTXSwwfxQUdbVNwK
zAbLkq6/FxYvZ9myyBELgkGpI5a+qQEQzIBm9eRqnB9WBs8cXVQ2KkNqlNdYm1YZXfEBB26q6kv+
DEeHqFrmcntIEN30XgxWwfjlTNKeSTQLXs5jQjsYYQVo5lGh1bBxJnxKBgPea22AH7KkwrvuiHIr
ckvfnVfAFvFAeZkrOvmkcWEEpVqpJWwDDUNynVE+nWfvZXLwALP0XWlWCxZF+ThjHLvQBoaEXKBm
BoTSS6nihklHbnmvqYcVomEbvBLYx6Nzcqf7e1k/8ltvEqNGjQrqbEhfgNevCu9MdX2q4qR1COI9
rWBDd4uSFAiCRTmoq0VPSkQa4Iz4qSFxSt86RYqQXxvEGGNctIoIbYBKOoyJkCB66tYQ/aLe+D8t
aD2yK1m/1gdoRjLPpvShffMwbAvPMBKBOyINqbkRlt6FbenYmWkr6QnYMc7QKxjjMFv67se33qxb
WuFTMRxvPIQNchFVre5JzTirQdMoDZn2qIRYh8aBOrnsu69bmu9rFMECNRI/qdkxwAkMGOuPxLgl
sdGLUrLWkkTxEb7eRQJYrkGdoYbdcVthKt0EOwhGZCPjiYQbc+ROxvu/ohUERN6ojwRilfNluYiV
wD2wPb4+kZ90Z5PkLVxajyKH1eQWO3GVDwSHM/Dg9N0qejaft9/1F7EBOdQXeSo4l5hmL/f5oxb7
RaTsI9C/dqNY96SX9GXEIXpPOljewF0dlTbyjiEsGSRhO0kHN2MC/y5a5/v3ObT5gETOI7/hXNRv
ziGSPeH4x0RsTVh/gQFG1MBFWepL1UY0jEwUJXpVqB0W7tF/LwwAq+wuMMJEF38pLItffHHNK3st
LH7GVbSwuw89il2GvXQDuRIirrCbgcbtpQaEC1uRTe+mS/XI2HNjnzzX5dYzRT4Wxq6Jq//m/+EG
L4cRbkX2enApKMy9YvSypAgZYRv1WxFfSiiODwvpJ3qyG+JewdxgMbEI3flaAI9g678/yB7GaIGL
cJhBq8PINvjv3feT9fa6Q84ycyZQ6iW5/cVtgEf+Ic+dA7r3C5ULSmyD+SoLjbZBQcrp9qu/hwXr
NJ23moPleN0fm6XcSSuSo7O+3i9SqXyYry5JAnQIdcX78G1g9CooGyhRu+CrJP88ygRrLFf+EFF8
hi9H2PY5hxRmADSLZIhFc9OOLBRfJQ/JoYzAT3pbz/KSmFfHMv+oUPkXTx4zesCWQFkR1kvNmYZE
drDrlW+cS0Lp/jsUy6ObY2OEXSbomtFURKqm5syvdDKB8kaCq7v0MfAHbsoFukDiE2t68yZo/3Eq
86xHvYxHdJBUmzXSkyv7p9j2u8G5RMkH+euHXe8ZjRvAnW9KQRxHCIrp+b4nkn6vHJ+su5nUaZsC
xeO2x7JWdziFO5VHsClrPHQ//nkyNWnPmNwf4shKaVzsIuBX3hd0l2FcfKIm+K7zSiv0zDfMpZmO
FSY9AbAd/PYprihwYP1ZcHgPlJT8DG7i1vEOgzJOGrblllMclHwTacFjjA0Vv4hYEpY7LUVUXFYe
D7/DejcPo0+V9/GokEdZdrkoWL4sQRBV1mDPCfmbpGXUrn9gBwaESWvVr1luIRQjC8zpR/JolcV4
85KUVd8JI5CK/pWDnhMmP46gKSul9gY5MDhqTSzsf+SBqjncoBGgVwOKydg31nirjNw/XzBgVmJx
jnA+fGFxz35sxc7H1EFhyGQPKIg8uZkLZEpvolM+jljWksqdKeE62DJTJadrkMX7Zc/kJx/jhD6H
yeNqXVlb3e1MJS0d3um74ADpDsUdRsguoTc2PHghwCaiwMGgWvr7y5G+Tn4DF1QZ4ZrTznyvUmnF
jE0VNoIkJ0KzkhHvvCXHYnNJmCoYG1EjG4CcyRsYgnFU+Juh5J3lF9fN+r+T3DTKbCwfEcSanO3q
w6ZEuthsPZD/wEk8IAJTb2R16cO00cl5E4sLl7XUkS3iu58EiQPTlFDhR4g1wkl3q5NHOGh3WUDp
lM6r1DbtJjH4NQoljf4pnkkCsKdomQfYqfBoQ7u1O2s0uBYz+H/uUXIJ69rYVfjFkSBb7F0QdjqT
IpyZF9HZkOQV8GDbfIR8/nx28TwoFUZoU8agsb5RDBL2jJ1dQ9c+vs04sGpsCTcgCAT2e2Sf+5ET
EH+a/8RwcZ67AKo/PcrF3FkTGI9KiwFFLmu+zql65N+BUZEF7DECX3BerDwXooLWNgT3K3esdutc
sTlITBF7+Dem2pVRxZYjZjGFQuEIe+v3H5Upk6pSn4oNGllQiNt3KB9Lxbzq0tHLCQ6Hx981Nsr2
CdS9noioQs5XTW8u64MXSvnv/nAAPP4TRoK28774gcFs1kthv2kRKdDLXorSk2Kz4S6L/c+Rvdmx
JT4qEmUyHYf0lLMGUbPsjMCleg0b5XPTtShQaTfwTtCXgc0DNFkLUOmMV1q0g5Mu3cnwzcb1w2GH
L8T6xhC1VCggbqEuSeFEJeI+cFDVmP0wKT/M9ivWXR6+AhRr3IY14tGI6Cc0RxOgvsS5AJzRovmb
73eSoB6AAbcNENQwOn40yRjRqWJ8ukIyJAZgue8dArH1bJY/hkyeyNdaoaczHfTjdJ6+DqsKbRfe
vqgB2VnqHwF8SaUUzOCn4glaGVMRBdHZ39g1ybB3OjRy0PkGHoHf8PrOk3lzLnFf8ZCkqCWIAcKX
T84vLaFOm3/qzbF1RRhE7H5nIzX++VMteVPXhc3tElN1ZmgCulwO3hLKtQLzt+4XB4tgdQZk9Nbv
XpjNcHkZ402GzGHAxnVtoknT68WfWHYS0WpBRjT/K9Er1P5N0hC/oFyHWBXJu2eKs/zmTLoF45j9
5VeRuiYCVNZiuViZO4FYlxDmLyiIyjQFFdCy1ZyaUk2ggT++cx3vlXX6k3mihiglZxVOPwnKX446
eykc4+CbxvEL6SXjaoG1JVO5xdSVWekcR+/pp2W3dP/f/l4ocyJZU69hVms063MgD08LVStt9Eyd
zYKa7H6bwjyq9kVJys5MSrxNbQmp8A79ACcRzPp/7tFZCuK3w9iqAxM/iar8/nyndBIAgFgW+BMC
T8JqZLrjOQMD+PIS3q//BgjYLdvLSKCTLrPGwx85Pcrn6qT0NPipaDWUbxACR1SzuReUMWrsS9SR
k1B1GOC1x2z6ypln6+uaUOJNw2BNBw37FPc9AcpNy9z3+A6w1Y9dOaakwWZVwxyil8bwK7gWdImu
hnIHp2J52zrPqemxU0a841Vj9L6qCAF74OvU8Glp+DPa3k5rNKoyoLwUyJtoVzCOpQYmEPRwEIBG
Hsw20kjZN9TUzOwnFy0lwpFQ/oNLtVYBH12lZWLDSVdQZ99LMWv7uzLPTHuTE3V5rvP0jUjkFZEL
EU/x6EpMw3vYk3nZmDslHP3G6AwbPOO50cDAufeAdOSqImD4ObOTwmrXsQhfisx/rvqXPetnzrTf
JT5Si2bvWrupcWIuS0EPupaA123qTv6lbag+IZ0fjwCuW3lwUlz6R3KXkw5/kL8epxEJCeLF/g54
4Yk8l/EZE3LUtuNHGk6l41xI5Y69uQP4RRY93ELpE2P1G8IXrhYAcFmtdXdWSmHvYcblU7JYf5wZ
lTqch+1GMMXrY5Gw9owSwIKe9XzUDNDf5xCFeUYzGDglSjjRMUUp+iDuhFhHPk/Krq5/U8egoIWd
gYv2S3cAwbDHSq5m7I/PZd9+PgHj2MINsDGMz8ta8MG4JAiav3pU+dhL7Z5rpro8u78I2Q4ulYnl
pSHAYrygvgGvRYhqvKmK/fV8WjJM/7qLQjtHYiXjMn0FfbWKZl/5S2yxyCCW3ZKA0GUApPdEL3KM
wviAXNWqHfpAGKkPxIy7TizBy+9Qi/y3xdZ4mRGamZyg1Sb5Bs5rjaHaGSKvGPM+k8mnRkP7sifj
7EtzcoUthe7MUrb02YfAtVcdfek9pavniHCIZzmuOnFO/h2FNv0JjAPsROHi5fGPa1gIpApSQxzD
MoUh++2kovjtCegBgtBE0DPK0Hw5AQ9ym1bkXR+0R6P1HBdkrUSERZl5jXPnPuDxRo5G0P+ngOA+
riP2SG6Yskhy95HI6YIpxidmvwWSEI5uc7I+yYC3VNxuuWsgNw7YfKrvZJX2yPDQ+f+hs2Mfynn4
FWhMnRCJjRR+MeT5n5jxTgMdXRvz2ciKBmNxqA8sZwJc8Lqenlrx9sAzrJbk99f4p6SvJOZv0Kql
axNVbiLr1pxDGEizLg75I8bG+1iUjSVkbWqCC5oxSaCcNoF6D8hrc6qGsWvzyNf3G01K1LFaM/HD
scDzQeuRfqSZSsJjLzwEA1SmkYYDcTFyzPok/Pdc0IyxRW64gUhe2t7rW6BeQtp0ppNEG2UL0g8X
piegbrIaUV3eeN9p3pMdmCAIdyWghYhBDjITx1a1zuoi7v7nrCpUoC/f4MW811LVJaYjKnbtRBlC
N08UhRU0E50d4jbttNZrKQ0G6iVZqAOMVhQzrNmY/6tjaiUwmIG2SsuO6vJBlxbxx4rG06IU54ym
jvTVg3VS5jnqk8RtdW5/RnghjadQFvJCIA7DMaZ6w4poyHRxYhWjmmTgsBLcJyNnvd47YsdkdP+n
/Qt18G1Ox8sOTyMC7CRiV8KScsQywPV6v1SYAyEOOKQNshmK0aEYskLcVjmaZNdwqKMHiqFSIrJQ
w7rtVPN9+d7XAakM0XFF41u7L/CMbEYPPrg6FM6ZwOjHORiCr/Vp+dV1W9inRCZTzp6nZhBFZvR0
1lT1jBVJ8uDbRJ9NMDh2Q/YIf5nF+BJ271Avp/w9/hFhHOgU7XUn8i8wXa6P23QjewSdrKfvered
/FvGVpzmDTmPCxrL9hna2VHFI630wfxuRc9CXsa1hBHmMg3usrr+7ab0Rw6p92mtEub8FI4jh4Pb
gnIoXgNKgplNP5PHQBfP1gqgBxWh9glKNNzBAtGFN3CNdz4OD/PNC+pBf3xLj7TC7peJerdNqox0
5rq6oTKv3LWMVkzHQ0fzi2b2epEuNm/b890Zml8/LnKM73ononqfk48vU84FoTN8x2taaVEA9DpG
SZ5JRGKHosA/MO8lh5uVRVjAHNEuYKu+TIZTH0f+FOg8+D1rWGFcWG7kJhFgmYZ6CSoOzPspagsC
dl3rDyUakxSiIfAJ87/G/Z+YyvWajzzhfxy0j4gPP8GR5fwAkDGDHWjGm7dM3b0v8O+By1HrOgK2
FaaeCbbi176MF+BH4COakqFvzI2z37qMw1BFb1nD414KVUjb5rcGi3YsUb66+SCUNqhXOZA1fkRV
fOsKua6D9/OB3k0Yut0siFKSQHjBQu8YseLdoR0gECr/lc93xgbIAlD6Ut/hOna7eTqPRJOtGzJX
0LbsJNcQ9p8kAYwqSXE2Snon/2/+uG8LrAU+6CFmadPvXlSWJUFX8iTb9XfHfp8dt9jLhwKpS4m9
38Sn2QQpeYgEKN5YL71E5iSdLEWNt75pMS2TeiYWZMlRfIgcQdhAamK8rOt1HQch+frRPDcbtZC8
lmL/b5XDvg7rEWY/V6UMoSnReInGxmSe8SKs6uf6mNUQBYkcRhScpmQKpymBUaemCu0EDmcHlZyA
sS++fm0oe4pVEOHRRLjwppFG2PmMn76vzjbWMTcGtdVO+ezZ0Pfaq8kHaMdzWRc3HViJAzGemhpJ
KEOkkcNkVYbIEjPPWVTIogTM1n06hpeNMl2SG0I/pCeuUz3bhfB4u8ddkTWc2y/q0KHQBzCnbCD+
9o1MdU0kzdjquXWWi0bYJJI/Bg2nzwsRDWLYreZ8cMXO/M1gBWSW/lodsa7fc1d9vuRFK4ZcPj+R
csuBmAivUGqz+9vKExD5Oo80G1MiwANtn1LCct69ZqcJgPW/F+FREPijQ6ipkRXqPSm3MIBkkPSw
Xp44c3C99E3phBhYFgz+QZiEqjnE9mvIGIOO3Qc4pQurWAeO8I6N6hpmHOnFFyDItQg6/C1A7mVo
ciuqbkhBt3MGwj6wtLWLBkcwQ7edKjSvaT1z5e+FqX5uhjqQ4tRoxAVAtH09WdfKUfZZkLJX/Lvh
+fNUlG3OOO0FAi5UMXc2XFz+Bhv/kQ5in5SoKWXbHdqITHQkK1FUMElcEhwYhrWXyHlfJY1G2a1j
TPtRdn2TbRHQF5hOm3xBTR0pWghvjoIXVEqCXf2tArWL/Af30W5pVg9zQVcjGcS+DlHOXWQfQxn4
Pud9DSl4cZ1Y553tksR8pG8WKHUZHfj4h+QA/bMuKhofbNWw04dAxAi1GMGA6dIbZe5UhfsAcCUr
toHlL0Glu5hg40jZwzmpWSQjuQGVqoCD7x5HqWbAFkKUroi7Konn9EKxggse6aOo5Dqsv290tLet
su2PCwXQEllc1p+cZ41UMsRRvGdisF2+tPKEVfpD8AdDQ6+U+2HXEpmBJZNlNQwKxwyP7EGVtXyJ
/UQ5ZswRlUQAalxxGBC9YVFlYmYNzNT2SGpg9X+vFzOhjq9RgZfTNKo7uqRua3m+JeDb2x0yein0
Y/+oXueDJL4FyP01oq+a3W803hX5+1kSLldpxnrMVS3tlc5rd9fqJxW/vy7zil2CqS8vh1gsW653
t7LrTyrz0vYF0a4CINKg0Fugc7WgKeL/ygpy3nsdq/EjWsqMUbcH3fxiTHRMwA8JiWMgO4nCPs+0
oCNyfQMuKeithx5wIOlaitzgY1XpdK35k5Mfkp2+2h/MycVy4iK14HMjY1D7G3BXOOSkblmRW4DX
X3f0H/CXPWe5/rtjnlihEO3l7aFOEe0Aunfie6PuMFwoKedvYS9f8x07VX9RItpZTfmbvSCvtMrA
kVqwmp5ZonjPzfzqZf2RFKtw3owxS8kAm4SXOzXTYENZ0gF2WSB14RN/JT6pnKrcrQSh4UjEWyGT
Fxq5WH1E96QV133IqmdMchMA4uDoiJ/kI8VJRT+Wg1HSEWN3ri2VAvio1rsVM/C79B7ngA4SmYNB
jy7RkpXbE/jrRrIhLwtYU8kA7UBdSJOl/C4RpJMH4me48cKfP+co6322WhhtIfoY/g0Lmz3eMpDR
jlIYL10BZr63uonWOU2SSn5uT75B+in2h7Amai5TeOKTK4uy+LWLwrXGyDDnIIPMb2jdnY1Yv4h0
i9d0slQd2Eg3LSaN8BMJ+8OmlDIzL+hYZ3I+aZLCuSHJt5pwvymc3GiCyTZyRTpkLyrGPzR0B+DU
6ongPmofFaKvaNRuEEs2EAOTySC+tTG1/UdvZ2JgWUIOzgdtb0vwPq1UA5GBgVPqg6IDYn00bCDE
S8jGfh/Jv3Ngc8fawT9FA2+ItWaEflFciSurp9Ic3LN0aXPPDbOb6k+fMOxSlizl357yBDZITQpK
qRjctFC+e29A6VDZX/wIRf8DkZM2Tcb0w3abE1btiTOalBC9+fgbkgIBAJ1ulX4Uc+fwuhvC4blk
BHKjTNoVD74Y/o1aBI8y8rCC5cYDb4qXQEmodR46FiUazFltZrQXP+M07cHBePzRN/p9/1vWIQIk
QYrjgDF5M6Q27NDM/nP8sCYJl/IJ/w9wrpsqTFLczr6hxWcMSzzwesuSJ0ERo+Zi+xHk9p/uD16M
YGjizJeS04/9uJ29H51f2lbB4bMaVzR5cyFXyIPALbwe1k9ILrVJsUmskMWhLdDvPTZSvOnXj2Zq
mAlUUcP6e8RAGFer2NeogCpny7EF4dKy1+PMmlQzOIQuvH1kBoXDURqT1gMVjNG9BS1ytDcAsB+f
7Nt7ifbkNWJ35zUJKtOxfVnEthXULqQc0VX+kpcpACk3DE0Hwzbfuje55OycDnJWoePT+HBwa5ip
4ma9fEd6syxgZQnRJnWN4OivvPxnX6MuM7EG4ahKdgu3dQ+Wvlpt6xQjPwiToKPb0KkA063l9FRd
9U10fGzYE4jC46c5JxYCVapPxet0ipox/TrctSTrikwLQpJmrcLeYCBhH1RT9rwnMOZQdm33i6Qg
2ULJcwet4wmi8RYwVIGcHaMeBhWJbZ5/3ZyJq9QYhbBu99QqJnu6V22a9mkk6mnoYnS5UlLYeT/j
G5nzHjOu+IWkno6gfxLRDvMeC3VSwOT2mTY3bVl4SKyzejaund10t1SRmHkK5ckoYiSTp9Lras/1
lVD+WsvYdrcJww9N0FjADmoLqITrWFwObgoQ6vxwU6fD44W+s0QR2eDJPkgZfynTuKvKDqiaopLP
cPJPyRfeE5NfTYEVYSTIXZPv3v/Z+GizGUsHQSWBQjLk9KsNYOP29xAwghZ2tUOFb7UE/9RcRNPT
tg8K2qVhFz5Wo9b5uJoBGtkj2HTwviPFGFc5tt/fuG/hvCxpYTXzJWrmrktHucoaWaIgwdq7pS3S
FACGsX1y9kouQGNWKNtLdw7aBOBZ0gI9p16ARco2RFUo27q1ZmsoL/tllNgahZQxkPoYMyPhfp0Q
ao5rBy/Uv3V636UJ835loB7iA1iTbbxXevQGBdCd4sSqHcIAf6g8m2FeayJEG438qAeH3fuJVOdb
RnpZf1ib1jWftVD56GGd4x2ivPEYsaYbIRciD2EqPPKHTK/ysyjOTRff6fPocidXXKWs+GAxPbC8
yMkDUg7bTZl4yLRCPsBjAmVj6jtDa8/39/dTv/zruhP6mFzENKif6TnkyQVFq96J/Iwe8aLx17gE
mNtZNxRZ1ZVQtExmYrbkOB6DKtVTPbsaQ1BYlx8tQwWygbYP5RUXW25eda1g4V/nPAJpadyVJZGf
WkT8CnJvLJWO7Y2R67BU1yPv0mzaTmmb4nuvbyZtTumDiJi5rFGi2Hb82pWd8BOOHyrSt5vAObeO
rhBcI4ZJl6PMiS0klcyeBv4Ql1QQvTLEU2bK4LbUbuyHK0/FBeOkloV3+QKZpKFP0m+sG7L9O0va
+SWJ/9FwlPgj6Seqkhz3WwrS3EGB3LQiiBLuM67wmrjzypbXBvWpqSZlvuRJ5OiMR014o/WMuNby
YsG7UWJc6/ecUeZySGoZn63DkJVHhwwd3KbyIvAGXPemxCVNBh8lSFmAlWFSkDI+M1II34L7xpo4
Ft5ix43HQmmQeaomsjJy/zZCgwgNCFALpinOjvQlfNBkNRpsjD6AQcQ6BQ/R1Na7Hv3d9OOklF55
Ok2AaNL1KYVKUnQzTo2KiQuK5CVBa0J8da23hJpztKWy+o1q+CJq/K/F4TkEZYpgdnHDWLMiGN9+
ASta21Q2bX//JHYZGtGZeuJbC0IOU3GzdG6jQR/+UcLJk+920ybA+mSgg7TH017wh4oqv/KCw1Ns
ipuai/6V1ymfKc9R+IZxcFolbejpQO524EEETsbkxeCPNQuNVYeZph2Kzl6L958D2CqHwXE5hiPm
J2eI1gr5JeYHYx0S9kdLZiloHTdYGrmbbABWz1jt2jbpQbNQ1/2QfLd2hULwHoJDu/iVcmnWDUc1
X6sCiL41+UrtzBNbr/T/fL20QaVNvv36iyJJ90a3lT3vg/QVf80T52ylx2n5OkaHmBDzaoRvFbrm
a27db2DG1S1T0y8O9lbv+9det2qOACoj2Tx/9HCylmkECJZ9S72GGQX21avfIALzgfhrYI+niMja
5DLZQdjujvIBpVO+sCnrcZKK4vjNtlCSORFfmj0WtreJkoL7D2furM8MP5VsojyoXBg8ByNn6/62
/E04r6lAZoOvtlPA4p6CExN9F+NCMe1LPxn3M9iO8KCVBhUlJmtyGRfNVucTBWWumnA8FE1XiHFr
N41iyHbMPGmIUgYMoqj6abZOoVuwYinu0BXlFyqjUe0tOkwkixjeoJtiv3ekf5YMB4b6icsgxsAa
e4TlRG+cQ4SaxTIWR0Whv6vtkXDR7kEOx8AK/HrIXIBWeZksj9vmWdqqq1cxBtah8UafkDZRvRI3
97PUtNadNs4hc+zd0UvcOEa2/YpFtniDH1G4XJWrzeUMjgHqRa/1P8+H5PW03PVlmas2x456RJLh
3srdrpli1oLyfowRTfmZvTBdBjWCZZYBnULA7bH/UkJIx0mjtil0ETtX8zvwbeqaYdQ32uHPbOQK
AiSGoq/qcKprdIn1bkRUeLBpuDbqYDsdah88fNbt2tATeKYTj5vcF3YNQFOU2z7MDbhuKir/oMX2
ln+EVandX6gt15a08YnYbPtPvM0XY43MpfhdelnI4EfFLXwa8WiaRf5J5Ico366G+9JZ7lR2EP6u
LA39blmRK4mpvmCZEOPOOhExc375Bp6S6UGaobP2of1zTKNmQwjNRnUBo6Xre0u4ansWqObCcaue
kU7e9qljKCVs15ob3YWFzx7m7EcZYhiE+owUhGw6a08ZGGw8rJ0U2AuZFwPBIN2htBq64RMpMN0I
ibeC9hDzvguMe1PESev26lriS7hdelyKVWyA05Y8sPKomUSjwN9JgWsmD9T6rUOL5YKpNAOj0OYl
8Z9ZCNOzcZ8Y+nIknd4iIWMWDmYzQyfXJ7VzgPq7BKzeBkjW74bubVdO1FGDdEavnMxWeph00/TA
72sQuIC+UbmQOcKmiux5y1LCyrPbEg7VGI6rj5FwK9EefdYe3oo3WDsYBiTrYvnZxJ5gBgF9fDSo
OJ/WToW+QnIdNAd9ZCa1eNI1G5eMmsD415iqznygtd57iQeIbY4IR6R+QVhPfCk2hWgvHx4gxYjp
+YNJGO8spE6g1FS6LsdWD80Xxjb80VTyfZ4WdmoY4EmYlgPdqJnOnGXnizmG+WXvk2CldZohM0Q9
bjp4yQx/alwppMEXQFhW+YkC63B8P0+X2Q3DVWuefNUWGIpSnWKS5L7HAB+KSF/549prXSncBpeZ
/qBMLW4Jg2BdaRr9vKHk95JuDz7LSB4YLoqVQFKCDps+0Xu1VlOfXAvc5MGCd1zcvXtfdAg1+LgM
pnQHYc2rB9dXdo9XrcsBj5rmpAiLpOys3uocYHm4/rbwoLy3pXW3eH45eLYp3zFM3zdkhw5ccUm+
nmyyJhdlrnLugZEo+5/AjaPM/hCcByqyDNpmEeBZd0ITAlnvlneI6hJDG0g//Kil8Iuwv6ZoaLeF
ZCDVsktu3xPMsK1R/JKj/E/CSywbhkKhuqAvsRZ9USe8VrprrH58in149/HHCcp/RjmFRvWRCTEe
cxthO/OQAmTfcspctQCHEBwrLL+QmjGuTCmkMeYXVp/wsJOxLZ9uYFLPzBqQbJ3V48szZXNeTfsM
eOIh4ALBpPIjU8Nps32DOzGiKdKd9nTPTggtVNxptCUMuWERhXbhjzoR1hwQestzbCKtHKYecbx8
b/CJD7+6g+g6+pp3Oiwpp4nDK4uta0htSTHTnT0oP+Zs5luQpAakFUdqU8zgr7U3VdlYUCyO0xuS
4/R3vc43m5+5x7cT/ab9XqBfJLrrd+7XSG+tNCU9jieCqXEuHRH6RkIqkCg9RIylnOouV3oRrtO+
IERkjkEWtYNF+QpnccQXRGph11XXaruKsD0uoAFNbW8RI3PhqpWiS8zOweuvEZ/HNnJGMhfk7TZT
MvS9RHYizqyTdy7GGiMhv8HEHGcYU3uBnQu/Cd7HFgjvFmsoZAZRDJEI8Nno/rxK4Wegn/ri0//T
rNqul59ny/AvebsptZ/Z45bR41fnZv2o3iOu1rPcQIqAsiMmPT315gI0ONgf+ydX8x+jFSVb73/j
jxuUvky7JdKgR6bN4rm2xrUtY5KCEDakkl44WBs5Ks3cIT5av+dk4AuJqu4x3tca3+3pKBY2fzqo
sP9rxBUkiBuF4rDa0d37BeI7uKYKq92I0gwzyTn5srH4UoCmW7jzMJ3116Pqnw6Nb5ZQIUPvyp8D
mo6bkV7I8ygXb41njGxnFyznlIv0w0CCU2LnazjzXtg+dJ0WH1jDaUGj3VscSfmQb0YI14+Y5GJK
kUnTwSA9cxdF0O/tkm1d/YsagXsUw2uCyNalzUMsVJ+prdtTbwUJh2MUYSLdr5sONFbQ0dZhdNjP
VKNawQAKnPBe/07C+USfm6jZJywVMt4Lkp1zaPGkpqBVhMOHzm2L3BR/LSc094Hx2TonCRHTLXLp
gb1ylwJ1cSfeyT9HqkVgyiqCuPPbXAOTLuOhs+SuRfZ6DqCNiKcnid3febwMyKmf+y/p5qktBUcE
3NMchIo8cqmsfDMsjdXzQLn7LnO1GA3JEZbiCWeNx1r8bETO/UX4Xyj90BYUUIV06w8jR+JBMGAm
5b6NjdY+q5mn5fp/WnqeCP/JEMPgbJNdqsRSDHwxKAMsXvuyanqP7kSm+mgHvzbPYmUCZSwtCklA
VqeA8scpsd3eUBfWE9BCPmU5KnBwKjQCgIiry3qX/V1qS+M8og+WaO9zoIKaVoaoFa8pbL5gtg1A
D4nRUPY/qQ5HePejUPzjtzqHHL9tmpjqTu6aPs/4KbiWc18h6to0bdqHppppywwg7o7iDxDJEBz0
hyJtAL4gMeydw8/SO85ozShG+beGGnH+kYdogXtXshJskLqnvQcUvHoDQv36y8rdHozxPAQ41bH3
h1J0COL1DOneHw/bmMwTXqb/MV9b2pOyVwXFT6faWYlaMR1G18w4WnxL8TCBqV3ywy+RM9uuqHxR
5DpKbQTjGr12OPbNzmC/qRwvMwMqq9IvDHbl7veLskUD6YYVGLQ6GePX3Z7mteoK37+kppRIHgWv
QCjDNuuwWvS0dMH64QF6X5VTsI8619B2exDZ7nqKnrlbSWr4UNT66imAW5lL8K2whS25+xICA7O/
kERi4leF8LatbMW7bP+Jw/Xb7dNsQRkXk9ktKCB+xf/NJYoCaOUfNjVNvsrgFsAdPDFIksV82H5w
aUGtZ8dvH0P/EDvMwsR7o0P0yIcICXnAexbO0Y+KEKX0ReFW0a60WpvqYrHtzj/H/XvUyGR4e3Sj
/MOyR3rPtzmQcqiz3YaqsAeTY5Ez3ErpywnKcabHMh38DcpQHsRJh7EZYxpZDTiVpRtlDYcbmgPu
q4sAJfpmcQ7H7v+BCnzKmtaVxGzJ88yHqb13Fsu+sxbvvfNsfy5y8ehbmlH+HVZ9seGiZo4J4xd6
dVJb2cQHytOECnZKDjxE/2p6ZIIfrwCvjDLP6XMGSSE3T5MoGa6v9u9FVTNoMf9UbDPz/cQh/xYH
zuN5u2gMAy4IX87BEFqaVktOE3HJ4jGdfhqj78cTW70y6/g5BjOj4QXKmTu7YdV5YXhVhyth8PVV
3A4u23764HQCWe8LouSyXKU/9vh+qsbr5wnx0hjmZvIKAl46hOE1SYXxCLQa23z/l/Nr8+hYa83o
QaOI61Yul40WMhBhPsXs1aU6xlTwuY49DMoTpubXv5F7cybvkA3ALGZaRRWc1vC0qmE+yagEolQL
yhn+9uXl/jpwkgxhUFP8lRil7VfrMEuQbNgD5Aw1MtXph/X0Vnqj8cBENkJi/81n4qNRW+l2QXQJ
l2lwiDodirgQa5cg0wJ5UraRBpsu606jGL/Q6Ox04/JRVTZQi+9TUwBWWaNJE9iZ7czLKaWbY73H
MIHSF/4MNWc0ouhbceieo4Zhypf+pYG8Sg6mFaMH5tHcfY1gZTnNLNo7rHaiuUR9GiWP19VXYYc6
maOkWlrKebAH/Xyb8vuXblmZNOEdL8A0fBwUmZsvj3a5WUKmiOgPZsva4dYBMNjImo3OA6Gp4YDk
lhmhLtGMzLQowautqR4K8YHraUJDhP7Ap1OmQfc/sJe8AuD13AnjhPZP0qZk5l6KLlqAYsBRvqoV
kwExGmQecHNp8GQ9BgVxSH2KOTeB4EJS49lmE0xjcvQbRLqAvLga3oD512fEfxpyP3pn5rBy8Yur
SBrcLgAjrlHZh4VHf4sNaFQW3VdsQzWmj2lseoq67cbLae8rBAZnDn54+/yqreR8FshR9dT/Q6th
T+5lxWOScbMZ5pgPKAHsG4KMuFkauZoHNm1Yy96OzAUvCVGvmhKfSTonc826WNVt/TKfAVRZQCHZ
+bwblkGst4QyA5THHh67j2jlLTEaE6ujI+qi/pi+8M9/m861r7AUbkxZgzAuwDVcQ72sJ9h2qVMC
22r1Ur2jTUyLRnAfw58v80YUjisved1vXZybN1wN2dJREBfohWPf4v0qnTshGVwFapeDZXKW5fIz
7cKU8PeescusO42nMv2WPnA2gsul5mKpVtbmIANLJ99y+F5U2JKEaWilEgoVFqYUv0xX6iEOVXRZ
AZvheqJ1x/PJ5QRDSs+wJ5goF2kXMTdGxoFBeAs5YNhK/uFtK7qMmouhxiwAkVqG0aQVzdFU6Lf9
TWsODiywLUp+uQNVNhKfsKZrGP27t+QS5jo2e0nsk+1GFpJYHpcOsVrLusV1r0cr/0SAw/oi3bjW
59WiTtBJY7QRfZXCvlGjaUD6fy1XXQKtZcneLGo+CyNESh+gXvYeKD95UZ8iKP0wIlrHjaDa/Fhf
86chGhVmlCHixdyz0xlYiFjOf1t8Xbt5AcIMN8H/N+yYQGV/65OhgjAPvbqvw7pgJoaKW4rAI7+P
+zc2GVhcj6bNNQ9MhHTkBbJF8+hXPC7lCvyQ7lVb2MeoDQCzMMHIe+ECi4PcCincobNIVeE+S5+s
YSmlHpvcF/RW8Z920zDoxByAif1km2k07cwyY2Qfr521hY3EQF6Ot0I/p51t2NqYuomHf6Xc62Rd
b05jCGJ3CeUVFsnQmHWAiXhX0tB0+UhZYRcCWB9wnlX8wGdnN/TXcjNVxZN7dxZcddZ7AVSyVCPL
QPuCPgUoWpJn6WXBqqAci5QUZemI5PJUvNIBx8aR/Jlfoefca8TcTA3jxVLdI/FjhJNAVGM9c9it
+SHLSiPPnLW0gHfP2n16MhKjfuGOo620ptDWhRa4QC1IpaPah/bpPKMgc0izHCa5ZYSSq8W/TYEM
q0FAAPp5XrsEvYVavmAS4fN0G5vV1E12LJNEUJt20Cx9iEEr1sDWPWP42+xrGLkxUoHr5ff1mp9h
scmQ2RnLdoos9optClaMjo1XxSaeJ/CvxDVAjOoJTd2AjycRtysd0h1zdyNBS6kJxd6xtPqVnfGx
HuPK124st+7/daWwB2QalORhfsdCEcitOKMOLlv21KGhTHpB5yV+bOGJZq9K/B8eBEErGwvpOKbN
KP0ewDdaMHRnMy9SWZp1Mrv95Kzjse4nQwoZhgbwHv5NUY7uw00HPIIuQONZpUkTBXfox9Ar0rQn
s6rfQWILlBE3UhCBo6ebv/3ORPVAQGXZLggkBmZQjcspS6MaNbkwmXm+sUpVDc1K4sK75K1MSFyf
IYyZ+bglRADLMexCYh+XNFZbGLXqjvo7uOTVANJdxoNf8lmruBOPpD/QzDS/8uG65l3etFXtkdsM
F/rL+0dgTTpwj8K9WJM2SQafwGYXTSpo8pMoeSPzkqZSJ0L/nokJM6bkK1oTDgzFeEpYxmnGNsxh
/9s9uGKOT4OhJk3HESbUSS36/S0KFpgr6x9iv87HIF6iYn6DH5tQTvEyGfQVVRY4dNFeZH66qE1y
U0Jaj2vxRa9T+T4jf5FjTQvXGP24xQhdSlYVfcKX9bcW1FoLGSTMgL2s6avwdIKDhO6VPT95Qetn
y4PNdiJmpRLyDoUQUkfRRGtrDUHzmZmzLXK+nMT3fLjlBsk0MyB8EgF5NBnyWGbeDitfVPrEEyF2
p79lEHEcsjUmB73TJ13nYRdPIf1YB6ypQr/CpJp0RkSkVeaW135Bh1cAuj3mWLVfigxxgKQ2d8oN
ZmGstabp+JzbGj+EtB8DEGzPCT6VtzxsHU3X+sYlApmAN//fqR2NKAOohBz7iGvyi9SO05Xb5BQQ
Sg1J/PxsRAjBqk0W3qFNKSdvnOmQTmJtyEicDwWmi+QCIqZFVs+MTgJcX71ajjvV1yqOrA/J6iSJ
rJYk9a8iFvZyKAUfMLtzz8+fAHnWONNvxHYo1S6NFCFmkdohfiRE4I31oOUNt/4t6b9ux0h3p9pF
In9ajkCQx9biQcy62jdkRu0sIdTVZ9Aa8UAVFAVQZo5jL6OeQaF/ZbYGVLiKEGDRYBE48Z39Q3o0
fUmee+8pHd56EtI4C8YZwQwf3HC/8Qt46lHtomEhU2dg5NKwSlS5MNHe4poEhMjRKOYpHy6x8mr5
zY+etCzQ2M/e1X+0EZ8yRLBsKaXjk2fJlv4F957rdsVK7f22dE5hV3224EtOkswguAUn81Yo9OY+
ydzjH4wavsKQPkqBY+cplEa5qu1GPKnz/n+EzReyi8szwbovI0IC7cZKhK1ru4MK4xJ89uPQ37Jk
/wnnlqMOibunUZmzpBHsvLPoQNU4Ms/X++q4mz+mcv/Qn769jHdscMxmFzG9NVBAp2wY86yE6kY2
r8p+Ek4+CRLzWxBt5EsLOLqo2xckxz+Vw1Xtcao96ZqWkf16TuXZdZr32cceDoY+lzNUPJC0FpdW
IF2m2MNzQZMemKUb8QUBogKwnqNOXPZrQCmdlNm0ZwFwv2v0XgEAo6gs95NdObelKmEu8XpeMUtE
G8nwO6W2mjlknxH7vke9KlA5KJyh/SiqMvYq90opkajWwrpuGP6F98f09SGeS9i+pXTJDcB6Lp9d
11blYEbtQIiUrJMg0oGWdMaoYbsa9pgmWR/FyYT368+6vcJK6nrXgcXd3T5RFD57mXN9WGnOhEWo
g91+THb8aA0xd15s1PfR039xKfXotieQcNo8HiT298Wl+voNJEWyXjbIp4vunKbrrrfO/vTdZ9+r
23P/WGM+zLprTJZm1NZH4rbMhV7SF1VOCOJRSAap2oUYlkdN94L3OKcw2raf741OFBIWgtRJSi5q
cMLQyWA2ayhunu1QQO2VF/rTTnHIf6W+9zvR9rDTnBqBIxA7BwOp8EvvKeGCpeobYRpkAj2X9c8T
53/MWWQ2CEUzMQJPXG90MOX1O096p6uC7o5lVa923Pr7q1RpcHZhNKmfHrm0Dp6oze8/MXLK8Fhb
SoDXR4zcC1pU2pULVOb8Z4u+pOw4X+hLQZ9QO3qcJLWbiL1m8RY1Mi3OIkXtFHE3THQyHtWGjsHC
a545RQyCnNE8tPjjby64MRNu1KSk8PpzpvqZjOpEwB4B4o/o2K7jvE+1da8TNVxKdQh/Qs0XCiPV
uMj0GldrOJ7WanWNclDVYgd7VG0/9g8RDaGynouLO83RrrT/Ezkkh7k3DllNhDjuZ6URr51qzlsZ
o9z2ymC64+i4o4HpX/uX3atQUVSo963z23E/kPZt55Qt4fOwoKOh4oHQnbbWe/lXv7PJz8bYZi05
UnI4IlkAMdQIO4R3X4P291LKT09n61aRTUkXlTZUKmEUYfXTIgpuTu7n3Bk8MWKPIHtG1KSMM1Ui
nePNQ/7fVkykDRo6RJ4jYxqEYnA+7hxCT7ESGly27l/OiUdpNJgHi1qE/VHR2LGf8nNY7EzBtWIi
Su2u8MCg53hJePHk+xNuG0rG5gKCGDm7N+z6nd1TC7MCE2J/KtE1Axoc3bv1+Cfdz7S75xagxJdc
diPRQ5QkyuI+5AHg9be4oDSHLf8TpuVqMbhoBqPHcfIk+ypm+ghqIGi8HO1mVthGPZenGZC4noJq
cCehYHHsgVopYjzpVhRpp0uXdUIYoTAdolKYbiNscTfZnBG1edcRf0F2P3ZnJqsUISGz3nylI2+D
YwtGTW6HikmNpgOfyi9aTEyaFliSXQKdpoaPQsyZA5autDkOMguh1uBs75sOJoL8zqUPi4U6njEl
qsPyhR52lk1oO5+fpv1PG5m2OhY+D8oKGUJ0EQiiuCIc7Wxz2K3H7kqRE728EXpBPr9mDv6wTrCa
EO8A4+sQUgDt1GXih+VnSKJqnQykPs/PPUk73OifdeQ36/aNYUu9PyLEBzA66M30Y5RfxrWfJ0I8
rwW6at4fP1NNVTp7A4X9EULmaTqJECYlDDfdKS6Yzxv0qESonEw+IIY6JcYuzGLadSMSoyEQzruf
jIOC7JkAbfQyUBpAS587fJ7Rpv5QPyWGWrRZSy8dLWs8sQQkAmWyV7jQcVlafcuPRozV+sNR9MZ3
3HKy7DJBsi4B169uHEKYIuwSG7Oa/SGNGbpd57nCUpzh8uuJCz8rtxxi6wVbh2iPDhwhn1aWhNMl
RavCnaCk7J1cFAf0q1YoE+aUIzYzPcaNcpw834fePpQyycZZB8BO84w1Aw1dcnZUQGoHqU+NhUZL
5cBngZh46jgdUXkERP9gVKCg2jZAk2UkKdbiiNGHJhbCjtPDHtz0BjuFYHD3cSvoip81kg3dHmlC
yL8Aqq3kH+SHuVSYu9ip4Cs2BA66rohNQe55B4QySl7870oPDdz/Ry7/wJXWYsQREw2qa8WvT7Fv
Huwph+JnprQtS6kZZp+reh/Y6X9oqr6sadq90xa5zZExEAw+dvLukVrukr/yGizwqCxLRYMAU/Nl
qWtJa584czOT09vFxM+wpkW+G5pjrIdHp6EDYKdL1HHJ72QJQKJDSS79BbqceioRlV8hDma64G2a
0RbgH5f8HJxd4w8mth2XgvR+UykDD0OzCEoDA+JrTUrjnpAn7UczqfsUfac7fe7zDBiUL6S8cqGd
1jN2e6wHjTgti8aQ16/it3bP66Y9u6GoHDKYzk0R/+OKEPPO6qH1vle+Sb7cQywA+LzJZlWOYR3d
hUSs1bTpfQKYvNx/w9bCndJs0LMFUH4bko02eFCFe4QcdJBa8kMRrshkem/s3xvf4/t+fptXs/s/
4h9uERPy5CABppPgus/Du0cD0ZjXrZ1uV3QRi9E07vUAItBITtzJoGqr2KYBmVTFgy6xqJUBxXaY
4FfhSo2otSl8J7MsPRgKrjZSiKPKzcYzE54EvkoGtNDHFW5MZ7GeVnPrjYwvyad//UIuYL6jX5eR
IHqSgRKcnk18kQn/nawh3zl3J7mx07IlpOXwLpUc7WncQESr+Q5jpOiMY8RMAlFaDytznAwlqm0R
aAM31K6F03iWG2AgN3ARg5v+dvxdAZ+MBgB0y7fZ9JT18B0IlTjgXoGNohlXmbR6NeIy9fT/EXNw
PyF1rIASl8DgleA6bEjmZvKyRTiu+nxrfXjQMJETLiD7atuANyvsa/kxDpv/rijbOihdle0cn0FL
vHuLkwGejZOSolwGXC3bBPniYNHtGYIQ+eIyAF4xU8SF7q+KVkeuvVXRrpu9QEJtF+TZ77o5dWbH
jfW68yEYIwNLDvMh/Nke7LyYL5sc6UuqiP5yhn1cLxqk3S7JF6bXXcOfz1Vb5JNRXinf2o6DSgPK
XF3WUh8exceGsCNdZieMsYWaqj1AZLE3cIfjkCCuUJ9dEKMbroFDG6eY3XSdAp69RcXT5jGmDeUi
Gxs7clUDLMNgCHO9KzQ8dr6rKA8Yuj6huQq0LKFG3qIbw3Zn8ao7w2P6A+1vFXPkHw6XpZWlF5Jr
lyHqAVU4IZRRrgC7Qtqq5T8pPgjIcGiVgisbkN2byWHayhgkXdC2hJjQMvLplKOTe3++iXs0JSe5
g0Iqc7c0TJ84Y9fdulNcZ7I/e+SM3BoQ38CmZZT2y+eaSMmRu03o3zrtD0/WbtN5KMp15ggemK91
4sHYlZXDV+M3rhciA1/mIIORmQI9wdahtN9M3eupOMCaYhpj0sjAqY6qt6ARiREhF5xwtvrSgTMq
PBSVpy1NGdjCG5fGTLJohS4KI29tbiYqnpu3HM/Vbn5gYXuSeo/jgSJRMo/dAaarcmi+0rbi8+WO
S9FR1+G2H3joEgeDaWiGlkImJBK0CNxmu23Ij46y5SGI5RnpAnXMr6NAbUOA+kawSsryx/L3OCrH
EnjARAr65krX212RCaEA2cbTLpeKg9HGiXdCRoCS0uWqGwN3tmdnNos/0Wswoft6NmZ0EnkuyN2e
HT3wj7jP0ODWLHwFoA5wm7hrEq/blVZ3umwk3ZoIdzWTWPdNUVnCICaMhJ35Z31p86RGt/e0fOKL
WeKxIBPIitPWVX4K4PDrtrxKTa1vJAxchQEWiJoDU4Ia2tWLkll5dj07iEva3tJfTNaocINxndo2
FW2Huf4Il8RHz+FxQqw7EqOcKC86U2+c+6CDtIp1EMFoE8PC/c9pyO1wlnB+oxhOvWs1UY40jhcu
KyqaUY51Ew9S7jLgPIJLah7XK2GizAe7mcSP5wwpIf6P0yIssbxadUB66+ikzeESZ99+iD3sPykG
c3FRkyqn3YG7tEcF6s/+0XOkAfUUkOJmuz17v9YUyQypbwrKNeWS7s3B26xQ3J+JRbUouc0WgpAb
hjzyw9aXYkahBqwMAk4EvHYNwStsoRVROyX4OAZd/W7BgE2nXLqSMshTJOUPRTwRPAB/TCYMW2q2
aexHwkd+0cxABEAhzkGhyFCFgm0T7lBULtfDvRME1Hy2esHaTi/6NJkXCuY4bjDwWPLR8olZwJ6R
sLbf9h2LkKgMgbQm/ylxQtMqT6yrLbjmca4fpIoTZxZKgcWbuNjq2Dh05OexBl4IlnrlA31VmS90
d0XOy3r9HH2thE5fG5HEUHMMxGir8mzQiPAIL26hQcQWfVPXLMmlzzUwjfezwRg0jM67DlIxRdm2
Twlw2VrlI1yW4lvlpVddwbo61V/STj3AtnglYPM/LsnvCvxk5eUmBotBlk+FS51BVPSMn6GEi3zu
plnBHIDVZSiP7zogGfvVBo8p7Br2Sf/pCRag6ekaRvXXFFbpyeiDpBe7Q0pb9ts3Q7Lax+W3IMwh
MUnq8tM6fFL6Az5KB5zW3TmlVPYFgxjdOY+2lJHkGbxH+jE3bNDQyazQ4m+l1DHAckdY/UxalZQM
wAH6kD1e185tECdRoHhL4hUHx4cvDrXfGIpQtRZmOQIRqJmJWBdOeuAi0WvOba4mQ60+DQyEfHxH
+t6zOhCSqWhajT0DUCnAOhv+EyfzPLy2yqXLBHo50SCflr9zUqHmp+UOWh5xPDPM4FPmbBNXTPDJ
1kmmbn69aR7ZyM9pcxnwYTD0eW531avN7mDcvJu0M/IxL3fjhdyxDQGrdWTy3fMlHcdJO3ekip91
cRWzC1bWFukNsXWWGG43lzlsbXxDHY0FH/l/IJ3oxZKHltbDKZJNsbFr/D3vZzDop6Z1bYcJkXZv
wNPy7BCycHQbKTUBRP01xDwCqsyqnLkQS54krWgZmkD5YM8oB/otVfPdFZgAKo/NzNxupU9Pyq85
s/gxDmb7Cu1bdNtbkgw0kQVfJI6Yj2i/GuVFIDI5/p9TZTD2nm9+2/HRRAhmquZmf3rqqPO9TNHh
++MF1Ctm8fBV4NaBZiShgD52cYw9na+RnW7LukGy7pVk+qPoDhr/lAPm1JHqWpBRlgPZtaTlKap5
q+RXWEwdXwwM9H0evyTFIwE/aYq9DMgl7kSR1zdoDCpOlmAOu0erRkh639fBytezXSETYb3SJaVi
8OQH/AN2C//ZWamiSlyVSmAIWsfUOCNDwjHMvhIFmJYp4KyGWqWsdGPRq3zYaFNJYvwd/BZFUl0f
J0Mnu36atJNlrAODcbqWYhvvjxSinuBZYut9yG5JO3616F6wZ2gZtPGbQrMbtYS4Aye8TruKiYvs
VJISQ8wtsXsUrRWrSfL0hOQiASu9HZjLIVR37P4xTVRjmJXWUvXZEqWVTCgH5ZbaHcgUbMHnY4NW
cY4M1kEJbNYHn5r88nJZhjWBihJabLWc/WpFKyeIdXnh7Tbvim5ztnEQLtY/8E1dvEpQiiXTmxTV
O95M22714EjtIGCI2DzagTLlRU+C+pg4dfCvotP0PlfLCAJer9A+SxZrtsz/gCzyAuKqEsNbSQU6
cVtB4r38emP6Us9M11MoV0aFs+inHrGORy8gQVBup3WpM5ICT8PAGKJbqSshNteei/2cK/oBWyQS
nmXGUOwStS/V8+nnXqQTg7Z9gxsE6+eQCxjP7xHc9QZpe99FBua7k3wRaeICmpZrRfzVpnroV9N6
uyG4wQ397HHUqjXCF8c5yPy7vjSbRAF0qn1hPcBO+N6LWHqlDCDJGi3jRxcnvHCsM+UrUfBHKFoz
WnTq8oDtywg9Z70kIo7cv7H1puLkTdF8NyPLCi/m4lGrFX27Zpz8Nw8Cvn/C40dZj1bRjEdd+rq/
FUU/RizfdZHh+41QNG3dSsIcg359rvMVLDo8f4x6s27sLpxH36Lp3cIvBb0ZlcHSmktDjL+1FRUW
eve6/QABKVwJFN/wXBGtJBG+R9wqTsy+3Iu92/5Fyu3yCLzJLDB/Qg0b1CD6MzNkxrmzsRBrgxpj
po7Ve3vjctO3xHj8yQeM7jCaeIxWvZYrhxtqQDh5Xzb9PDZUHL+SkSTfAmhbtYVG+tkOR6n8joQ7
CRS5OTVAoawE539AAHz0XlMcFh5YtiWys4Zbr6Qika9yrTwbzwT4ZJvXcEYWd9dJrCWr0RcnEQUn
DUbN6nArYRZ0gqVj4JovtZqzaayFtKfCmIb7uaUAjA6NXo1DvQ9MDcQd+p3wgYaE47WKW35KVXD5
P1BFeX1ptkSQoP8XYmn6Tk6CU9EdebTpyhGv2O9oTejeeTP88qFvYyOR5G0NlsV/FhztdsM7AkTv
l6bP+rRzxSiDmCv6CgX6C1bgOXTbqdyr+Pznn+02piLf+T9hF0iZt9FA2KQIZg+M5lCf2VaLm/7k
rsqC+Xb83DgpZb2MQJpd/G51Hz0saYFjoGvICsL2VUFqgI4spwriuWhje5Kab7bU9vGbuHSU0QO3
uPiLDoHRqR32zAcwHITEcZV/A/DUqvzK7p+UTsA3CankKy+6jLw/XSfV+vieYqKtFfkDm1ub6cfn
zw3TlkSQtgQQ+X2Y+SSCXSJ/rnhdcOgH7M1LCzM1YPd3zv7Q+Wfs0V5iUil9ur9C+V1lT2Y+KTOy
sZt+8UPgVUSiXoXS4lhPo9u3awZSBr1jmIaKR20x94meqXmoEsnIqoHXp1ZlypOU8aFBT3HXuhbO
if5Yt5pEFZCys4tKBglswbMxWn8POCdQqsnGpA+2hsJs/VIC+JxX1s+r1rizhTtPxMNrhqw4xdsU
9xOm4CCxzGQODbRIxx+MfcCVEEbXmpl2GTPwoOGFNi/e+IwgmFoQmSeuvK0nzUM70d/B9f+bZz/O
moreaZQWuWr4QWl4NLHzNmPwSLJ2Mh2wtYZj2AU8ZHJ2egaMRY79+QLzKHLdR1sM/dsJk+xI1Ql7
OH2xiZpcnzExNaeNE7MqCXGM3LKfYqNxN86ZUvkr0PPN6izdqdVGHSOx6w4S9FFosTuK3rnlqtlT
3lFKI7jGWtpxsUJVeljuoCGIVEGK5DncwRwWUl8cEX3C2L9xVJIVMyrrPFQOrNZKZk9GTKXC8r5O
vdCdkg4dKjOrWfdYtGJSkH6WEqymYBjG4Xm70MTicFDrSE289VF6uwIqt+8pEN3ruG3RK1HeLiWc
LHGoIjz76u93mjH5q/cdCkMuYnlJtwT/vq+m8/gYkww3a/KWNL+Gserszhf7IqYvkATKzB5b9uQr
bQXgMSZzYHUt08Ig1pnTYWTVGC+LHfv90S165L9jz2aMntqhhzQSWeMeJwYxmBP7Jx+MOREuBgNG
vtCRwn2ufglTgxN0WsLAQVCkJSebsOI8vRj51miOjP9FSFbuCP++Aa9laSbWQ8/3IbeTut2N+/IL
AuKTzfMH8JqlMh09X7Lv9wxQ/zDh6t2ZOolimjHmI//yQebNNysrFh8jebFLTztDI3RUQuXAw4iP
GInaSfGdOdtTpzRpm8RIguyfWDRdGQn5TC2x/ButWY/zz36sPRCnipst6UYDWdPHMQCvdTC2Ukpe
wkQODRIrGw+1EFtIBjaCV+gi23gLeY43C9B1wCUdLUWHdeZv4UgD1iyn3IBjtEjmb7+o61i42+L4
mMwbmD5ssgO+yXAPAyJ332jyNU++PhhGRYThilFCrrh+GGWBLRvHTyM+ShVYYtK0P4KWXPQdp1Os
Wmgv/Dr6BvEyVWZUbTpIbEa6smHM7m/4rPKEA4AVvlGaLWlOz8sLvsHuVLUkxxwDQ1SMhTZ+opKw
FeSXumJtgh0qwtYW6BDOy1Su+ID9BBst4VnShHEPv0D5IyijkWMBXGIcjGMLA87wGVffv9bJb4Q7
NfN623gOWaVsJJxGtwD4/ty0CpNu1GruLeNYvpa5Tb3K2sPRzMNg8fptllYTTdzY8PDKqVkADOCu
qaR5R0+kW40jvcoIifrYXJRxIiFdluqBkfd4HVRNPPAA8PFx7qcU5eCM0rAB6q+uGA7F1r3AMjzq
finSLwher/O7FpUgxfx1jmXuIhyDiVzZ1jDk0po2+RJGyOZqUHazJQsTmfjOh0xc4Hp9tLoub9sv
VUqu4Og8P4bNnOmOXsFfWTkjvrDNGrdee2+OwA1NR4nlRZ/BgYEnljTmavvMkDhB7vovY65h86YF
aaf4IzhemVsDKnhEsGbKPVyY0yUlqCCd/nn7mDTLSZXY28bth5FkEQ7Y+4WPK4CT27aZHF9dEMp6
DeF3IUx2h/xMBbuGlO3VKTNcNtSBWxHXu7FT+CZa92sURtYqj8w/Qsm8k61j0oR5Uir17DkukERi
d+l4Heh0BdUrZyB/rLSCyoWeuTyBGkXOHHyxQjveFrdk7wXXrtM3zcD8UGt6cXuFl00bsoosDPX5
WldpgISa3iZQwGOQgopM9lwa2MHtI4qN8OYw7iO6KL57mOrvngd08HLzX4aA2Uduamhaj78iEwES
ppY6XiPMnt7mwc3GgBZF22FDmLkspf6FREk9fYKXYyEFftJsd3ccVcpHq2Pv5xF+huRyRtiAN9mh
/BEsQz+db3rnCMpNo73moAUmy7xf2v4UrYZdM3Pn+/0KD2wTDz83RzJPzq+nJg8ndKwnTZohvkNI
1M0Buq3B3msbz68MRXtYmEph7el8lzk9LcOYFtvjlWQrTtLJ3y/0isXV8mcHrcXaPaMQI8Mdfp4l
NfnThila9xgrk+QFgfWJaaCNrqrXtzSSINsNC1bf5bVCerEvs9zHKMANtGwxfGetE4jf2wSwU8oV
b9u0xa9UM8EW9OkRJ02BbWMBfOLcnSIWxChxSYhSy6ExmHv8ksONcS8XffgrinSPVVTAvobPhdoA
5z7BVvmTbs+wpej4CCWoEeREJfPqoZsg7GvT9bXWZTSyW1/C4lqUcT7QUviEvGJ1kZNZOwBv/RYX
O1oQtwosSnO5q+0NhoZ5BspVE3ZKHk/ci758kSK3lC0f+uXp6fH6cXOoWuGpdrFBuNQYpGmSHXgU
mwX4V0mr3bb9z2JxCFalyGhYQubJuHS1F3K8QVrmQlvNRVriFHSV8GuhLF0gayEKIYsj63nLlAJ8
cOfqOa9Ngl9xKjzIaYElazksHYaHcWbqeNJn+LTJWGwdcqeGEr7hDq+g0U+Ug5DoS2d5NvS3Man5
tBbSaqwioiofHpxHesv6ovlnimL0SbMCZd4wItcUfMqi0uy58YK2fm0FlRh2GV5D871jvInLpR5H
6MNyQI8ZsUITtDsy4mx7HiuJxdxwBazGFpBf8vctXUv2ss5ERvDa2HH/LEXHHnISKhboujqQ0ejY
BDqMwdt7rfd6lPVefWf4lgN2ALdTqXJzjROmHESePHvHEwXVXADnryHDJkcv73SBBmnd14+3212y
hdD+ypxXn7DE5R0nuSmHdsIawEi6E8/oW/1cdCPIpTVwjNkZPqrtAHgibkTrVOmwWiea9kZORJi/
NOSUnHy64XGXM3/Uz8zGkmzhLza//b2VqnyMRw3BorFNWAVp2EFEBf5FOCZS7s219opHNJ/WSZdY
gmbM3XsRqEQvtaCNK2Qi8rHtUPlxGXOno+tmkpYk/rdYNLFbQ1m3LKYhJwR6yT1bidd05JCKn9dO
otqvQ2DaXYAG0KPblb4l6sdK7DxXXl6sw4+qHNqZULoJRzPLU5sTLzp4fSrRxmmfZVdsSvQzsj5J
USCkWx34G50Aty8Awx5sM+MEg2dAhKDutOcsTuQvBYZVFRpfN2JKXU1/NHgHxk0/kZ7W5yZwV15Z
ANGa197I3Hf7SyrkjdbTEccSi9XR0ZxDM0Awcel20T0qal0rCDxPuTMMXEEdegENKue5ELeVLbIR
zniioDF1Zu4vt+NTU03Tw8/EVAGXQVVhik/QaFzH9g36OLGMgLoHnfPu+GuLhgzvui+B9yXHWL0T
pUB9t04NMPgQDnePC/3lLt7cRKrH9TityEK0tlukr3MvC7JoFlb3V9HITQZUyVuJgi06IKoaudW9
DatYYlVUQioST1kJJHF82ix2Yb7J/Z92P07U+DhDpRWwZgFQ65L7xA6xDw7fpSy78EtZUooSI0hr
WCYJM0PWVqpPK2uwZRnAwmZfXV9bxGIAL+QuBowgKaqqSxYXXGUm1BHlKpx8+kThLYkuipYrl9Hy
MamBcRGpVkFR2h2EBFOanxirOObrvfwzBT47NX2u7Rpvzuk+4aa+FnTmZ2aR0RqnBOClRFBPNIrp
/m0kW65YLwf0bKBEt6OgDXIXABD3kxbOdefTmAYW+McBwkmASQZO93w7QQrwB13475WM5XPwxORX
FYXhI31Z7IWxHu7sy/MeInYc/BMc9SDiUlmh/QnxfkGDMRZbVjyiyCD7YXrD3F+3CvLUxEA8MePM
Q2sWZGZ38Mj7oxxCdYPifTz4cRFggwtOBK+RCyfHMy6VicO2BoBdSw5FM2IVWha/AJDv302eWLou
vtYxBkId0K0RSN2+WXXsXFvMtPzPZ7YBm1Kv+WSiUvcHjeWwxjOa/EVthsoYvaTdI8dxogYVC33P
ZhOjrdy4G8bHCLXBQCIRTYQod5sLmCB0hJT7PPnz0SXehCkeYqnbHWtn3imx/66PJHKK6Gri1DeJ
C3gXuSVz6f/EahafYyBqDiJ+CTS9jvIhEB+lMoUJJZ/I0GlMaNRoTAQVEefC0/zErwY/oIB+G2EM
E0IwnDj/mEMO6f0vDCIQu/aN/+Zp8/KMx0cJE6bKLCi72xDg9rE97gWLa8zbD7yOpCB7C2pGthLJ
cmpHrqzf61yIXZppqS8EiV04cHLd08euup8PaIAwqFDbvupEaOKakb1Yk14a62wjoRcSJjvRQ9m+
v1VkoRmA86JnK17PfyANxMVqxhZ38DC7zXvwly5ntok2nO5A9C71Fk+aTy88ceDJ6WceU4q5WK3O
bZJnE4MvNOcdd4GV488FqZxfgieiae4TWeXTHF6ZjXEm6HPw9Nwv0GZhywWm/cUbwaH1YNWuPxNC
cIRH5Qhky9avMWd+q5Js9FSltNLrrSaQU+byWnyBnh0m86hQKRO/rrCmx+h0/WrARZCTtdN+q42I
9DW7UuD757rB2wNdJVw6SxGL2zCYubPcwbnJVVKsv7rwHh0pN3S/DT+R+Y4xjsH6eiQ/6iABqq1O
mdD9jEK5iXrgDum3RRDCc9bY+42R/yA6zd1jf9Hqd55W2ASadbcf8tm/iGo+d3fU24fqRgs8uW9f
3DMtAMYJj4Vatla0SFyvhbDlmY/zA5YklRIJDKZYoA9s+3etNJD8/B4R4H++0vGg/eq85h+bU6FI
n7kjh55Kwt0JsecfepbH+FAAzRPelH98FLkRuT9cFZd56cdtbEJjhkDkz8yodavKdbW1vYsrGndH
8/kSENJwqa0pUB2weZYVGMV3d8qiE/nJzI7JmMOiuP4WlEWfuy3PsFaDHTYkjQS/lacpYvYhOE/h
Jy93PQCH+a7SLqa8G7F90E00tSzENf1o6Yctp7Ls1yqLCttmcOHuAyRXQVZa0RWmrZWNrnNmCKFF
JmpYMlACOfCcQhjXDS4JH02f12p3ZrRZi0ZFjif2oQcQOPune45HvokUCNK7ZCC0xWpIK1JeiOP0
egxm8OGnWlf+9nIBw2yqq+aGEXg9NRLHUJfQiOTr+KgJueAUu8j3XlOxCK69xjht+EtpVEDQVlch
kM8FieO/++TC8H2Wd2oxFB8iry9IBYppGRiUYb3C2Uz1K1Gwz8LmzvFS8k3jO31+qsJDJOOtNC8G
9KmxjuFRoTNs2bms+jG0lgMlheTCXVhtAvGcrQH8JAs23545vICrOVEvs6DSK92ebZTE8LfSEe8p
PoqLRuRA3gjoSZm+F9PSUnkKtcsxvDk+AAwYTr7CKdzu90m8TgV/Qp6WUXpPWWhsMLgn8Xie8V0L
LeWjU63VLhWjDWeQBZ/Ahox4GBzxDwjoGIlEe5d59HizznyYymuPZ1QxDmjT8tA2VlYRhnSySyuT
2JO8/+RLUc+LZ4tfS3ObXaQ7W13tnG7wWBvpeBE0rld8LxnE7OTqfR1hs7IuIssDYGTJ2aLu4UAI
GgJafSkv8iDHza+ZdhZDrwhpwRmQztoi1DKl3LjhSD83U5om8mmt84xTk8zX+z7qf1+I1RhWVVBW
cbQNXWdVeGI7na7JxGAnyDeODYoBGhtHlLc7vLWVoNadamlWcHqVq7CjNm9/9ppNAAcJ858Bx7u6
wLHK7O+D2yCAxYpK50bEs2FtoJKuvESbAjZezBaswRv+fKuR8Aq+tGJyMCr88zaozHWzOhs5/JAd
D2IY8XHulnOmJsoXrzAncwf00tqUmn2cDd/xddLRQnqajg72Yjm2tChQQrxudJYIM6ghh1aw57t+
dnvA+kh+dcMytCTLd0zklorrgtZey7MDZRA/wfHyvpDmMpkgos7dBZTPDMW3wn6/GnrNvkgnGh4y
FO5BYZpogpVpzi9KnoNeELiLSApVVL3+rjxF/93uhPBCWMmD956ipi4HdacBmzC5XQ1Wg485cV02
J6tkikCwGNvkfCKw51geC5V2YYQXZZUXGC5D1/T0UEVKfvE3hqqtmO3qd1hIZjrMPR+WdZhXxXNF
8/boO+9zXy8VQooZonlG0FOu1V8gXrW9b61JiyozgyYnKuOjGRNQudcRDTA9LtrOziIFeIA1myyS
Yo+wBXY0yZJ3z5R0R41cia1mho4NJLYss5p9HMoGsXfvltCRd/eKoAJ1JZ1/Bsqn5YvQSoJ/i/Sh
6ojGykqbZzLTZ8ZYi52YWqUI/6VNfc4a/vDna0NIT4rv3vx6uRAaZL4ygX4ADige9wP/2n33L88p
D/Q+o2TxyeN99jQeasj4+MoTdenKrGM6hgRZb9WwtDs32i9s0ZwZEvPwIMyeZhYChMGcEw5mIg4z
ujn4eKsRvyd0GZS69R+HTu1DUy4bkK8oRlBjywCHD4QvyClFoAF7M21KNMhdzYXsIe10LXqa8q9R
WqBbXK1bSxKyZu7L8mCNXaRIBBHfCIhinJyMs5DIq/WF3spKk2CjWvfx9k45mIcpdjfvPHzHASdh
Oz/+++KXI/F5AAYorLVcmB3yjqn03To98h1/eaQUi6ty3ehqFZUJH25LJuDF3C4JFD05sktpMWyx
Rf95Rul8K8TqzmvGfv0TTkQyggQ6d4Bc6XjEb+QFi3TZ+eMB9dXRPZMAoGkkMxf/7HNo9zhVR/+J
WJMvJ9qJw5ByIGXaj9LH7yJ7T77sIzHtmprNUzL3Bdo8FKjCvDRFW9NrOsDm8i3ISu8QJZbaVOKV
+56nHsoZz8TL5dq0BLja6LHMaUpvkFbmQ/nMcEy8ZiBRbrtN+8ka4vZngF3NkGphnNFPIC+IYm20
i7i9gn/MBiDITJuantU9akVjuR0Fs5spVd1jyj73XuwcJMNugSarHf2UxJonokZJS3vwglU7Oqpf
cuU9HWVpsP27zl09CB6yWVMN9ZCiXB1F5GTpDrudfKBO3niwIvKNLhnwA78M0yrNjqAHi/mTNf5G
aWx+K6vsfs/LtoMi6zgtUJQy1qgIU5O5RBC5K+pWHe1wsKCJ1Ae1Gqkdoq/kaU20z239AgPFnFVC
boTEAdF8QGaj3fAc/VAeFe1ewHLVC5g6yrDJNAnGT7GAkceiB+OMm3Pf6kDKafvMVUjrpaVSAHHJ
80zQu+vAxxhdzQ+XWsLEek5jPtrELDF1MD0cD0X+lBnoWM4VfIEsCb6ng8UCNdOF4DJJFyqP3P8e
ZCyW16MjFkim3XTMe21Md+wPkit5ScTpJOE/eX2R8hY3QOQMnZ+3wy44MT3hgrtIvuUgn/XCwi8L
TxIWAgjbccWnLFZqqjF0x25p+g2R9agEXi6rCQulDEB3E4qMCFaKhgr/EBchT/GQfKvRUubiz+mF
tl2ARBn9k4jJrKC8UL6iE+/ZjRsV2QGtXGAeoN3Cq4XeUZdmgOLUS3ZsVzBRdpMmY6cf8xBvqxZS
Wd+cbAfauLiUtCC9umTWJUK5gqzjVJAykgl4ny2GvNuCsDu+ceX5zA9iotY5H6v3QPm300+TGqoe
aoZuGmGLUvxMMVvMtGcPTtjkMZFCP++DUW1wAuMZcZEcQoB9zO41TgXDQlnXbZMPjPSTGbwNlaYl
9ZufyUs5ytkwpHbb5AeImBhvfsTnVcbrh0d29n+Oxa3AOX+G8YUSnEE/QSBI7RkBrN71gohBJfYc
vvdNFRQ33/iLVBH5NTRvCCWZoRSUvneETE2LzvbePQqeZyih1g1l0UwUh11FrivB9QTlKyYd7amC
bs2hElnmFGe8oVvfUZd6r06qo/2e/G9FYLFb+7INNwq2jqxVm91ovfAVekoWm8FfwvvEfFqJlVkB
fHZlmSMqt697thLDcq+Mfd4e/0LvOrDOEY7j/cduF+ldCdU7gYDjVxe6HBZh+5w+pch6ZJRpQKYo
0ElSBVdwb4RtY+j5Ex6T368OZXJCPW+uAtw/m5RAaK5EY/cREADe4nOr+O3DdFaXt82PQcDQI6n0
mns7A2VIljv97uSX0PbkKgMfpWqWK5E9NeTpK5mwy7ygwRUxUzE/HtqXdaM/C4xe6LDwgY+KKHlj
NImb7PASRCUerxg9Zg/i09zCmIgX3SfXObUPnew3hU9oI8jSv2lcyd25u7rRICFrfKEPedSUVp1Q
Z0hnURWR8lPBfaCSj9o+JUi/5RUzTldJhp6jzcz3uK8kpk84L+AvaT5LqVLxd7OMoqCNOxRzq1kJ
BgSrLg4dTIqOy9zTcnXa87u4hfrYNZOKpXbMx9VbsT5Qq+Ql5pSFsWJkuAZw5FS4XkJ3BjZeOwlz
kwd5J4V6tJCIibX3IJJFuqAVd4goEE3W1S4j0g6O7Trf1bEUDltI0Yq3AdTZRuoeGtupKFBhoGMj
gcNAVxRQCumj/xjhn1bqFEY6TkpT+BRIfLU24tw2QYfJbQT69QJI7VJJZOLRNv+G2heYzlBdSmtl
h2jbMcrkXH3oHJYQA6yeS1J1RkiVjwtlIi6PqSv1irgLzAAWfLxOW9RjfOpCAVLkcjEHMnFQdPwk
HooyqIRVTYbmQwrFx6mMw1vMP6j/RqwZUMgyHQfMnAVA9LbGua3mBkptw2qo2CcQ1hfSINDYaHUF
tdR79ba51OVQrpnEuiloITSAfRocnYbjdroIq4s5CXuYIUH6Op7Wojn9cAuOqoHYNQOZRMfP9WBj
EPqasyf45CcWRc0esfYCXLBKXsQe3kLAzgDxjqBIUObgD7kGCxmQm2q7NWMPJRLJLOay0NjeJsdX
atJVIrApOqPlLzaYMV48TlauptU3PLrMeocvoEDlf6WKzHyAIiacbxCVm57zJftPoqWdXib+vKFm
xAekx7l8omc4UkkO8NZ3MKT0YMF6aoBZbfuwS/HStBaEgNJ4J5ttG4RdciO2HVfo6sp9aii+aZ0n
Wgf1IQAOU305uT2J5EXTGCIWn1nUB30rxeLjun96rR9LGJqxP4TUHvLXV1HeVz5Ks6gHV9Q8DRol
rBjjioMJ2w3LfdPVn5WsddLLtPdN/KwUrX4d/nEbHwT7fTwypFHUOAwLNzpiSChoiSX4B0k/Qmya
PMHB/1/bUMbdpuQXJFR7fnP3y00Lrl3BqqcStonsctVmCTA67z2Cn0+WV/FKuzhrYZGi2XeWuZwq
vO5uVtjr+dK3AIikAAeOf4rcPMumBVNZYyFssN8ADPbQc4c9aGQb6Hj/NsDPoe1Bf+Z09y8JJ0kf
uoq6dwUAaDMw5Sxk7TxS9lyOYTfD0BDOVPxgktZRQv7oNhcuVrgLBAFjGIZfo1GtCNvhG6aCcWc/
YOVaA64H6dldyy084Csguc1YwEkZz5Nuk4G3+4QnHV1sAX9sYFAWFAMCrsvNgMiTR55FFVzokHeL
gEwkvlxoPg7PM6aJCxGeIPfG7aToMIpAgsd+7WpET2onBLnM1sUkHi7OjVdU8sqrLDNMRivxAFzL
9oMQIXuatT0al59KNijZHWLolCxZFEnmdplRdgB3yfJZJHMZPyFxYnj4Yd8eM2XvGUvLc7il8f6v
r0rBfTiuZsVht+ZAUedgsJIYIVkXxwOOSKkypxN2KyVQqDSy19qz66xy88hViXOIl/uEU8IJ+LAI
mRRI0UfCk37xoqyHPH2ubJTql2Beak0FAbzRq5+oDFc/YEBnT/E+1ZAMyOyQgogvZwbVnoqKAkeD
CrgUpLNGwl2j0RNbr2D6muFn+8nvHi0ScKpqPc0ONjNbgnGijxIQdazZlp7G2z5OkwSgQpM8T2Kx
prw/r/FCE7wFy29NUIq+ScZtm5XqRSMiEgqyUs6nVdo1vNHQhMEU9gzOuOleFLLAQ7v7BDI+45L1
mXfAKF6s90tLZOimp+PhBwyJ9cxeqXH9tBqgktPrFLS5qd7/UIPwkSgqPkOG4Eq1gBiM9pFt7WAz
wU7xZBzd4EOg8N4vMa3bvENql5OX8+jNT/9VfD0Y9CWXWubbNGDzXxBshTNLYsAgzXO2gikx2QV/
MxDsgCjpijlLfLCfvnp3RMTrid/+u6tNWciKSkYQagVb1De8jyAYmDmNAd+lTHO8VeVA/RGYSvjb
P/z45L1qSYGmw85tT4wLBRzpe4lKBci0puuD0kcDjeKSGEvjGo/UveS5QjIyrvnax4YS8jlImu9R
QpN3QNBvJPRHZXloW0tbCtVfiG0o7GESx3rskkNTqKlXvY3w2KJkD6oozfB5fPa1iHRwiD6w2FmA
zRdht7PU4dpXqnOwLqWFwlPOq1CoReSOIUSDevaAXxW2T1BFHPK2plcBYNmUJu8/vr0retu9Ey3z
ujqWh8a9nMJRt/s5dzmIElQGkBuUYkA6NVyVpznQ21Dat1UtVoXe4FJqF1ePmZPNdwKFwjVPGccU
iWnoINgK+9N1+3BnTbY8cJPDstDcPAJj0p5QJ7yrG19hTQ6tC1sKiPfWRoJK/N3GdPx9mGg0LzYX
dF/726vBduO9eS/fAIaRTypOcCZA0hqZv0vcOLudWtlvOYAmnRiWcicqkdZBAUmcDGet7o7RF8G0
OlvsumIl5cClJAPVn0pyriLuXm8ZULwyP4dSWr7pgFRkJ+Vr1abHRXeoJDnl6OqWKJrlb6MUPiDJ
ifSaA8zQgNJ/BEaSYgBKu8tJPxiFIFxXelP3+xVMKFJyRsbbCxCaTYrYCaHZFprEea6VnBbafffP
aWwQqp9THWJoh6YvEhUf1FF7hdqCtMdqd2FCWhp596ThvmOhKjafr3lhbgRSv+RASSzwcWf2hgEX
rwDoBlD2oz/m6XakR3ZYgVhEJHaraG1JuLnWDRkRwMAFeG/kQhJeH+eF+kCB0NM8765FFC+A12IN
kNb8Ih4Hh5qU5Qf+NToXV/dH/hPyMQLzbIFvRgt74Y41HMxhrt/omDsSvdzv7jnR2awiKqYtmz4X
HAufJcmZ5Z2/vHyrOBhJh5KnCOeSJtcXWhQLhVT5Chpjk6KzVyrLe1+qwfz1vb7GWK4WKHwzxuLw
rnUddLDP4rfhfTA74aEo9Qkfxy9UsJTt3DMa0vlxyawuRBdec4btaHw3FuwF7WUeN5UwZLO8ymbk
9uX//7ovXgfIPWSc07NW5Sgn0HERXa7gCibC9JiiS/GfIbpJvRjCsrYWWb8qW8Q9eTUU3S5lgqSN
CUlum8UZQ7ozBqUFnj6UsAIZ+Lqaxbac5eYFJOchUsKOLzY6HzD2ACg1oasXlXfdo2stqIU+2+y8
xR6fF9J9vtJOnYbwdhQ0KQleZ/aksZSasx8Ieo3HVvjEGoiIcISbDPGXqhiBlS/IoKDv8ry4D8SN
9+G3YIKIIeg8dLBLfckk82C0QyOMGzLuFTG11uv/z6DIlC7RtXR/oZr3MxPJ7dcUMDFCxTe7L++J
/Gs7C6oXuHRTDVmSgXZuMysvnuzdpwwTSMP8yKIYyIC3fAwKrRldnzO+CkDL7rSJUpuHNSLkhmIr
bK9PfMuvLGLDh1JQYb3B4i1uTlAw8CMVCMQWl+KFK91uhdCCflulgcsmzufcPxPwVPJp+zYJJE4I
UOpLM/F+6qvyrr67dJYJhpK+l7FrjpviwbpoBoX1aoC9FWCoQIHag/lv2Oyihp0s6lYq5Wxd177p
9F85UAsHbAhX3bOKHJKdc+p8N03zkJnEXDmhPJ3vveQbsQAI5EqI5qcD2IjXfuvNkWH0ZIsW0Dc5
w02F3uqNmx/i2XBnTGsXDHhVR6km/7F+dSf+L4aMnpJ1nL3z5dPwYMCyyTM0TWUw6v7WwF9cCH4t
pHGGmlA9+1PjYrYvbrKvmOss5+/sO711EVOsfJviAVLML/9SKCCJHEDnPBjwlWdtSnhOivoOq1Yv
TOiBtYyWQtf9sUWEtL50jZv1qDsWJnFOMCkoxnwnpm5DJYMgOUPfuWFUtDVbAfINzdpNbQOK0qxe
A2eFxtJIvM9FOBgCmlc6CuZWVcEB1fxKLDiJgpzpnTaec0iFTDIrkU+K4F07jV3KVtdZCr3O+OhV
vZcd2r2Lju9Tlt3WgWPw08yY7Q1lr4QwUl2qH8KWsH5pS5jTRxrElrgny1gVw8SnhlprQKtMbrXM
GuaH90qEQO8hbqaNsX/0WwSvChgW5v2sMWLeJBdXcQyz6mEEM/6NsjfgOpG7nSZ8BkdoMZh6Q1x7
WeHUqKG7zvO+fVdrt5mUXX+ylX6Oq92ierg0BD1kpBF/f3iFLnhrYeDxJfuTA5QSucB6du/4YKcH
k7hgRhEKSqPUqqVto9EysQdAB2nTfXE5kZ9g8ifgmYkH53ofX6NxEwiU/nBpqr7TBKRZEH81mmDU
MiYdFN1TaLiBHxaJxqeJQ+qi5V8raZM3Q2xQwgVbckWwCNvKJYg/v9YW7JOS9YZdyPjCBlqTsNvI
ia6y/boqrFIht1xVyqvEOqVBey9PbEpTNXDd2R1gb6ZGWir7H98bmU1tSLhoE8PCJi5TMR/6I79l
ZihovWH06MI4hhfvCxD7nHAO25+BAYOxUB2HA6OI2nLCAaRr4yzBfEcfPC/gW6tZBBnj2jU9zaWY
TPq4UIZrHXAs61e7bLKl3+Def8JToAtzgOimSxg1XedYfBwHE55Tsm8R+AKcOISV1yzGttl0EDgS
KS/gol/xiN6znLBxQGedpfouIPVudpi838WAOpy2VsoOmLh79xNEEE+YDn+FGJcsP5R0qHMHB4uy
g7V76Z3Z2kF76UwL5b1hn/T0i01Sw63WXD/kCzoMmV0ooOUd2+RAAnSU+mzuWXqKgube++xQ2ZMz
ZoX1B5suYVqY3foU5qjJfKOB1f8CuCAtzlvYo2iJzphCWMLnEjlgNN1OaK9JRNwkevOvnPjYtqnu
CGWEYnlmzb9faTFp0bUFpdXhe0uKcUIarnIaPTgne/f8gXZ2iojnegropTZOCkfg8UzdMUDUVEqa
QVcmjObDJ6wIDAsqGY41WBjbgDz7gKwNAEqArOO6+uspCquEDi89a/b5b/37mLNDqlV/HtP15Zg+
RVIG9nQv9GVYnakCFgTD3owYlD+EFy6fmASCigkqiggKFbwEqG5y2RS33a2xbNw6IDOYL9Cbukgk
Y7Qdd5m7a2g8bnBh2BcrhGdJXfKwihNH2SG+vkDoX9oE1IDsDcztP2sRHtAl8l31x99I7ZKM5VCh
Ykuy3ubgrCNz8MnJzWOB4/j4514lUFrThyG2vzKE9vbU7fXAVuLgSpDwqZTH3h+GbfhguMUlkLdS
hMtJLqE1JzIzjwMaMMkAn0Myntmy30qs7dCxo1DZS2S58dN1+6LFj3XArP8rKiKmuVOTsA+ypKeU
XEXh64ka668NuunIKC4HcppVc4HSAC1rjfDj70tL5KikKa6yLiyHMQ7BY5iYikvo6FcAXwa0Imls
cBcGMn5zCVkyMQeowvflXQvhq7EyxGH6woXG0KfjwgQm16ZWdV6B3ngICHS4bXvdjTQSc6WnGfAj
26QvaxTHPJIrchGbAF/SY5R6v8StXzBXFMcK5VN0JTm4qedb19ZQv7arCJYpHWM3sn+DkHN/MQlr
++nlfebPZqPcIlUo6C1r/8iuyj5DMW1/RmLJOHUQVKZiBUpttwndi6m49fMU6yfsPmbtkwFc06Yl
p4Yl3GmSHPZ29c3z5TU4wzONEsyrEBEIogPC4gy17DdXYSLl4ZtZq9AVTNSjR65MkrhIHd4oVvJm
TUFT8nQkyW2zbUjoT3AD+03YCXyuRL1saIXbPywiwGa/+YTzJRoThCmLUgdtBy1zKlob6wizY0+h
JdND31GtOll+Yu9TpmUV9K7PVJT1mu1dOAo3xXyrnt5JYttfwkac+c6ZlWKTtiMEo1aQxWu4YoX7
7S9ZPuWlYqyRBouXWmDA8WQAwgWXrDh/bVw8OOsnkW6Uh9AzqZqTsMsRIgvPm0J/3qucnqbDo+r0
3stIyMTBVJfE75BArPNi5951llBbrvnFfK/GUecSHq9fwUIcW52JizzO57SxHANnahdhq6yNxB08
+E5OSUotbADLty046OX5C+oSlv74TGKP+epVMCrZPCzrnKe3CbwkhAi8+A2ld5tEd7eCbHKBIeD7
iQJJTu9Bfbs+5nskhTiADjF0wyMTJ4XgivTlbMoU3Uk5UxYCyWCwMKm+MbC8YIv9WIJrO4CxLR3W
jNzGdzEdTCKPz5q49FiwdFbQABIvgCd4RxUk0ZBvlAIXjU8LoTDbYfGF8pAPZHsy5NZMj9bFZ5OE
hJLIHClB+KfP/5rTZQ+8WPCqPOEJoXWrnsyf7wxAuad/p7oF+mfVFflnfyXyjgQZ6I2t2WiPeQx/
l5SHa1Rx/wdYLIyADA4AQHzFi6X8lTygFxqEEiCoEQ3+a8c9Ix8pC3LBzPQOKVS3U+l22kcAnqox
XonDLECAKlGaLoEOYT+KTFSfPCFmJlO8wYyMkPAuJfUPQadl2q5QzuuoFv8HB/jFzI7t7EOhHf59
j0Su7ZxwTlXEKnp4LjfUEgW7M9HA+i7pMcHN651+R7wCcC4WEfVDQlZMBKqPkHqb4eCrK6zTDUiO
5LruD/unfKZ4nh5/3kOOiyIdY+lJNDOerKSgPu9RxcJpiNgYBSViN2U84nGSmyYuKioA8sWsPV4F
Zqc6jUEiKulv9/6avOezXFoP00Mr1pHZtbTQLp1nwY6AWw5RYNSKpry0wHMoy/9nE/iL1dxfuesP
/Geuz+ceUecHhsjC26Z01lvrhkSK66msTWPJnT6Akd8ymxRJbhVbx6EAPXa9/ZRQKjP7LWJ0Zoej
9T/1vnQlpLZwlDzUhxgPAhIW6ZAilOs22eoH/YrqR9+Oo09Bkyzt2brF3YbNK0F9UFB5nhW3siuA
uoc28uDzI+peMQEpn9kKqKBgQl92UbxDuL2mJA6cl1dyplpQaqLuyNt5xDL+c2bM9nKUSBzX3jt6
BVswTy3Ob5x4f3hX+IgnhQ5J9BZhIwvTL828dY8kqUMZMfDDAdKyLhtn0x4YcmJ9MOrJGFHLEsyZ
iIYFxDch3ILEX2EfZeEinrDF8P2YsDxUvjrVx2DPLAHCD+/DV0xCWcsqMu1B7hiPWp8r7+t4Qqjr
l96RBx3Mt87w7cVmej/U7yfg/VfeCk6kRGHYKGsV3qU6iDHJYnaH1w8j2J1CRmefSK8mSF8QCPke
i4Noptdm8GuIrbvnID9tUO+ke5iI5cKEZqXlz335pcRirrFQLP+xCeGHvdLYI+D20aiP98tl3PAP
e5ugpiqF+DvAiyT9ladHA+BJgnH8KiXUE2kcmMppgslH85DdPtucjmYwCiGRk0vXqynvIvD+YQDR
A2EwH+99zvrpgm56JP8kr3hBp5TY4gLODWSbCZ6dElm6KtEXh22I7EvkWmD0u9F5N1CSytpJg4ab
ZBo5Ns1iZTVZ+ZWIi202wM6m3/gr9zOUR6HJgX+yyKyvLqjrQSNlpsuVwYdcelt5VVk1NRcmOGkR
FFgCT2PoJ5tdmXwSItJy2vpcEghGxsqLkWaEN4N1IqpTHW7LXwFTyaM4nW5rx+sexkCSKaQXFxvz
xCWune04dHfvnPdGkRAmwf0PHKZpdbEyA/sUXgCJaQ33LlJRnmU7+e5IRdzt68nl/9WOpoQ4avUf
oamOq+KhIk2sa9z3AHvN+rINYVHKAQ32BldzIQoRfkOlGchql/w7WG4z/doERS45jow7yea88te5
CBOJoNkG0W+crpKeI81FIZTGK/uwDBWOIf3t0H/YqwMbzrcD0mKil18a5Fj6zZj1vbtbLswv//Gf
dhmTBIXre9eBPMfbocah9vtqbtBavPHP+4TdSwvVMj29zw6ylIXLZHVVRfo6YWZ9iHayYvbLDl7e
e/stISpTzDPZXKZICzwVtwNYlU9qPH3fwfeasl2BxfhNOxY3Gx/UkAR9xv6GRsIYPpkThY8k6nYO
MERGCKkUNLpqwAgwr22oOdY+CVjoUuf+rF0sv3kzgo45LMJgJ5Iha71+az5NkjKeMmL1uHi93z5A
h65OjYuZ4ZkYCdbLKM3AE0EhjRoyrDUs6a+uUZJZVnMNAFuAYuNTlp3vjhjwF+yrfnjDiAcOtG7e
NpASYEygk8ehlwIQa1GlTrvKQcI2YVGPpJn0/xGOQrTZMUziAHC0MLapodSDxisiXlK2U/ov9vrc
lbdiYDIQOlRCGmnHifCXfLmn5gx/9qH9ADimt8Eh9ECgID+3gxevgguQlMxmvzP2rSrs6+KT/DLv
322Q597jI2HdP+LtLBLk8MRNaL3RWADHcEva9lsJLL1M3YfxuMnBvZInCI+3WgArI7h7QRnEX8FI
wjB2PS5pfOqLdTb3xRcnaVTBdrurfEkfmd37nm/y/gXVdx3K7imKtD5QEcPar/TLsXipOPUSf4OX
keQxKooqtKInAq0Cp0IXHTx1IQifGzeLN/C8YK+TXLke/1/9O9vIG74LK3/CODFr7tOLmQN8ytJI
Urscvq2AtweDvPpvWXnsV0gtRclBowc7xq7f3CgejFXOK1TM+f3IYFk3DNqMTcORP684eLcq1mR+
uOLEXzOjlOwFiytTlLaFUL9Fn+dvPb+ltDUTT16R76LJd66nZpC3I0Nu9j3Sk+D2rRthzc4UKJ64
EyROo7vCHa2rSxelx1EkDSuYINi39ptrJARza2hju38Abg92j6qb+564qvTqk7blri1YLQy3KQ0W
lM9ivQRku7r8AC+Gk/3vT/aRcdQv3b8xFgjMAMYcPafIkb1tDIoBPsO/WMSzB6jHYnHwL7pJbfdI
M1/i8swVIAMNW6N+DCAaxIcxt9pkJ8Pzb3PCblgcNw9wv6qOBXVzpNoMsHeny/ePC7a53iQvQaSQ
goHWxrfoUvIJM9xNGFNgJahUFHnPYT/ZjT3Xp7FvBVgWpHx9+PjV/ppFbaFd89bObmHGZ0B5PXCI
unSYRn0gR66XmXLBYhr7o5W/AwSL7zN0onOkOb/8bcTiLrZwTG1P0P++10vIpPZVtj3KpUQicWDq
3eZepRr0/CycN7bk+RQ4B7XiSGjv9JtG4GLAWAQr5tmBJVhMPFF14mPz+2Shy/LUVbfUqNkKtZUb
P7NmdjsoLCSYzWX6fySMogx/cwFqAn09DrzMbBNN3Yb+NTFCM2RbT8YjS7DtkA+X3hzZQXRx3Yci
U7fRpl5cXcIzn+0wFsU7gi3tZzunvNyT6V3qdGrH/ex/j3pqmmXhPBv7XpK2zVicD0uLCuHvcNZ1
41q1KYSF4a9T3LY5G4ZpH6MGtgsSWHvCVcVD6JC/Ti9SGNb+ZVR0CsHgOL8VHsBX1Fxmw7Vi/2vj
cko+7FJV6EuUvOXDBv6RO/wNg3dFKKW9B90n8aPY0jjUT6oMhM6XCIC9HA2tC3WV1bOgWenG097P
zG038HKxKLXvPkM95KUpeGx4KR+dNzXtf0EJUADoCBLcIJwKnPMiBG5I0HjmJ3+Hp1LtZ6tDf1G4
6gS5OO4u8sdPC4wdGS6/KhLJw9qCYFtLhvVuXSvKng5bAwd0yVhEnCdvBaSIO/VJEP+H9fy96E2G
aezX4MLHNBwLHosPSg/DCGmox6P/gSSzgmatPctRHQE+76sAr3ZNk9hGiRbPpqRZw6gxgGX8B71/
ESiRbyRrYB33vhfiHDjdR7y3RakoKsyBOzuLmh5iK0NlqfbmjTh5HTMY/ZihhmXoaZU4x3cE1111
E/4j4RGnBadrV+jSv8Gphglf1wIv9Wjg/8trBqkZqnLrUtGzwL0RF0nLNgqT7rMzhaBsMWowauvu
9fAZTJwZn2exK2VSMM1Ju7v056VbBN1HRRX0sNGfUuQMIlpIwDMgapVz6ewv50ant09nSN70Nx41
EaqiOinMtlc6fg+4gaLzq+9yJTUXT5Yl0ffEyvxWpnMsjSGtYFXNDShLEnlDqE5UcCfkfXIb5KYB
iknF4k5hk560v6qyGE9mmcGoCjvqm7mDG2PTYikAlJZkX+Rq1HhuuKBRlzji8g3b2EVZycx6Bk4n
Qbw5jsJSO5pIGwVu/NVcqYU7bm2u0Z7CIld20jG0eIF+JbNpNWc86UaxGEfpqDlLgcK0jkmSUZ3t
rMda1qfuXjWoIXARwvsvq2NNdao3ppUJtntXePSOm/1PEkp2a0GgQsebKtCidWEG8NNO+lhmdRGi
YkdbCWYoiTzUlKB52UKrep09g87G32N15eai+7D7/r1/MRWjG7CcCSpSeN8c5QR4jrncbBmOOZG1
COdFUZ+PTbpBtEcECpNie90EIn7kqFlsTKmAgGVnstb2/XAT99gDFfU1x5WQs0DaQcjL+1x5GD5W
Gb2aNuZ9xTUNZW5MAChKiQGAZFxpN4F41+t5qND/7vc58frNTpzSrAhMwl6RaiXSivjzRYydGZuw
omXDzzUvNVIUCCxlAPSIyx6DHXDbkaEjLJjYDqFmSSvCn7aBPFlJ7zUTQjZfGfORwYnPzYxW86AF
lnxraCo7dTCLLlwzK1Vat67EnlN85RqaNBk9dgixjuiAfq60vqwBQpAloHgkLnkDxqpj4lqGRDkx
KsbZQncN3K1Ieo33nk1LO9GN+aqCzhPKvoY9fCY4BkukZ0gWWGmjeYbPMSCrXXK4WWPenEfGbcQn
1SNo0nwce9EyrU5HNE6cpKk46iHxPj1V9wU0QL0TJHwBgBTSFPP2E0unavt84W6wH1mTpmkCf2ki
N29icTEUNrA/8PO4cQ6n6jznJ12DaG4mZdn0+MPvYSxWmp7EhtrNWVBDUxMc79CMmc+oYCtrFL59
XfFXwnEBImIGAasoPKnZzTRUh+2UJYsNCJUekeWh2uYqCMoBLcjW2nLusHpvpA1EkfX6SyVaVTSe
nunLr5rPChRLPcBOBA8CToCfH72NxWKY90v0M5GyCkbIQR5Nd/gt860gYdv4aW9ggkV4USkrcVE5
wLySBqvY/h482qf4zUxwe09gdqBxDZv15Yn8gPhK46vDYkFGxeY9afTgxmB68GDpoTBqJ2z/2NER
cjD/cPP3g3lWRKnvMpIPwj7IvjSh/3sTZefNl187wJuevhlGiYfrUZKeoDWB6dIduvXOz4JC844Z
MNKTf6CGi95xK9qGjUx+SxTtzkr4YqlldYmYz/OOwZl91oeZ8ij65kzJIoOrD+HEmBUzlNidTtQJ
NJ0yzJy7uEh1VgAtfpUBzEgfOkj/Y16OwjXBO5Pd+YTFxTLo2szF1OxEAgz9M3Qa27yTti8S19JW
j9IHrvAfhiL+gIqfDdMom5W0qByqaaxKjskaPDxr7i7ddZbyQ5YfVvm4qMYuVKtUVkbrowohQtw+
+XjGLzbGSUhkPlMB/uE6C2+fatl5DhUnBpOApOb7Q+8rSQabJTVTHRlCZUpLMFXig5o5mcZtH7On
gwzzR0nPklvAEsF6sFQYjs34vPll23mwp/AZh132fcKkb6nt4ESSu77y4abLdy45UIUjiwo5uwRV
uls2yhACY3bO9vnYoaV9uEe8eYzlcpYMdKE9kZgw6HMPv5KgtSPpEVEQA6T/QuSKhSMuEVs6Kq0G
GOz5VyE+uiffgXSC+MIVYqd2HAjKo4TXUs4riduNpzr78tsKqiN4QlQ0gS1iHtaKsm0eh3CdHeGP
Ld0bZz7cxHZJktmQKMZjXwe+NiuBkcX8Z9dHmOQNMgAc0kjullIBFhkzVPZ9H6WsxhJG+7+8dLeT
hNM6ugaB2tKb+iehEjrZFD6Vt047Z20SP8Xc2j1+KThBFGXltAMcp2O36O9FJ+SS9VBAs3UfHpAH
fNWY0kCi0Rq+/JGnUPiihPOWYmdJCfVrwrRX+UWdBLHD2uyEWRzgpyVAcfMqZWcslBXFMIHvr5Bc
X/p4Z7kkVz9AM0iC7H1YBXEY1mj4BGd/+M7hpPuRlptyu0FqK5Du8WYmUGwu+eVcmLVqf3hjLKqa
G5kD269A74oRmqgwXVjPZ4CSb0rGpjIHAjcB3WI9gT63QLr0O8UNimyyMwc8bQxcDLKpMuriMM9K
uldhEB+SzyLFFAxQvU2M08Q/JOr3R+ESOZNWLEWVDavgmwPeX9RNKI5NlqjyMpCAv/Aq0GoIHgnV
68xYzxIimmOohCSbpcYY6fsRoM2RbgRj9QBs/Dpm1cxjdsLRWU4SYO8UQYCYFJTdhaOBRp1byJOK
KzIs9ysD41G0gzFHyFNdIJXhicOPkITLEqkZmjqyE5Za3mcbgRD4Dh4z6UShLOaJa0d+lSDFrpbr
Y/aNoABY6J/H8RUd79gntKD9aDDVliggm3mZk0SC+gbk+wrCH3aIvOI7kuGi4fMfEWrGm02mB2ug
0oO9nrp2koq3Ey7xjEJF7nVhNuW6jwTNkqxHSaC3eg24hAS+jFzqneOGci4hkcC73bv/Ba7mygTt
uFrw7c15rFpNx+LhGG9L385pIpUxeN8TUK75s5p/0oaU+qKdjQoSScc2+m5hI9PVkrTMA51gKlXV
nEE8NqTymt+Q9ba4x1vXnu7+xfKyMuWC7zKPt5pjBJgEAV2dqUIVpInRgp3DMpGFIX+ksM0r0xEx
TebXB6RClPbSUP4CHhvDsINJwSto7IEAEkvjhgZTVJkmAdhG2gG26/wMX1oq1xhmeDlk267wV+8T
CVPJeEYkZZFcbGBzzRfm4mgyH1zOjMog4Zf7y/1cCqq5t+xiXv7B9maLxWiFX/yLwXg2Rd9St/YH
gNgE11LmuAoQFKHcn+uNzssQSUgOm5nXRo277ATqqhd3ptncnNAcmrb98MG++7wxdWf8f0Z+yJmr
UulBh0WHFb1piB2dQ3PstFGVLyK/myovbj5nSdCUAl5ZQa5Z53BJj2Bec1tNJuTt1XGS6x+m1bJb
gLK8zL+oozIBZhqd/HUelbs92EU88WGs6DpaIhdi85tTyG3bvbrPHDmzlWTie8M/GeZ3gckkiPUL
qmkUUvH4t48Ntq8DQLByL0OViIy7W5lk2PkcDnNQ5pyTZfJbNHgF8LgXxziTTHxl01KZbOsGw1ax
0KIzlKChH/vzlwalDNWMnWdoH8AF4zPueKZBFJgkvzXNkXnqMmxvwOa4+QX/k7HRpMQqgzFm+Yqb
WctMYOH/cNk3eterOSp4HVtj5IxMOmL0Wetn5JFpOj79wBSlQAzgsSuGRzreHBUo4aqTk4yt6TCm
QWCAzmXWnGmkD5rbazTCwqvWasaWNyxajhhITBO+j3TsaxGk/IhhglqgQOmRKuKYLdohnijE3EmL
e/ScWY4DbhRtEB/MhCL7mu/+TVSxUSTM3POxymrOMiEDUL+mtBykw4wjyzo7KfBAVl/qrxHCh9MH
kse4p6w9MQXmBoMq6voOF1/7wbmX8f+uxQy2zxICqD1qIIfdNUmf8GQNx/b8xE0+wP/Wzud843gp
SLMJVsdd4G9T0LbkHZc/uYOz969atcHb3cUXAN9ndj8ln5q6LIdrfVPtuwC2VrHTGA9rScTJ8C/C
vMvzhQ5CAmnBr9jBGSzUWGeQWMMyNOCkYE6fLKx2AL32DMpHhMckdSEZOp5Qh/Rfc0sHmVXlIFWa
A7IrykB5RM4t+94FrJ6ed9ndQQNjXO9ut1bXlVpaJlJwdeBMJ72XdUH8h8gHZZCUCHFCCehuswKW
q0+8n6Dd723AVNr522qWZ/7jhZpmGzEGN8iz1XaAR5dwpHKnMLyDIziDTuNrVmMU/J3jZvKZvF5c
8VhQ42DYZ5nnY4TUIXEl3ZKpGRcNwscU56CBCQmGtgGbtBl+8U4S5bayS4D3/tOo3Ny+UBX3LLvJ
PDHyIAHEIouGywiyrozRlHb+jP+D1nPYcU4LarWPDPHdJE5BSdtpkFV/jS/Mw0i03stFtBZ2UZqp
ZwyeeB6l3VMrsWlAxWpxwgGHCqhH70ufFm6sWSTuiI/OThZLqqBDVytW+cX3GdkzePEa5G+ofpEe
CeklgTdC8yxOzVIZToMYCYLMCeRZ4Kx7VQbZGuu0wB36fbRix2nnUuu9B2Ndm2vAQtvQ2TUlD5RV
WX8br6YNSBEtfi/v0e3J5rnUJGs23l+2htg+y/L4RuETEZqPhaEelAadeiSiomLj6tDX06T0Jhn4
purgrtpzlFe4MYcPy9jIlbE8qQZeWZBSd4PKLRAN90E7ERvXkHWHzcPvwvMDAJ6tiWx21Fy4uxww
ASfKoXPLQ0p5/oi8Bap/zAF8qplOkfDGuKO6bcjB1x+9V6WgHqmaMVPL5LspyUssk5MiujAK2Xhy
lnUX6i5IAsodYQ1o/FFcEnKS7gejstU0JrIBIcv1ULEB2jy4LjVjhXdbD2vmbhkXtQi0q2jA6fC2
jwwxx8WkUqqY84F5zehHFv7ggVOYS3tLJ0qvQKbg35CrOrLmnNpVpIare6wTkfV8SMPJ16uFhBWT
ZIq+0JA4/H/hcIyJWwkVu96dvHAcJ6KvNzxEsAX2XLX0U8ELISaywG96177+peCehzTswhP2cksj
JRdVARUjY7gtqrtpO7is1fOsFbj0rJcbV1LSJhx7C/3jjfIHxxmno2DuY+WTi0+d64Dnn7D616yI
+QkkWFgrAr8TUepa3FwGDr/QlJufRtaBp28+81Ocnyu4xzCPnONlHJHXMHlEa0iSSIfR3MBFr/Kr
qh3meVv1IKizgS6STe0zAAdk9zXU5Ci5rZ+MGomePyPtSprTNQDbGe+yIbhDRxs1u6pnM/AzBQhj
DVLXDZQ3ULT0L1cDEY34oACgkrJUB/cXM/k1fpN79eShbgGsUSqQBM7sTbp6cHo0x+ojMPVidHkZ
G/mYP1wSZspLUuhDnXI4WBz+Zv9MDzvkkO7qfB+A6IvueZNe7nh6ANdylZK5rnpeUAQOfjllawCF
/9BhxPxwmRa6Njd7JgKe42Vbc3ck0BktOlulTGqOr672JhDINhrpvRaa+8elrQmp7j22EkQ2mTTA
Lz6IePy/vVhNLxJNk04O9QY+Dgx+btCD6IvONNxHQtpZZ5fnkGvYEYNYt7wqX0M5tzxRlwmBNYYi
J0xNV5cMkFPKItp/DiB5oJKZpxML3vtR6qsVI8yCnubytQhYq2wim5BOjnuJnoNaWTHHv7RTg7k4
XYNZYvxCnjGNvfgZTHq6uh81qwgrXKlTIqE8BoUY4d3DH/R6l7zw2XQJkDAD1zGzLtX7i40CbYh1
IeO3Qu68XlvN5SFtvxt+2qgJnjblpcsiW6eTJr+5JyS9MPhq5/fciDein9/QqVaDRqCTdYYwKSBB
IDmuxDZYg3ZlfvLIaekkBuDZ67KPZy0wayHpVUJUVDhY/rt9RfU6Ui6zEIxm9yIRESLA50QYFysJ
OYmD3Qd5ELfCkxDh+XG/JIsYkS7Lq82CZ0cf4FuwvudGkX7x6IA3MDE2ezlofYoHQcDzFQa0X0+w
rg5G5DrZyAb+fY56knxU9AH6RiUkoldBZvLnnn15Ap0tJgj3XgkqMmqwH99PKHfjikqoyORB/Yqy
oRNbIdFt9jz0onWCCDOPSSncjsfY8zUfrFaiEYL7nt7MJ0snmLrNEI7n2dJga5+7PJ0H12g29vmU
NX8ww+/a+fMwsmarKg7uroI2U4au10gfqSeFimgCt3pfMqL6Ii39JF5HZv1V+twyu+6GGFtuZJhj
hYZDhxfJkAuxDd1bypGOS/7D10ye88wj82QvgCErngFMPFhDQA1aixjGDsqdBqXRGQshohtwOnzP
xlTiC4iBYZjbZ98S4sPHoS8Zx5Suyn8Kv74uEEKrKxrdj0/qMz8J68gKabCjUZgFXfBN6zCfevj2
6lTnaDwBdVEzMjofscA0q/Sn+QbVuQSgu3GVwDYnOs3I4LW2o4dc6boIFZ7bw/Tc1FgqXQ3CM16D
CmTECQ8u8GjXI5LEewGCImQtnOfTyUj2dALDNzwUUTKYAL0KrdtpLLXNJCGkE9rbFusyNk/BguE0
JBlNk0m8Yn43xDsMR0QAy8Zrmk18lNLqKE9f9kfkULFiC9iDPn3j4zuaLkiHOWE1/oGcKsWMTfEP
yEQU9Hh0yGShRLCDVA4C0Mw81xi0Wj4STCXM6B5rifXyv8Am35hW/Z84Brau+RZbrOnLzYe42ScN
LUK7NG274pKWeuQ8XlpeHIT6mOC7N2v23cgGschb9jwILqpnEZ9+my6iYA00jflASStIhscQjgA0
i0exJl2KRtUtsdDivgx17rLEF/+IXH34UlWQTU91xxl0cJkBTd0pyl7tVAnWxVZl8wv0iGzOH04/
SGPsjhaFlN9kstDzR9HAxNpCMIGIm1EYsGPXGncVsCYcEeseNZCnWFKwJN/dpS+k94JBoJhwN66k
eLtvJf916bV3N3v7Trsa1D6QPcKQFA/6/evLkQCyKEktEQdSPniKwPDRJ3U63XmKrZ5mW0uH4ad2
1ougMO3bszh0mos73Le4lr17RRucgGcTr8QKa+WSM8qcV+gMWMmOLoa/V/VsJCmg0XxJGSO7BqJX
LwyiNsSqZMvN0/x0YrOrZXh9+9lBABm6Kh/UmQXMUOVlbr1q0LZ8qfTOqeW4xbtU82iCMwT1Kq2r
JU7rYCx+8FpqyZhV4Nl8BzCNTvQZfR67RLL9Id1+2OpHp4d62AhX+I/H4CcY1lC7y0RZJGy9td5T
bzxP6gGiqidJo0x/5pM7fdOUyrjTaQ2GKTacOPkiHj61iE3sQr9O2CSJE2zBQSIbYkQNy4Brx2X5
DibWPU/dU9SkdC7HYvyYLi+SWLXVGpvqzpHvZ7ocRDG448suz4E4ElWKuDQmt6BMUC2aCiq5qgbE
eynS/xsd+jvsAp2G0DqFAamYNSrlg16c9og2dPxxJFGM8GBHzLGRQhzaVtCYkSrzBikdJQkSKXkY
JLjXAS34uAaccp7ASDTr+EnwZpLYr3iTdfS0yiHX3u7o/3laGknnBuo39qo8fIndNSEtAD1PFbMh
7tOaBZ/ZtQGgATXEJa3zf5AaYhOMKLthl/w5FNHfYOHduxFhrMrYeL37xrV97ehcNvB+JEJnLIp8
1Cm/p9uHNv3YjlwZiLwe8YJTt/sFKh4PGi5TPwlg7jD9M6KsiBfLJG3ZY7l2mX7uvffIbDlj1O32
9KokzRr6q6Ey2GXLWnYKK2VFVV6UvcHgmZlm6K9qOTaclvyxmjS+JrlxFok38gmFwYkui8zjVvMV
q9p7iwDyvV0MOtVSTFeIUKiDUz3GmVNiLzDA7bURri3V1h5XRXwJ3kkfa4jI9jsw8zf//U8dJvqf
L7mtXwVQWzseDhTlxMz9Ncv9OG63eHT3RYyMf34CzPDu6W4E8csLTv0GqRCTTvqIIy4sWS8SzC/g
45tjlTLtfiT8VA5k59BNgsfdFpjoBO2aCdvpyHra8FlmX3Idpj6WejsMqgfE0PzZY02pTWgRPhqj
eVnEMBPsBKsuxkWy6lgQaoPg5e/CSjP5hVJ8O0qk+uQ9U8w+3LFU4O30XgRmR+0nDVIIsRGt+HBl
GM3MTjSFrC33fuHapZkpvHOQAkXEN2BjG2N+AEzPOWmsojouIu98FheHSEUyYt9wXrqLXjE5QSWS
Xmy0AgVpX/rDj9cNQBCJcYnGUUn02UMPCEuVHiL8hU8yWyygq9oWkLsOqVhuNRMAWqG7ZZSfWKqL
lma4fDINqVrXNugSdCks5jQ52Tkek0ddkBU64VNAKbPb0IgOyWg/U6VLZPAYN1a19jJHdzSIvuIb
M9vDXRyeeOM4H7lAjqvFS3U+MtA2dSI8Msa4WzfaxiDFWWt8EfrUddbBYDjRdwNNCd1df1jCH34Y
uF05KfZsMpbK7aPhQ8LIYDq3z1EWXTJc3Y6Y3T9cd1mk9wYOH3yAmCWw5yYewcp0yUg2mB0xj7a0
LdKV5tQZHd5DfjZnDwM5uDwZ7Cepg089B83uz8AtjwLyE3I7MYAY1qFJanlChjMzYFnF4VIOFscM
LTOEVzJvS08GH7Yh4p9FFcGJQWI3WlPpj03dpxn80aHxxSNqfZJcIDZc86Qo/8++0MrFtW4yPwii
zEMqPQ/Ew62oMPOZSlbd9EInQZ23ixbtgxm/FtEPV7bRwFPRuyFKVlBY1CeJUEKGAH2mR5MNyH1W
5LVv0IRdHK8nsgOcM1NYdvuA8keNJDfpJrjMPqXP1fh7u0+uncss269n4tugLpTkRYgzGCuwffR5
FD/p0Z0EjuYuhtY2eKbXIMGTCm/X2QL1eyUEnX5jmdg1137amHCs/vGuFZJp0BVVZBsiljLOdfc1
g5Mj9seI7E5dBr1yzJaLePd623vVBqFpQkS6KdjlIA0WvPLW96/aAlibtoJ4YELQfPooHJX5FIs9
ClUvvENjCy6zkkcmt4+ToJXF+49GDjdUAc6TafV9vGj0WiJWYAZdZjoh8kqFbVrNUs5HEjIQyzL7
AS+Kk7QoWzG760fhT/hD+45naz60utfBQpBCePlrVUEGIxsSSdD7J0FBKZM7e/LwS6d8Y67w/BFt
SiFYeO7O/N9DyWVijgbBghKlVTNyd/IGU1SE0nTxWCJtz/Ax52qLoclBCtOZ0cmBaP9emCEtsmBF
J9mwDrhbnMUwlAdsdDz7EEvt5hM6ASGTiPeXuAXCwQLQ4A/5RhNdSw2wiYcs0sHHjyvEfgyri9sF
1MFJI+Np1fU9ciBnllQwIhwhtjXrdzmrH4hjP4O1W5XY1mTBOEgDv610k046FHBXs44VBG7wZQFt
QdryDDPYkYp0Kc9CVdKk2YMrNd4Jfad79O36sxtnKKFoN28oADDbk7ATEjT7ld87xsWug3YVkgQR
vVfDdNDVJ1TkBNATtwg+mXegUhGkw5RbCdoo3Ikm68becIron59W2pgOgHNozHcxW5db8Ci1d2Kt
Z5Q8DpW45pj1n8LRPIG68ZHq4E8of3wGJTgHUxTJ/UOrkjVlEDI6u0SOJj6CWQmRvLDX0J2WbzLd
H0qUuoR8+ZD1/f1NVR17O+si6nXA2WEuHjrKYfuXWeEeg41fi7xAJVJ/fSB8qb7kSzqS7ufQ93Dh
ER5xl96Dir9sbNePbcSaQwgZc/ejr8O9fser5TxX73vrDL7nsG+CZh5/XA/YU8QOp9zWUaIqqUPI
3gXNDl8lp+4Y6iCfsLCulpNbY/rhwRtFF4Mj3Z+HB+fZ/yGc6BDjqvNS4Oyv/zGiTAy1Iryj7Lr6
dkhlO6NKnf3blme0CH5KJiuGuERXbEk6gFUYHkpH2aUt3IzYuSi9C6Cwd0AVGpG8QDVDcxxKyvIP
zVkqCmfnadBl/gXQeoinkdS0zmIGAIhtOVuHZC4FhIzTn0SnfGnwNN+WMRnpimPxDnCQft90wB8L
Su+X06to0PA2vdHwMcq6qRbuoiKgmvibsX3hThJQroRQkyan2rn8FVkf+fM+RCbX9Ipe6DnH2IBA
TaTzQGU29btkpmP/xihahq+8J1nJAw9ftoOwQ6XQ8K3kZ2/+RNxVue8qlmB52Ws3AWfcMnuFLFJh
JqgD/OonZtS7CM2Yex1IS07fYXhn6zPbfINhsRhTtnYX2j90UTQTNGHbXSIRwmgHgzkVd2AxZ/mo
yM4tNbcHQ+T9ONysO+CDc6W7ZTjuXOCQfijCkdkVuwCwGrq1o0RINAgnRyBLFwLi0q+WRA/SN3k6
opDFzbGbcOjUuwpRRNFemN14GD0I719TONlA8hANhXLcE0f8Y30oBnBIuUxtinlnICA9oZAUWMwN
2JVJOQePiJ6Z2ecPGIEjLudDYg6BuOX36khGKwf7N8UlCWwT28DZWWgdtPftdJCHSsxwKBX4J4HF
AFnASeBeQQF710zR7ZOQ/kaRv+4SgsnJGbzHQrrUxwsbJ5/SNAVjXMVSc8doqOqXREZEu37fup7V
mJMNcFlO/E+8TOWHpS5s7SI0rK4Ct0yvdSt99OYoswZFy/QTngACH4gKYFdU+KyccdsEcCNRvEgh
0n6XSjcKUjO6KvrIS+hy+//u4jG5dmuRmb8vqljOyQNY+gWqU4ipE+e8kp7wOw+c0qieqtNkLasG
gZCcAgbz+dBVxZKscZ0Dp87N4clmqMkH5fCbiTskHPfHP4LBjZB/D6EytSnKB+d+RRiv3iYtGFb/
IUuMXMaXu/OOpqzgCpd1u5u6cr6JKdREKUWQ6po1SfjBPNhunJ/lhovTL2nhMkJSoBkukqFEeAmW
qGcqtEQCDT+mAqpfd5QY58OI9Q0dAXNKQw0KWWZoLLXCvgCZAV4SOzNbpW5NFl3jghNgeDmWlhzJ
RNpsisrQlZmYlh6OjJvzFZXxkuAJsMRYq5p0Dv2s1VWBhi6BkYVd+oK87kjAA+QRqTxBY+uW/GY8
HWpDW71Lhihd/x04RQ1lRJSSiJekH8zYaSxjc7U9vWcXt2ifjVILak6DLfZ1OjtvZXFulTTrd4+9
1z1ZKa4x6W7c/hIj7gnM/0Me96nrOEya+3cy64k82mpX5LK3ufGIAcII+JTOQOBhYB6QaT8/+jcW
A5C6yyFwkqQ32hjkTn8Izlkyt3mPL6K+G40qiXinZR1hwwAwE615c+ly4qoV18TU7U0ibLcNNmsC
vfMVsvJdTKQvkEnLp3kIh7sDG/sny1lk7JirMVR/i+36erivalH0yiYhrkcHzFsO5dTaNZBPShYv
YT8MRsTkcLzZC2qNs3YwzK8bbzcT3BvZ2OA/DGoJleHGi0DT8cqz4De3L2ojXF29U5V9p4Be+kOS
cRrQ6mHtWvZmYGR10QTN4/vmkcWDxlaEJ39ll2BHuZjKHWxRo39m7V89RzuKmDeydBjRCvQwQiGd
DxhiYhTpaTYb48DiliC685X5D8hE5cPUEKcTVp7uHhYPAGARJZkBSZE9++S6YS+2FOeHLW0dmjzX
5cBueWQ6J1ndSWPwVIo89llDQm5W1LkkYhWh0A85Rr77oYb/x00K8dS/95jE4PvgQh0bu3Flkqpn
O2OwAPn+WZWjsiYTD6C29M7cLO1KW7glGFDvVVqMuCc9WMGgYU99UcyUWF6ssT1DEhdkWbu3VJLy
cjBxAwOiJ9Q7FPhVWTa+7SE0Va8vmiA1IcYnHHpZgN70Q4qReJAnqZk1xZ7vJraWJpjP04egncjl
pSPHpSRGD0PMZExM2bRHXLa/G7n9LZRi9vy4KBv+NyqlEbo7Gzmvgxqibz3uFcIBmnxd5sE0gR5y
72knCv/WoRCj2N1UtcDJuYVrLuu2IDPCc2BkMLoxUroCxKyINLok8XFrwN4LflZ1Sy7NDhDczNMF
VIpUCVLWWMY6rr8Fl7GFnpSOUTq8VXqPcD5myCIGFjzJ7IXpeMcyJlWON3k8VkczQ/14OTcdGBvm
O2ecisibcJCFgcjglnFPjiuFRv/2+7WjlUT62Lt//2KrM28E/S83WF1Tl0uACHgq9Oc2VwuuhIr5
laA8LKLsoR5XGZ+pHg7/DbEHlW7Ej00p3SfR/FnPQE+mHGQpkLt2jyJ2Bhi7fA7EjDwpYOYP7LCs
zKul1Swm08kXNHUUmady+jk0+CNBxnnh04uLethQijNfzoFX9bEWIZ6V9kWvQ/mFA8wffwR5Fpf0
mMquidOi6FL+8DaaEjP89GVjGhH1BXLKY4G91Dq0XsM48D//hIrOYYHz2Kxrry+bJgZsFbofFN/v
RzFFkLtHGEfXITXVhHsyWtbDvtau092Cplz9zf2CU46vDX0dlWSPjXRmsurTAnU1NSD5lPUizle3
wG1b7hKtxwuDTkItHuV6yLXuJEdKgsARO1CUNRWQylo2CUvEdG5SzLhj++PcbNIexBe5D6LcPfXu
maXVcwukUjA9VmvyC8w0ZgGR6+9CDpSil/MOsskpYfSueBL4UnylzdnbpGQ+HpQ4kuU8BQmn1cnw
vdtKdVxYwvyDdoviQRAPDRa/M2ZaNVwIEhD+Gzt260DYwhpxGR1JFvPeS2IwGmwPT5+ZofK+/lKq
w2pHNicoN8RSMlY2Ns6sI5DSNXIx7crLo5gPr2EV74StZl1Z2VS+wno9E01sXXB2ei46JgoPmQvk
GjkNJEGGdxSxpD3JV1SAUzTbcTtXGbGPUwJhxqkigfDwq8QhwwShDXG5pm6G3SeWzpwImCww5FwJ
v1Y4zTptB68NzSBaXbYz5pLSKyt+Yprh4TbATN6ZzM4AXNHmEydKdmLEUob1gfnfYfwGmxofFaM/
/fxyB/Nl/hYJSDKSm56bfmbpYO/Dn7z5HHtQEFH8ZJFnGAq3889Y4vuZJjQnDX8h0ppVcr1eFSMh
R8SxKn2NOqKo8Y9M78L17A41+IJwugaxCqWbVrHBGZzMSXASH9yYvzKHbR00MkstJES+tH7qiIV8
WWgcE7QTQJkFcG5J7BKQLlv6FmMZ8JR/LthBIZZdrfSLfcIe9p7dh1puxwSaRsAWloDsidn9C1NV
u3B9d1J9DB5E1Eprpq/jna/4K+wq4wF7H+RKpx0l2hqwWItROZ28c402hCgCindSTLdaIZnCT5Zd
ouU6TW4I3hQlcc4o/X0g+gB1iJLMQ/UfBU43hoM5sDdfgI0hZsNCdOIwyEiMf0Q2hcD4RnHPa5FW
UuKcYvx4h18Qklm3wSsEKy6IRXDlT9DN6ElmQAf6K/n5+3PNtqG8EqNt1WCAfOEGnMA3EW8XbPCd
oM3U1Gc2dEHlClTR8wLet5exc32KEN2zvUuK0+FlJFGsG2GdDjnUpmrDtjOOySKE6KUjeSeY3AvV
ntgkqATuVpYafY8BX/z7o4D47p7HQWqFxD9ihFD4w7hDcetPuqEPWOpsukn1m0GmnrpCd1mNdS2s
/WmxN/SWeqKPB3GKVU4dSfZD/62lnHN1dGvShe4KlUWwCYKdC+ZbvG3Ak0R5+DgOYxYHBVs8bJyI
A+PJcF55z9jT7likArlmy7UvX+5CigEV6yg1+0OWGPQhI2oFESK9LwSDGznTFYi4XU+8mmTmMv8w
LfQB5IbgJ1CQGH4iMHXnDuWgMV9nlrV1a/xxzWu/VyK97z8OB+s4Y/T/lItXddtbqAAd7o2fL2fk
R3Q6jGK0WYnjO/bCTWBDa7i7hj4to7uJvQf3EUcNyHSXbwVMXYkxmRIjWM2xekv3q8OoZ7V4JleV
atjuVIq+C4UwO5n+Qn0tYFbS3cagIBtEd0njvOWt1QJHySVv22RALTM9PzG+u7GNe8AmgNUZnGU+
Vm3qhQyK/1RWRiqgUBoMek6p+jRJuESM/PnJlA3MUoFEYiCIfhvcsywtwGBzMNYfnLaVgnKUMk+7
uyYjeT0f2/XOPuw6wGACs3lZb1BXDB9T0sLwxToIuVhfQE0jIC4Yky0QbDqxZAEXCUKqPjoNDpUf
OeVeu8TSUwUSd8kHxEzslAankYfNwTQquIPx5zntTNzc+J54hQZP3TwwQ6W0x7TIqFKZ5ByCl74I
f81hSzb6KHfWnydp0zoXfyirZuuIyB3+JPQxPtZc+zZ/gAC7gHVJNosn5OYgVnwViGwfiEamN3mz
IE7YfTP4CUCp3V5WeHIU8cCaS7BTijE++Ok/XrSAnxTDYqEqB32Cg1xyou0gahetAvVgvDpDWfE+
HneNOBU9rNxDPmGHV/kV8P3gY3UKHI2yiuGbQz9oe33YlqNv84jFLOxitAMLILx/VPgtykCk3EEe
j1vLh9rZhJWpoMi3PqkPsGjIBvuqoX977ZWHrnSrkHZ09ZNTDHpy/4+W5GJrQ0HRT046lS0ceIcc
RHavQc/+jsVT8Rrg7Xne0m06ktFn5HLcxbjIDIrCIw3kUgJ2labbqfhuiMjQlRHeWTf/L8g6zrQL
tmPaxQ8q7OZvICWatHCDiOiVqvIKDy3XalWonlkkCT0qaZpKmm0FqTehT5sq7KORUOg7OQVUTY8r
/0ayDYE0BLA4g8C0/+fVCitToadSOZRs7DzO6HqNiQiN8L1nTCjaWK5e6qRVi+VSRHBU3DZ10m0C
eC2Mwv5tccxON6qoKK7mMyGKO1WntraiHxlv8k/PUeFGcHDU0KDzw52XzrW9LIlMGtqq3BMgZzmg
yFZW2kpi5AvFNNNT+gtYzlnJahh5jgbdhCpgeJu253sODfnIB4hmDGhldWpaq1zhLsfw7bHngxDW
H5i2kNtk7k65gwXzC/wLL9oyUpXRzgpNxFqIleVzhc5ZE/5yvo01xe84t44BUdT08eIkLiYa3h+H
XBTI09VnsYAfPubg+1Syrt7PTNhPZWJj2lc6i5lYWk5kbPn7REp766MJewnDSS3Qi0qOBKgOnjkH
1lHEcbINjStHtUZIhexYOxUthAxCWM1zasZIf1TveClyQ6ViYQJIclzBFhH0vn57RzHX0FNB+1Nm
gaoaJs+wEALygo2iHXlTbIt6590dS3MyskvJqoMS/s/DZyj0Vo9ADXS2eLupeKI/Vfjg0U92Na+0
/A4/yviz7+WtnWV/2s9rD6d1XDqUm2iAOAeOtgPHcGfr1/MyM2TExxmgqUMo75/M8JQbr8fs9Ozp
1bBiBA/RdTZb+Wh08ZhmeHaW2JIayQEL1j5MF9+3UPZYyUic2wPOcG69XZgv4nRQb1Rk8xs/rkeJ
Q/tkLG+jskOH/AObxt6yX80D7+vpGayaRObyyQpKhOt0+kySXv1o15aZ5ljPVjv6ILr6DjuG+lJe
sr4lT9mSqG5pDMrv679ulkTmiY/VvRlAUz2gRx5tsRp5lAiEF7HaoL3pgEILOeXehDLkzjecZeJg
snZhfCB0AztHPyr3l8Hec9pmfFi8FblqIaketA4bkZixISq8UnAfNfHGUNheesr4I8VswqEzyXxn
XGxURYCK9f4xJc6i5SAGT2dCPS2MRz2Y+EtsBGagDC60t4aLaJPNTXV5FwMjrVaIhnW0LnChEX2F
c0PPVMOmLAPatKjksaSxHbdDmOkT0Yu2XmWXu1EDLm4zosJLa+Xr2TGon0YNpM50HkZIZd1NkEFH
VNjaiVVjCr4dyQ/dBJ5Vw+Lb8W4sw+zIvx0b0G7u3+Q2f8GkzPqtlevkwAdB1DWfkzScelJYxvpr
Pzj0XZylWhd1UIDoSV8CombhJ5Xc9EAp//IWcpv+LnJqNvsgSRM3NAhsvQH+8Wx/J/E0y9lISIug
YMz18QV08qCgVNESwjybh6r8Z/7nSJ9eoLylqoKZBAWM2Fv1Nz6qboHa54TOqge1STbCZfwsLu4/
fcnGbI5gkcANAu0XrA68lgSZjuqpBg1iK3ArLWvKjzMJOt3aE0dbIyfxPqdnqVIUiyDbI2tiAg8/
H+z5S7XoLxZKBWHEYkk8alw03LnC/6qjwQnE+YUGe3NgDpltYHtJZThEGZDS0QrNvCPUMVpBT0SY
aq1NEy3u25yL9wmUMa+sMDzxYYNvVXy6pDIpgrdiCVapXqCQgcnjA9NDTiCgA2BaUyXCgpEUkVkp
ST5x/0ndnC7MYFMEXYBVAXKSngZX3BJXLPHvKgp54rpvWiVELcXpzi1E3ZyDN+xGIpgIovxmjXw5
P5YsLeQvikdHRzRw1A2rSVjDb3Kx+OUxoJIgnRH1B4pkj9RKvafmd4ehNrzXuXFppNK6s6UA2P6+
vWM5LtAliRn8Aobny6pNdzUDuQQcdehvgj1cHzG2pFivRYHKhkZcezv97MSqWpFUljPQycbBrKTO
L2MjEV/LhXKmI8qSwNLUX9QFUWLBNBADFEnSJZ4+4i4RB3lCV8lfw/LltGWslJuXjetFi5dnHgO7
apE1z8wQSVgoMWzY587qs6FIKAIIdZxqjzY1YjUQgCp872VNVfq2BQbTIgbvYtFd2fFyEcd1b8Pm
QLRsxOOLVWgnxddRl4slBymxFVNru5LecjQd8Q0LD5rSOI3mUpjRlImyzVIktvwyzJGdZ4+u6o2t
qW0kloHrEgY6y5o0dspEcJ0+d0sXte78z42EWtW6CIWO3wZh0nuqHGco6aYRQ505XKIE2MXeKdDX
VUeGO0Vcp8XfY+KqUwp2zV5hXxTohP52rv3ufovLaQJQta8zkmLuTgr5lNi8vu4PRRjfYr36ez32
Onpzfdoau0Q7HwzOCHyjQpTL/yeC1ZgWc57Oa/d/82tRXwkRarvXTiYt952qhNdVcuNkang57qLu
Qf40MQuP2DhCNtm1ITJCPmMJuS2PtSqr7B0pn1oPB/DkkzxZj693MwDXvH7TjjlesmJfoCKJhFF5
6wISuYQA56mnRpwXzeevSP5yKSOgJv4IGo64LuJqgxKP0psi8qZ4phB9j91u4tUdMGQAydT/yF0D
Qenw/wERwonFjdbXrUYL+qXWv7OEGTVnP6LsDYutvIex+zQiIofvKNtyvFTDWkqaMmNYqOOCBgGk
eaV9UMWlKMlnoPXIgX4IjqnnDK6fUpxFp0WPd3BI7yqr083KTWalyPAJm3ybeIy4gnLZ4u9AUbgi
sWEfKdEUHFCpo2fCNnEjUvtpItahzF5t+8KGoO5fadn7kV/q5TzAixk9ecWQOR0FvzDCJhFso0lP
5F4wk4r35tKRm4oZQpAwTHXo1ibndTgzA1bqhyTYrm7De1w90xHYiy9pNFVyKZt5NWLNwMQJyabS
4uyQumGEGp/Zka7l46Cbtvl2mCCvVw4gqotcjZXZekyX8v5x8BlZANbBKIlEVoRVqsx/wZHkqj2U
/5uFAU1IZViqQke8ghGbc8chN3/Kn3U2oTla2K1jPvwgEvqQRHP6hP1ZFWWVjhCLkoGsC3AoQzLx
NipSkDoVquxBdcHxONFIjfjQevVfECL3TUaf955S5D1yzZSX/8mSytDVVy4cgdquqxt7Jl36dE1U
MRPac/6A1eCl9vogUideZYGwGJFyWAgaXSfvPkC6LU9I3AyPW8/DjQOlXeYFURoiJ5n+i6c+JYlN
MzXa25rRw+Wzmb7L11kamCUSaGbGeSXv/CmJnJgtR0l6yinDRz00i1XCWZugSc1P47Tf6EjNFThr
UEGS0TPsT2OTomvppy0+4GdWXpH/z3Y1LU9kIfpFzNTEQMFXo8zrxsfYnL1S3UwWx08EawBQxqmg
pKqm+RwpfJobjQapA1NY06pDLHI4ST+b4kuC8wWHhaG0JEvdK2OcGr7mVeC4UT9LLKY3Fw6FjhoI
cyM2gTb/zVh00IdK7ClRlQ2ijlqWIT1TLUyGeN/c4GBd8tDhJc/Fdpo4Sf8mJlwiSCAeuFf6o+wl
lVqAz2BIL3vEj4tjPhe5nJukbcr1OqV9eOWiFRA8fBbAU2Yq2cPC9/dqXXVQmAPbxnbZZ82h/qH+
e+yeD0Xs2U4jI/BCbkUo26GrsNz6pwkNO1pGuPGvD0YJRVG4spRuZgVzV9csUI3gsN65Ok4TiA0A
ikyuG34deWsLNmaHNO8ixsqBQWME3FQq9Cq5Qw17DvCxlx/RvpaIfxFCd2iq9fVtq+u9pCaRPeZ+
OrWPM7IEDNq2EeDOzg7OdfsF830SZWLT0wWKLk4TTBdpjEgyZMXtXVx0zH+ouAxTo+ps+VjNNIE6
TLuxPHIn9WXWglJd3G2bASxKOd9fA3sKwJDx+RB3b4Oqj/KFTn0U3ALjnIlGhsW9swaF4p62HtOj
TwPDJZhOSiY6DI2hkXsB0WRbV5IPX7ijSEmv99o9EUNlj5XCx9v7jg1DhweCqfcc4e0/rwpcZqCT
kGL8A+r5xLnb56qe4ZPSP3ou3kKKMCOC0r8u1JKj2ny0MruyuHVIKmd93WxorLWpHbGaezRNRe4O
6O4M6oCBXmByuu37KuqtxriBZAN0nY2wPtJiMoEc5Z/o9RMyFgCKI2SLnxZlzpfQMfg/uk00LX+2
t3DBOjY4eg2jJula/CeL0+b7hXSLyk+KZQ5UL11F9ffYdydUcloaJBi5PRnz5x1d8tGV8g8ZdU5b
F9X4BbsdzhsSZOqW+FV5eu3+T5hIgGPZv3lyQpp6qrEYaHU8s5Bav+AaUCosRhydxb8QxFpgBpkk
3TtBKv+zFlsJceqV8+mz3WkhEX0X0OyYW8ZXYlemJzMNDQU2+Nna4IEJYpryHMLqBmd9gdLeND1s
wOvxxI4Ly1qeSXk4xuSJyaUJx9nVafVRBhMchCwVSdZn+ofu5lL/jsBaAC3f6yIYYhMy2BQDuXjU
VBmXXcEeeWGEAh80V0qiFJfz99e5nZ/V3qHJqmYqbkh/xYEr19SCRl9b9dSrWTwvPehgXJyIm3Zl
K0ESF62vvw1mm8GKjpgwegVql+bsz/3HVfuu+8yDsSukg8SVy8vJ8DDjdpMMEAGHvk3aCLEAMMeh
A5DAKLEhdYUJtQqVdgRvXld17Xg/tfrKp3UZrJ02oD/I5lK+37pCCDbO+LETtZxnfa9UfDfKdswX
HP1Y+4pKBdY0C7KxHwKFInvjL5xwP3NA8X4KG6YLDdPcOeP99EZAe4n+KZePopv4ir8z6n1SsPVg
1gHLpCrYUaQeemBp7xI/UJ3RkO9MJZB0lQQlNl1acXop1hkbBPw3YeLVYdgPNLw3e3vD3J9Am8fH
Bu633lTwZt/oEK492N/OrVCbO19/H3BzEVJV28/O7+F2jBYS+qDvD+jWqEtmn86OoERF8AW4G6tU
jbRIgAfWg03yxUbyedlKCXytzXaI8lr5tNlSpplBP7X61LMkL+hUXuwBRZXzmRyCu5tUe+bcrUq5
FlK6kIqikfP9cPPNWWHpARJ/sEVZ2viIL1OLXExQdaUkCZVGFw/bvL9Nvpky0EMvJ76FpovTT8VG
Qq62BuB/rNTJTpvmSY/VFXjLd8lDnq/Qk6VgJnIAU+oowQ074IopFJuhEnYz+3RTiF+YA45G61d7
nIjIujutR9hxArsFVIJ29tIuP/i6dZNvlekHU9Y9IVPFffBx7oxVEPIdgabmXssd6UMrYbOKxlB0
evPNofHzo+GTg8hCNCLO0eP5kQVR5t0B9n8SJdQ1mSDd5mtrN1ePSTi78lC3iZ3WAbTq82ViaATQ
GH8FlXqih1ksiRbe4dUEgCV7Om/7miGbXuCX1tINVI0uuqV9Z6yydXsIOh1Hf+KQcVK8MpSaL7Tf
CNm/ynsVki4AEDD7/5E0ug39XhWiXQFXNmqf4qnQe7QzXUFQxD5D4AUmREL6ZhJEzJ2M5kh+eLmu
l0mGtTuLvUZUHOCecp5N7KRBytoY0au94sqbCZbQMe97oFXclwTFzgrtN4Y2s+l+ts+9AKbMb6bu
Kvpzk54E9frrU/Ns59/y/T6omBnv9Ph6X4JmKBuPNNQd5tNk5z3RvJqmqRkSaQj7QpDAbT5hp/1u
ZDmKOfTkpCelYBNhlibUDmkx6iBD4LRF15cHYtCfpjP8edMClMvFiBPobsZCGAO6y/MulmbhWxgk
ASk8hYXS/yAarJSsUC80NXzjSJjMFwrtTblIICtjnG0qkXhjy1X1nSzBAlJUAMbOA+/pxKB2uBKY
decNpiUwPBHFklgBZuunMbajjoYB1NgO5QWI7jso0LO8nnQmmdo5dJ79dinzSx3ljdB8Tz9Vxxdp
3q6oAPovtdU1kt5Z3XMl8A7remMXOztzRpImn+RYwaHjPUZbROCb1ao+3c7XtfLWURvWdBPD2P7O
EFanEWIEbFM1C2WjUwcayBbHpI9wWnJKdhczR5oaUaNxn3z+NWKFpao1H1KJq+ITvcexnUxBE/Xo
yl7KlJjDmZREB/81bo8th6PwQcQBqPbtl/Om8Ur0Z9X/YL6JtPF9AC4/3HRi9Nosx4AFhYxwsfXW
qSrI5tJTXxfbej5KJ5LouI7irxinAh1bkxadeRNS6IAlogRGixThR+9ww46CRelwic0AyNLvrQ9M
dYpjTL/8BTQSEfiwjX118ruSx9vnedQUaFIGf1fOBxtjYeDKr9SZCv1qTWnRSieouA41WRkRWYWv
kDmFmTMb5AJNzagfWtlK1xQNbeYqcsWQMTrnckb6KSjjvsb3ZZ55lUcaOkKGojhOrMmG2dNzTqQa
kgSZhRM8ji1qIa+aZnp6gSoLVbhF64YVTbH2cx0Og6bOgMvTmd8tl7QatBkD6Bl4ADtcw5ZUmtwc
7VV+vVElwJFSIbm0sxeR6fc9fA4xxSjD78p+ru5vBPYsO+4tA3KBGvwmiz1Bg1jhPbHqJGoQi78T
2arEpBRz/5Yf2/BK+cWr5G1nGuNuBrV6zWrcfaBhiIcKZIXdyZGEtJOM0UFsaUFP+uxZ1Aenehp3
VwKvHjdfRpjdzK14D9Rxfhi3AtR35kMqNsIpGy5KwjXDwZqZJpfTpnRD+fb2cPqd+hrPpi42lsRR
Bwzymo8OO+7NJ2lu4VvFVohMDhO8m/LnC6MNlQ4gwOc3XWT4z01EW2/v1o7K3IKVqB6QAza7OzeR
Qe7HDXpm1fpf8b/VFAKSbLaN72GNZftqJm3AecDQEfEOg4cgFNQOPavtOnjIpik1Ko+orw7Dqwqo
Oj5PFzr2UEP+j5aj2nbFhvltYIcTcakDBi9eARtYX4+cV1HTDL6bVyxiANu6xiTwQYaN0N/SzpYp
/XkR6zay3fIrAstvAaXh7ITULJopIWyc4Vg6Q/RuDrqb1fogVrAaGld9yudIUkyt9irF9zMH5Fez
t2kOG+kwoUMjNMTv53LyHMhj2T+rYTBD2sBC6NWsFhknwd9uGKZsv/9RidoY8bf/NKFbPXMZ4z+Z
A33/h0PnQP6rNkRay6q8S/HtIUxkXs3uBqwClPilr8os0Be32AWyr4ajHF5FwJ7FXKXOdeiQlaTE
asafNHMzYBWRTKfwV5LaYvLMFMpZmKTi5cpV58ceolPV9Y9gduhbYq0kmX/oZ4d9UApXguLY0PjR
T9NcruHdCmbFBHDF29jow2lkK/7iI79hUex1Pg+HhYwP915Qkzpk4TBW+KkgBqO4cMXv86KjZZUo
gRqEkwUbxDeU4GJ2CK/VSVziSThcRwsalrf44SGfrQLF7Bc2hKlNp0EcjOOPreI7VcFnxQvpqZzV
c5fSfLpxOa0hKzyzeSq+NECjXgsyNK3SWK/u2969RaA9rqRrvrxSbnmkr3MZGVZyaoQFGgXdd6Hz
du7DYffwHs6KTiHdUrAjHy06jVM0ITaU2604aKqtlbHFGk+KVoicoHzANQZVDxwMPErFXXpmE0Vj
s71b1x0Zp0RCb4ak35DibuH/l85rPNBt/Xxwmj6cpW2voGimRmgq+RmrYbeB6VFb21+AldQu1aDV
rxpujEV3BCjZRqijXKRjJvMR8dbV4EscTaOxxb2FjG1aPuXkanTjl25EXJ6z5FWyJYmzNgYgkKDb
K5tn8GLm4eScGtwYw9xc4M14FnWsH6SffOcTqlnlvjwiV3sXiFdZZMH40vxn9LvmVMy2mYNUpHnk
GKQTA8qpGJ7ApJmBTx/iMf0+CM68EfRhzJeJNEVqaRLMwWnlE8Ril1/uzVF+oRsV6jgfjAlpB4GS
bOoPV9Mp2a23nPjmm4gXd6uM++e29vD2FNYlRAyAFMnqSEsySSJm5FId8GOuQt2Cb+sR/MdAL27x
xh9RYIJkrExI+qvTLE1EsvJn5wIqUk+WwijowTOs4XpGDrHY8Gxdu+RbGQ0ve8FhbTO7ZK2jyI7F
qWdtZe1/13M73XnyNBgJygfHIV5WXU8WGY35DmGs5tH6OYlBtVNkCwIexOEj2/Z7CG7VaiaAkWjl
JQNMHPsCwUHwPoX0CAB7zmSBsKo91puv8UA09PejkmSiU8pPHKTa5t2xUBVCSzcmnjdwDGljI5QX
bT33BV8Kv7/HWIoePphCEKUxMJc3xg/KxSw/r2cZ61HsdkkiuMcIenPj18g2bBYVYpm/NhoHe8Cj
QYS6Ghq8zHAPbhmvQusyVGFSgIigxoJrtGhTaOFAlSFE1iBKFP/Jtgw2flJcQwJpCfAdmNp0Vyf0
/nmVWSNI+cUnZkn083URSu9rgFbmAcqQqRO5ACgNdUpiEeJIhScIrlP3EblExsEl2ZPM3sUxcXO6
x1Wbe2AgQTe1af5zrE4sniZzeWC4MURsiH2hF4J5TSqOMoZKUzNCSOcrw26v5K4+g6qOX5mMQyRA
jDA+08KkjebS7AgTk/is+30wK17YN543J5E8ZItulWtekFRKkOcs1V/8b5csJhEkgogYBi1Z03Fe
/yNHqAca9rrF3VMF1Tf+97RL64qgwmfz19bq8LDq/iEUIommUvJro5gcdNybhGGE9geKmZjNBBz4
4Rhuj8tcX4TeaD0ejiQ62YZrZeTRx3hLLicL4FCIACZqudwqvlTqe7UgBVy3m4GLyTuWYdbzdFAt
qHFVEBeSul1UbD9Wg0x7QGVCBZ9rEjF3OIyl4fJ9NvR7iYwbr9+rZM90x0qxnK9nHwvaLE2B9pCd
Usvk24Wdy+1CFridQa4CYMYLqssfBqb5bLv7bBny8w+YnOeFn1H0RNKyZbU1H50jKfk3bAoz0QEZ
SO8NYnw1P5fWlOAtIC0f/r8xAWQt5glum8p6/a76Cjs0i+9dhV4HE298ipJNwJxhfttyjhYNWDlw
cX1zUmsUL4byvAAhYzojk6LgzRLnG5XgODuVxmI/xh99l5iE0/oUjEZTroMAZxp2uEqhRKdSAs0B
CZkVVYuSxlv7zKHHkE4AqE94fKddKSjHoXXLPjELFWQguBO7wZtx7J/24AhucGYHIfecv/cdASUV
FNsXgDsZxZtcTfgR0ihOWNe6eJAlWZlxB7iVcxl2kqdTTHO9oKnlrJ3gWlTv6WGYy5uYRwxulxiC
YIgxj6SyIIpHzV743H3ZaZCGqgFOndanznmwvAIggodVMfHe6dKM7VxjXu5KQzOOTP1nf6QMx6wU
k+RM3zxxszMCdSqi+a0h9zHLK7kGPxqOEI/4iIcxHzxVj5yX2faPFqDt75fIKDgNnVgi1mk2Wcxj
ftsk40SBUYupfGhn63dZP0EhN3i3J93SSRaHyl0dOar/S9Em4bhle1Kwf+QRgYvrHh53ADoDFqsk
aaqbgDQLpIeaRMYMWGXsAEw+6URHymakXajGIefcyDxu2apkHV+R608FMcqKChuu0fEBRQPdtDVH
TKnYWSHgeJqOEzAGBlZ31EUjT8VVQIlUaQavISa5xYHbHUdbPeuzLWgtn9uJKwXt1jq8wLCYKOeW
LjkC5kJUNChlHuoAoX8m9NzsqUIDbUWMOpohN/p6/5hDHP/zX6cFRcBTPlq5lS18D9cDEbAxrHW1
o9p7HnMvunLjT6eGjDKrM0U4v/RXl3mNvyaqyRiTZjAu5dyS2EGvyNJoXKVjxDJRKNIJcBEihRGq
BFHiu8poUgOLvLY1/jbT0miaLmTRJinX93ml7QY5S778aSrv8LdIpt8tgzgl+o1geyoihs9hVUNC
Trxwe/S0hBJUCA0v5JeA/kACW0qrKPfFhVYceuuZY+9Y4sg572mQs3uGRnI3Ht/ODwved18VNcDp
u+N9YDkvfl9lNilLc5GOUWQLX3MEWMtKKcwgdkqJ1e3RlgV05ahqPzzaA37WK1Kd9vOjB3fLNyM0
VSn1oV3SGTzV+83b9I47ElAac9V5WIO41bs3hvX0klMJqFSPJI3x89AoE9wTW94+qJ6rEuMjEWDL
Mwe46vfcZYTZ3lI7EZZQ/nFz5W2BUPa69jsWg1mgqhCcZGJ5/bIIuue2cyrEE50LFRkF/HqTjLTA
qVkzozES4mBAPz5d8Ag+lsxDT0oHFJLRykNEUsBMwh8QcTU9vZO07oflGl+ktioqSvnAszqgtOX6
EPrQnzmg9XT0YJ9WMrvB0Vt8EZhLKDd+2OZ8P6agQ9ckrAyP4N9tCgkF40qtgq8eXqkV7gotAn7p
xX8LYHq9KP9xFVnwpf4kPiK+QYM6Y0z7VUR3yZME6oaoaPn4yEMe8YMDUEIQZcmytYHte7hEMLDw
VTPIsmNulxksUXDHyCMVYBwcZuaEJHAZcFebr3YXAlKOkumN44272bZYUEGBGa+LduRjB6m6I2KJ
RADMkYU4wmCMes8jHbXNj9S9OCBAH2ZH0p3HB67iG5PB6SrZwgF47cLPW/cgnjDl0Cg7RW+rRp27
7mM9Ka79CiByPQjRCSs+kR+2BWvtgdYrT/vfHJcj+fLoIaUr99RJRgTUdpHRneL/a2H5WVD5GRBl
RMrV9w2xXU9a1E72IO3wTIQX/v9BWxE1RuGpNFDF2NlNI06N6DZ8CzLT4BoRbby65wvg7wuWCzS5
vb620X7puD5b5BqQxxaFERFF1Gs6ieBfMnvFAj5t0PJsiJVI3Zu/NQCUAewSLUaJi8Ej26uJ/QBh
aYzaAZlwsU+F0iKiPDTtjkVv9Bm8n60NY4jW4cVzKTK9J7ZwV9wIbxBFtz44yIK2aqdOe3GglH4r
4BQT0315/OzCHBfYpeeqkF4exE4vKgFg0lALhlVI6WS8nRNG57oYQYI4osuzwb42X1jT2zB2nEG5
Cx0VLpu7lIMU1GNtwBOj1IEMstP0Awp1hFjv9sLaCY4XcR8J8JefCJ2hEna2XPvbyOByqkel1Ys4
eiIW9wvIxThckhCn+taiLzkW1DhuDNY+YbQJjSLgxVkaAVqEcoeV98niotAYB3sDEb7zaWYLULtj
rtZTrnd6tEPTmjmk3Tsh9E5Uceq6n7NyuQu2h5p3bGQOkqKZvPI4TJ3ibiRUEOjlZXYVf2Pjkk/2
2vtKXFLG7HS3dd2JZoDRkrAJShRaF2kx23rUIxxuTJ6M8R9U2E36elE3CABPhobYXx48wIIJ7ov/
uTzYRv/dnsVjnWX/7GWaE0Vba/1OtmMRBTG3P4gI8+H93gTUhFyOpYYaBZArXjXEzgu/qhZey5z8
/BspmWmGBXBC/xZRbBUmvvLVnxh+MsuBiucRjr8lSHewjw0MMk3ws7bGmduP0Ykj2tAwPug0r/eW
AG6prJP8tIhGln+xM+Shg+d9JSSly08xfd64pmwFZ4g/CkOlstekR1l4FwILFYTLWp/ZCtxU5CPg
29CUztYbqee798jgrjk9/Btf62SuBwuRyJnJAOKglucwMtEG4SDl01AD2f87X4l/oDdSIlFxvBL4
d7MsRllfNFMei2nhrMxliElclLhUVD2Qc1kb8Hp2OuCIYopWc51HgviXtFSeY8fXUFZYO+loa3dt
EV9BriRwIrZhqOEM5SQPq1SEm9h+Cltiq+LitdWzBBuHQOoRc4A1p0ijMNRqDqghVz6R7oCax4o7
bgKcKNBbwBNhPtahMC6Lj1B5ingaBQHX7ClqCaVG4nKd7rQMvJ1nJ1jr7GCmSKXweBBYrYawXGI7
vltemFNQwur/AgKNdqGSQ1M8VvR0gaf+obdEUR+q14UkXkaZmuPgfx9mHivvAnDlx5SDcdWFF2Jw
luzFfJyw7qlJq0nSyAPOhgeK7giRG3KIr9qj3zUPDQNQUos9f+ngaqHGXXs7t6O2XojSw3WRkTFE
r8ZfUh7Hx69DgNjyua6OZpPh/2hV2yTjzf8SxjTO9O3oUM8HmIc17lOZr1ruPRpnZpjvyD2O+qiX
LkaF3TewlvUSE7vJLCv9QZWhnZUmJWN6AiN8V5K2w0m2JWFLE1W4cqU+e3NEX+njcjUQnqnhrkpO
K21oKAMAhhOEN3ZKi/Y5sS3IOz7F+Hk5FgcOpeBrfCaAToje2or0GGMq7nVCrgpNQXcsXcwHKWNh
X1VYqXzx9inPQ5d/RAlINVVkiFrZQwb0v02f7nWGa6s+1Y7pteMZ7V+jdj+n3AtVYWn8sVbcwFts
bNKgSgdMW9NMRlwktm8HtFUmPYi54aP2JZwVaVSY+RtPABmjPOEPhhFjKzvBXEAHDiQKxu0l937I
u/b/i/tbjHcw8UTBAooradmimvjCj6j3flePrGurwqDnRFwTMh76Z40C/8JGk/dTu9N5yn5pHwSt
d6nlDRfDisBbRfHWRtYpHNe36aWahCOL9yguYCNU8QZuZNnDcoNC17sLdw0u6zJR92hvRYrpUlDl
JX2LM3eUgBMqvUJTCu0qNSeeHbUBG4132UH8GCFChmgFMUskRDw2Poaqo1CdpS9onwqrpFnpslH9
xIXeuNUp5Ye7Hvhl7plx/zsD+pCAXYyiL2eGWmuM0+tQ+ulb5ei6kg9QkIpP9NfyptT7iG7Lm9PE
tLzJtmp3lD43HjPJce5qv0aShAzdR1ofhDEwaNssUWW2a96rIxElPKJnm+RtWIrnq0DOCtnnpvfS
TRy9pyPIOzqqSMsAbyfnIbJKnDznJ59RqOZQcGd9KLg/izu+66RmqIpvHwdJOV/5Y3pjxrXvxQL4
ePYQoyFPMeTDQ8TeYGnxVr3hGQ3JoyubhO/uycbQoWKYtUOzkhTR7CjVS0UHuhqNzmYN6XquhLcS
+4S6hF3cT9CQceeabTeWk76xSYU/Q89Hgu4Hn55nvgzc4ZU2LvqKS8OKTQNcmJlJbuWHAucNFHEV
/lgVM2A/WhXYwLACbOIIs2CZ1hb5PO0tNl5lZOO1ubrmF1FzXD0p1jmAoy47UbIlpzPI/1voQezl
no23wltSit7DkiBOqrR9m1K9nkUXs6qNiGJYdzWLA/iLKMM/hGjOkl592RXpNosVjZeBU5xfUKyK
Hw50/beL0VtsjQmX8uUEYYa2l9WT0nYt5q3vgmJn1SAlsrNghTlgQIO1NEwfiuVSA3Qe5lIGTMS8
JkD8YLTbl3LlvBCzCIf+H5oIMOfkRGrhJUDiQtAZZuw9tME+bGGufU8v6+HmKcKQ+uaTqX7vlL0y
xjDA/12X2yE6dqoqfRyBsG66Xjh/92fF1DoKUbqv3z3RsT34uzQ8aLBIyKuL6OigTIUmlPrgOTFD
FUFJ10v4RMg+wyzUH57HSAcNnM7YfypufhIFlz8AnNzLxiQ674ZcTwprGxI9dg7knR9/Mz+paTWv
hdZ0sYf4AbBTYWFFweAXzG8JCAFHqrt878qt+oC7vogiOlO1GRA9EfgAOWZz83Q5GdEvAwL+6Sh3
IrinfUqMYosJWt9V/4pBkKmuM9bhebYqRoAqkKtXbT9ey6yRuJiCfeYnigIROlmMN8EblY08RLsN
0E48TZKLu9v1q6rKmb8yypHFR9IDx6d6LycP8yN0/Tj5N97hMx1O1R3BbFuZR+N0fXBobQGYEqxd
59j8iMf9E71xMSxpuIu3xcdZb2cSZnMTHh4pszX5Ve3k+DpXM6VuOJmiHC7WHwVsbQ5lWPYWraM7
4Zc4CshIXu5EHiwuaoawjir9a9crLNJGA0FiKBCOsZmTKa969LYEgdwdQJEJ5B1M5wCnZZwq1FR9
ssQKJ2Ntu5lBopVebtSxqQY7agVthPbZNZxsGcSgrMQUSldalzHojV92CkU+umxeW6B9zp3s50kO
dPwWtzsIt+aFmmwnzh3GzPUzZf9tbNLPn66Gg7bOUtEyn8AHUQx2ny+zQTeYHmkrav/zotx3uzp4
ieb6tEa6oaGRbpmIF6NS7Il6V2GiVQAc3wiJmRJUsbJFjzHesnNHHpHeVXGcK8LBzrp7eG83CFK1
nd02urDPY1YCPl6GWiL9DMkEpnoq0aoHty65zl1vWK2/pb5JEfRK6UDJLTjN9FPoTnkI2sqgnEmW
bJpkFcCmCOcT/U6mdmB14OAgvnJawV+2HGdMENfuu8g76q7TiHXTNbnxA680yIssSFX7+rgXWC2Y
0GJcTSYEOPDvT3qNFYsUxnSwdNZZOKraMWWnruA4RtAzYcGMe0MAkxfqf/u423iQRVhPlriaD32f
EeUhcnSUBaGn0xwOtZOGNbJPgdaiRK+UghZAgVJ/NMwILXRLw/wSyAIYMzS+cKQzySFSWFWygyiq
yFgMFhbEGJMGyg35IUfA8SdL9K2P4UQm1LB7Mk0akaF4tBFvTtCtstvPK1ujP+eCkJJy9gYZjuhT
j7YjdYTU0doUgcxdw6oc0Bqueoiqb3xUQbQNW3hjHFLbWkGhyM/FxIo3P3A9j1B2CnPSa+Of9BU2
B/BZgwcmFNv5xyIniaYEo7QEiTjy/tTF3rzSBh42dsWUo+S4eHtVrg//imSBYG9TlqMTUfxW2PKB
ti+PlEG8zr0a55WSkVUz4L8kgmR96Z6LA3fbgTuRwHSK5DqMEoLKjXpXmQGfuZouBASNUgSayOXx
R7Xb9FlT7wu3KB2ZK5q6B5mdclf0mfHCTRWDseWdlsJagojEleujT67EJGavyYyVmqNvtMyIlebX
I+QN5lYtetMVTQw/yL/h43ybUgCaq4H82Up4qW3CcoRQWJ7AX0kr9J64qN0iU/Nyfo4AF5tqAzJh
269lMq+m7C2YJE1xYohfSNuY1lWMaQpKFcZIBhb6DQ/zSRPlBOnqv7ZZFDUSJ4Ic2GibPrL27Qko
nOCc08p/ywPyvnewQJ6o0MLuPWFkiNYEXydqcnhN4fNhQl5B/h+PUIrsM069Nkrqi2jbgSOCzjOZ
lF5fEPEGBuBWlQG0cZOMR35S2OvMLRDynixih+mpEz34KvM9mVMJ83qWNFFwpreu0z3pGWnxHhES
bsMWWa5pGkD5/+GWcC63S++Ih3chHig/Y8ogtNiEkwJGaPre0XcJSriVHnDohJHTlmWWVjTJ+DDy
Mj+62GlHY5QFYVtkrTJDv3wj8AvSOaCXqku818azZ6m9ZRatoKBkJomEPznoT3FzezblFKG0L/s8
hroYRKrwk8s4rC3TZZg3C+cvguXwa55kzZ6/3yfXDjMpPEiwBAL6TCRQ5Z60xxXELhTMv8f6QuCA
cZPOTTnzgmqk2V3ngyLlkFyFjMvQeQGcmZE9G2Pz6vZAESiKPQLBKcH4gUCWoYSp1WaFhqJVn06Q
cgoBVeKT/yEToEvovZtugZtcOEIJr86ctyjBgbajEUXI6hvUcLQXwf76mZ45a//HKCuZ4L9JANtD
pHspekC3WwUwCgaUfNDI04ZBxLjlvwl6tZMkes4gEIJ3glWIFeyptaw+JiWKfM78jMeKGZijiz8k
XdcawjpFnRRN6TT+8h61qHIveQ75dGjZCVmt4r9x7/JhmQ4ZfyyW07oXEdhzekCUd+2bxhDUHgV3
5/kvc2h+ohfnP2FdX1USQTEXpZ7Yyr2fKoRKlJt0vfmaAyNBmTSJN+ZlF2zdvib7cCII7C3/Xa7A
MYBg22T8c11BU+Da9xIrTfBqX2TqNI1lmctoRJ8lpND+PJ6q6J17mvad1eVzSoy2LzBfxCFKBuii
07PK1TiyRD+EIg50AywedaJMIlW08tne00rlTkthpiK9QzYDmz1nu7PolSA8xOnhKFz0cWDOybTm
QhipLTLAD14FVovdT5nhazSL3M6/d2xKRZUk5uFf19OdCZv4w3KLkCpXFELIlN8L+yutylIsVquY
RwZgA3puXX40DJxZW23SuIWrvdPutay7jE+GUyqexHSW8UICJBT10oU2CJlkNALaYA/CfhaaEYDf
5ZS1dQw4WhCXgjFGJDcfbqtjZAtY+j+1ZIbOLoHEkux7QdDgPSnHbBC2XAPgHOzliQm3reUNeKR4
Y2xNIokyTa1N56f35U0Pd7XUcvYtZ8KjAz9QeNqAZpP3KWGb0Xs1MwMFRGWH0S55yNOs5m7Cn7DX
SniLfIZDZV2YXmiIj+rFRbeksJmttLjCDGWObMYmz49A71nFxzhfNroAFnWgyokIGGUX6ubdDS3E
uVpTo5xhuMLsuGvWuFprPHiyywHDVMi1o/hqw4W04eAfkGKOHoy29eG8FCtUxwZb64SjDkGpYar4
5+x2CmpNDs+7IRYEh+UJw+3Oo9U7i/6v68l/jJ+i2RTFwINAM2LQYv0mM7pQoooT1DkBSA646Bpk
mAaIumjlaxlJy5V/Kdcvow/Nbu3PhUxJuvs+Qgu3qBdAgnTqg47G/5QguzD9aaJNmF/Fv1nG5e3H
E4mk2LvBk5eA/D/dHtinovRN9IlM/P/lLNA/+vuzONmGR/10UE1zUBWruMdTbdFC4WMJwUqT5xwj
SLgfNYIlbnIsEBj1eOz8djB3N7SOeucWKUULLBBB52C5OSaNzff0wEgBx2pTWL+RjGh+gep0D3sh
rmjQRCDOxzK6uMVz/1/iKwYPfvI/BTdTelVTZhXows60brDvBK4l2oK4KXfx3Lw/nNV7jtOZ7no1
wSqUs2sZpiRk/iUuhoeHI/bsFNMV+dmpzeyXWfRSgxzCq33IQ70Y+SddFsTNASVPzW3/R7boyAWt
RwN2Tob73NeR4Dl4NQ+wVU3K/7Lw37cSwVEAZpRn9RPzVD+nFKoQVE9V/TfOE6znPnDxWLKUA2p5
qJ6Wx/0A0t1STnWpb1noKUIhheBZez1laEpGdtnLXUvPgGMvU/qKmMyISotIjGtNg1mcWmqsUeU1
WMfTPXV1Q3PjVcjXKCJ7anMpPBZpQki/cuhpQOPZ5LYwxKsVTWoEvbsw2sLGm4yk7nvyRC6YgPXa
/UJGyuJa7pFzOeVe3RqIT/AP0lwydYshRfuMYarOXAU+rQaMDq1iEQ5bEVaTxrkbkFFBodAxOP6Y
jNtx8vQbnuy4SPV4d7bCk+88I5EM3jxkzcqOJJNTpLVF2px4StzdaRcSJuHZAoA9VEd2193pKHud
3gHPV0q+wvQdf9FVJZ3nIFliJ6o+8ZLJPqiutTZuy6F5EKCfPG4TCQJwJA20uK/MmReBX2Agi2OZ
jgnLD5PodoCdujlre5TIJsSYaMIRMOcBcF7LeX3Y6gHGEr23KbvUZ+pFnXS0rMtakMu2dyAjDSpc
vErUU0LjAV7HIXo8Z5fNdl25n68eSs1gnnE/VrkKuRgAGywn1TbTZpKU9w3cp4OJN1caspnh0NfF
z3f2WHLhCos2+q0bR2Wk6oTx4lm6c1inhCYdwsdiQQSHu/BQlqqIGRKE7J8ad2YqfEcXCEyGjNON
l1eF2r+5g5cmCQkR8QzICeUqBV6u0YyAhZ5n4FwJlQcexH+Ayts8UhwkHD71Qp7GsaJcxy7y/VFp
Ip5WCKjcFcNaGPqRJj8m8r0YyxOh+t6FLS+e3NJCRWYnjnDVWB6o1HB7x8nwzHRByBMWH/Cd8oyq
CRcaZ201ivh0MJX3mDAnkRTD9wTYaqn4ybkmds/Z8jFkjmhr1WN85S5BRFRkwHlfUimHwmU99sDc
+FX/TdfEEmhMHcLqDeXzEvAA5COMmAoIJb2NSDCBB3S2je6ZStRTTCnUbMWLjF77JKDJqWDHA7cM
80NyBvBtm+Y6pEBRtKNfy85dhesqh0F64YnTvTWphTdUIcA7KJsR7WoJFywZf7DJCcBQ+13PJBe9
ZS1sux9LUh+eJXwFsfadoLsYaclQKZ8MImLznO+tWvDo1XwUDLHVZlw8UmykHIc4eitErtopmylY
8Y+Q8bPCjWui+q1BaTcLz/pKD7yJa5Bq8eMenMXc50UKj0/OPeFryNwt4tnC+Sye8dd1owPmhYQ+
YH2P86BModtnaP+ge9K2zub1TSaPOx4TNED6g5rupfkE01YFIDcmif4yAgSp8kMtMST5pBVlJ1ez
R8MGEDh4jWhHoWFEONHxBhJ1XtFaCgzXZ5wJx8/993QgeU8g/3yQ+On8Eby7XdBBmT0aqZQ/dArA
jAUvghWRHuVLi1iKXshHrZKOv7EISOGqctk9uerozpbe/UyFqzk3M7CaJIup2HEJJSfjCVba9IOF
LG0cs4xttFAtjAtjXyERW5rI7iAyKivi+jmObjRZLx7RUxXwKYPJg9unBcArp7HcDKX38z4mbYSb
ErWie6WV8OK4+kBL9xoCE6pMKMWgv4s94gZ7XQMN2xS7aY03BPkkhQ210sy0GEcAnvkiapuFcOE5
uhJzR5mIptq2I19jULpRumWwvIFKLIhTI1XcEV5JDaH1bNJx3vzThg2wKebKMH3sI1jUzNBZAJev
izlviL0H/akF8ZTuh0itgXMf0BXWJviv2Lsze5bKkvwJV3oCZ5+dtF1UJXkbFb5X827d5nmoGyd7
JQ9cSz1KUAHc5IDoRuZ0o+2GnH96oT/LgRlQjs3SUyiY+D1zQ4CqLEkve5+TKT4SbHrWVqgCkRDC
Y6gW01aloC8K78CTke5QsKqoMlZcQvluYUQ2OMnM9OOo0CWg/pe2Njsda4osqJroL512DIdmuGYi
yMw6/7hSmFNl6GAWxhyBHkTCM5IaNLwhLJE30Jz7qB2gzeZraoDzWLTsNmFjfd2uKRIob6Id2rsP
xzOCyziyQTgOD2rZTitY1gk/Ors80s3bl99Qgh4IkOE2VnoD08dSEJdgOGQEmdZxjTrGj96ngfnc
w1hGoWfguA9K/BvIuXGEkNKh84eSEN02xbpJfJNCC2DF2xzPoZ1YpqrZNLAt7mE1NLi8VSiEY53l
734xQqM+8hneUOB+33d12r9Jty5HiNmCL8B4quNU/cJ16GR62QoY3D4Ky388dlsb4cZFNQEaJgM0
R4+qZKlMip76kMk9vAJD3/EOCZh0XfMTR6WgZwgStoKcESVaI5QjeLM9MsZ/Fno4dHx/ULNIy4o5
wg01tdTE2EOIKhdw1C4TIAnGM1TPNCosdvYSdDUeX+pSspkmURfTBgAT8+orWO6LcgA0SflF9ntg
f1JyAYdvHasBC4p8SYTmvgJCvO4ANOxqdHIVVgXfnc8hlEselOYoAzrNnNSNATogb7+exbyVWnE1
htagKPazaVgBaQHhiEitvB3ZqgUMXgXyAgc06vP/BW+Sl1usoaccS897wAFeK2wzE6+5GdLNpFV1
gDfRav+ndjBwaB4znhSJAI0hlw4Tg5V6jxWT4HYAGJNe6JqHRt6KVPTblpTSRAPcjzWke8zzhx14
1F2mpXAwY8RJBUR0Fsn6iHnWng3AZXIiGlkg6jXaVsnvyeeieJnx6yAV+c+UI2t4OHGTFfTyg2Ox
j2FXNq+HyoWCOR5Ye1JGQy1wZwBcQIko7h4ZdZ8VJL+cEAXhh0kcqAJ1jrGzb10B2WQnwdxGCPEQ
yfCJB3gds0sXNO68Ufo1CqUHgE7qCM/k0iT/a7oKqbhjabXgWim+56p6Ax8ucJJoWZXrMsvG/jC2
Rf3Sl2QArcUJoEjY07TYffHnm9r96eM8DpqHK8l/xJuDG9L/bZX5efaDuXGfjKs/FJHpL5RVEDTi
vR69XRU/6pJeuWgc/MUc8NWvVMMAo7NN86huhpz3ldHiODX4P16o08y0AkpItlp0VM6u5xcgU/G4
RJVgY63t+w8ZiEWgSRntLScgL6cs9x6v2xZmOLPAvowmtJ4fqJeDb5gjkHzRQowzgUVY2w3R2Xew
Cq++DR5P9sIEXhbMZZQoCoxrHBv2+rK9yXdd26RFSQ6NFErvbXS9JwI65i+/+T0HIvIChHo8h86P
4H0JXFBkBlPKk/d7aigMM5vzpqpqG5Ert5upk40Qi+RU8iTNpwb3hVi0Ytbmb2a8mQm580k8qTM6
+R60yld5V59TZL+vZ16iFnoEEQGXjKLZretT6tDrHM54CZzAuE8WnqvHAJXf5DmDC/MLYPVfHazq
pd5eVlx2duVS+HClYfFHnt+HLFMRyfi9xX9BXEn3peTWxEtrlVTY6UUamkINQnyB6/Va0FDvnTTs
jLLXope40nAVwzx+qIAI8E4cRZU9giHdE+wSFv/fJg0lcrDzTgXVOfz559FefrF0yJps26xz3mz+
N1+vNoKrtoqXrU0naz5IhUzHjL8yNIcBF4+zbwrVGMiU+n6EW1ja6CI6QNrZMpqb9jtu4BWJ1X1f
CL/0VyjjYMT4t7Hez3tlEypgixWLvFyaNvnLLZVzuthfSC8b6hyax6ogiJ/E5HoYzojudGBA4TlS
SKwqA+nNFi8j0p6FUghwOMlWt+/Yx6yq882Lub0guVMntNhUNJ2N3NdgxokkNQM3+z2W51zvIh5H
3J/afrVKlXrWRcxTt+nHErPCPpBvzjal2TE6fK3469awDKP0mebDYzNSDqJYhDnNKDCCHzhvLB5F
Dga1C4HaZq3ezMw+HYnhfzzVC6JSfHtTniO/q7n5wIyXe6bzXANU0b2LbgAAz2IFqonUa/zElkKH
GLcizO8BK86JKCjjDmd9J4Zq3RKgR1ZS/sR2ZP4yRRQZpETC0z/xsyFps7amiSSB0c2WUPjdxC5p
DvEQ6ZlCEosJBrssxk+/hQrq/75MQSjtNCmrp7gKsZx5GXPfnIwTeAr6xhqnL99cejBelmQJIS3Z
h0PfMWm1pAGuWtfHbxJzVCrcS07J73ThhUs/XCUKl/z7w0rwX4kwbYWrDwTyqiFsLu4fpqa0kd76
qxgL9LlzKjKXtR2tGGnXWoT4yDN5V7wQTGRatwW/PFm9eenE+lETmBoGuI2BRwOmUyguWHc9GsGD
TeGOh59cv13dWNQhfeTzYbByi/7FfF4jNVnXTe0Sf3zDeE10Gl3P1hEe2m4LZhaMdhK+o/ESgtyx
hVlK6SmqGKxT3ZZOYEsdJnyvFCuBihuqqeRFGxKdS4tF7r2/3zBCr+tTgTmUTD+gYEV07hLKK/wL
8RYR85feuH2e7dBOLKFYBx/wIE45p8cZCkyw2j7+N+jRXdAkFwHN1mgp78WYYsTBSOayxc19IRaV
GM7PKgzirWt1m+XVrTHRtRDViI5E6gnaPZacnCLKs+CMDXAVuz1V9zoFIYyOg2ENPRevUTk3zh28
+/YCv9H1zpA5akjvyFLdgyavM0n0jLXP3dUFFTSYLobsYECP2vqsjy7YpcvgSt7DbSB9M/mWqLuX
qdo1jdVzLGLS/UACjbCt3+yGdsk1Z9Pk+iQuZ84D4Jm74ZMGjiCQisA9MpkCqNC2OPeaqa3GmEyn
G/1zZNV/4197tIFbIeCMn2Tpbj9iHCiAPrdeybcSt64DHBgBQO9Uow/Jc6hFCE3hOmoIWGaPnaHt
UVbfaRATkEq8zjcVnKbQYI4g/ACbW0Bdu5hpY02V21dtFUabvw3NpwBEppmCAuve271692EMhJIM
xKuTcQ3bI4GirwIq0vK5goGjrdojLvX63BVUpKgeCVinEZ7p+4epkeWUWdudDhEAdEgnwxLxLSai
f6r2IIX+RwWi/SuTt/LOOiFVyN+rYc8XoPOfRoFrAmm58zcCNyFTghAjBHxc1JitTVomUho6kG3S
YP4ARJ/DYNesHXgvAUTuMIxfdyV/ydpQBFCM2ztekCLTS9Wf5KCfUM3wDjZNuohHnl04EqZ6ceXH
vPyPRCjVy4BSEt3vYeV+/txxxuah/gReK1kB0a2TVrRadX/cHkCKAJV0FlQ+g8fdNDLggDpJLle5
bBxwK/TCqH7l4JH2bszvc5grO+SbxB9Ru/pqFqgFJpxG3dj4qbi+TN+2K4DLq4APSFIw1mMtk/nt
lxXPJR4VEmySZExGZ/oCtzdt3RrEpEgnn45ILKjSqiubBdLFwEFGp/H+R/0zjxYPZc9eo64lph3b
oyLBB1T7GE/FtNSDBtai7oFjrA2F0whmK968yvpu0L2Y0m5yzcyoRgf3tBFIkZpqdIW2bV1THx7s
QB10JpjuDUcvJcNTT/sMp9JvPClfuamuVu54jbp7+KF2tUID1N8lGneCcMSIgN3gEfXl4P0IeLed
XKqc8S0HafzfSaTtDpPx0Io+NtDvKa7dCYUWNPfrUdasiq0Zz5xYIHW+GmUZvFIz0M5l7v9HAN4M
d/YovNm1ZhX2Iaya3VyMwEWTB0QMfVkkofV5wscZrOPvfL6HdUNhahmfmuCiNvtCq4KiUOzu3DVQ
gmjyh+3aoIAZMknTMmHHqQ/5sK/JIp7cfb4exu2e4N6IZ/RYSHFQMn7+B93NOF3RfL9ZABzzAu9m
fV+Jvtjs/lPXkCAFS67mduv/pMPXqXtp5RsFsUDIcGAecKjwV41a5lMRkeo7N28jPWVZoG4bl6IX
3crkjfIZcAkAdR7zHm+esSTNxLLHbIi4H5jjVIrT1j5UmNTqD1xykkBf31n5vXyg40LGlttMmX8u
0uU00r2NQNpL65OkAl09vYu4pE/Jkhpb6ix503VE5oDNJSZQMF2wLkf4ls1BSewlyn1nScuM64vN
5LqBEeFdv/wkhq+gwvcxI8Ye7chTrtXhGWw+i0bpx7RxmUCcoPg157B27DUUtPyTiJJIt2pYjVvg
kod/zT+GfP/xoEbes/nV3WIvnbzpmfLQtIaC0eV+yIt64r4B2aLA5iensk6olD4yLxwL3PopoBhW
CExc3U3O1z3OKQ9qQV/nEDN+r+6RzhEfk0ySv9esyka/9KgxP9QvwlW4Uo8V445w1z96jbe8dJal
i+HAvfyZPsfNKqlrujIp2gklNstxZ9qYrT9ea2/2+3VRwgyrKozSo7sS8WHZxcoyqnFIz1bcYvx+
LOXyT9FH0ZvOCfRpfEhamzapO9P4+bhdPTIqanVD5fLMhFlahvGuDscnSGPyFqcWNVoAfmVyA7Nn
U6csT9fvenXuAupJfS0Ig5ja+rM7LuskV6RbZKZYqm7e/PKtxj30sd+oa/9kYqBZg/mpg5jJIR3I
HnuF+OnL2rBQC7eJ4pdXvdeK9ltMqt5565E2csX8ymWtUcK2iaj4vyNJvwwoxnYUu/qui5fMq+Gf
65YKBW+xId541NTSkNnXBMR5hsNvpSZCYLk4QRqLaZ5kpUT3RbWqk5a28fO2xsykL5esw5lmcIXP
ic6TPdKshVhCWPgp/Wm6fSk72r1IqKI1bfGU6StgnQdd/40L2o6vEsfc2VH3KNaH1HWWYOiOagpN
0z/oFHPi2pGF0kyXWIdLx2uAEc3ue8lrDJ0M5fnHhuxYXFz1OICyQBN69xa3XeTAFAEYf4RWfM7d
qw8EsF74D5JcwF3JXH04JkJW2EramS3EoRFmdVmZLRKdwu8TsMs5xNhRSh2fhuPARADY/U8jofOu
nvhOjSkzCnnlvze9ug2SVK1JkTosZ2N+X7ZiZkUdBAZAWNmPQnUy6JI/g9k72sJYpy1GzP6lMER3
Ez2Z3L20ZjNAfptmm0QsboKhIURejDt27e3l1nhL6JLbnQwF3juh1XpmWd4lRrecRXQIgrjtPcFb
aPWJTJE1N3McZLb6AJEqoKNWqqvBI6m+yxxoEv+DeBGvueaiTQ7EMykW848TsIi3fAFtWEgUWPlx
qmjIIgEjQXihMlhdeIdSMm6GnoKTl6gBJH0FcAjxcvpgy/q9u8RUWxvUpJd7gekZ70gBpXeEct2T
hlTKdWZ7bdgm9w/eI7HedQEqiqZ8/hRIVUrF09sg33UdpM/1Fe6/JUF5baPBH8kVoGwcPlVNIF1b
D6QFdiklXIQDt5QOAkaBhgufH+tcNItohn8997rbD4LYJ4+POaPZ4fn+zb8elRX39nQQdgHuljEt
mc4Ba5APc+AADaukS1QLb7yW+x6X1xW4fien4j0rnFreDYFsCJCW+8SWGZHfQPvfSeibsF3OXEDe
9YFQbXNaSRGNXd/upNUwRFn7Iprnisyyxvce5lhPJ+hg5EAG+y0x2zxgtbVwe/5iM1IwO21l6hTw
LtNQf/lD3QiDbJNXzDsRQhkMBtj9mzfYGJUImgdxFp5TYrrto24fY8PaA9JbSZ3qYne+w2DyMxEP
DslLPQZRo93lEd17JSt36h5Kbbsw4W4cY17NHGEUIVhwZxPbofLHDmiJO/yLHOsvIdIvOpaoR8Nr
R4MRWgGZM+Fur4tYez+N7C+oniusQjEi6I/ob/q1/akwsQzIpzySmpEIWoiKKLIoa7uwdAJ/sFaK
BaM1z0jbrYIJDCPEpC3363Dy2C5UCA6Jhj5go2l0YVcqjxPz5OAvCUsr3rNToOLJjb4D5pdkLNAJ
c4Eahh6pgKrcvratrO7oiPr6ptqeUGdW57Egl+G+MRd5lSpng8+Zn1CK6Qkxrc+SK198Cs6mKavh
vnyp+mRzQjDl5lREDyoQ+aPeXdWJKkOx1xnNLlkDzHdVr1bMnyvrQVvvWvDrySjFYzqMhNe384Ut
ZiKDoPQbH3wvIKtV7zoODUgRsZBAIwcnirwWH2FvIkbCZHFAooOUiWOt4yhkX4QQcIxUvwfXjnJf
s/LRSB5eHWhSsW9mTyOMk05tImZGMcGXgFpNaKfMZuXJ0H8HdTyFQFnvTY5LFagPk3b8Zzg/ht0i
uclU8BEcVjBLzzMMtv3F5D2zcbLifg1tNr2LdX4e+hs/k0nxq+7LlnDn4gJuwV0lMd4uLzNjiBJk
muTH+iZn8oSUEYmifJSPWJl9NcTTLQzSbD12RntzuMoH3V73d2phU/8lG6DJQDncg7nk+aVwOLJ5
DsEeL49kkTOtNVNMJ2NupO1gF/QY3JYkEz2Ha2Jg/p1dJw16TjIIiMxrQ1cqB7aWaaxXsmNprwla
d/I//xtcJ7MGAf62kAt50mo/DE33QcT+IbhplIUIs48jO/HQWP6UGPr59uBVfzFLM4bjAlnbbFzy
vaffEnVMQuM3BCyOe3paoyFZD//fBQUva8KVY5Oct/gHRj1k1QYw52S0QDvOST8aVq7qSPzje6a5
4iilGaJgcBqu9Cyr7JF9DwEWm3owpLcK1w3K/Om7aUc90xMVNeUKSKSRq8LglET86DktGA+lUrZ6
ZeONCJGyBRVExOyw2gFT/b//320sgU93ad3uKQfcyCFXj2szm3cSZuhg2c2zEuOpGEPQj/kyR1o3
3OAQ8qhFLGF+2HR1KM3F9yNwKY07sjNvucKeOKiZcBjUGHZ9dOYUiCFSuMNv26vuts3V+T5+qhLU
KBCzjoJ/u2Tq7A4Id8NLetbo9h1vDSqmFgabbIdUur1ILlp7IqOIA+gn1fG9stOAJPb+RDYdwq6Z
lLVUYcjRxWtkIi1JNbWidqzdppZR+Li2TPniJ9ZWcOvD6+5f2RXqzRC3p7xD6D743VacCsMQjrG4
HEkRpIuh6XxBGodkkbN5UzvjnruBg7d5J+8XD1Fpp0aWojV7O145YTXJNmrovzQLFGtneDbbt5ez
2U45zO1XDTtoaigmx55ysucS6rhoWaLfRrEU8f5/jgUVkxMTnwVDOgVf9OLWxqDyZbFnTq+iTadg
UqkdhF0PWzx42EbL5jS8PPbO0YvEu79ZY+KUAQAEo387OOCQ2/hEv2+BNkRDs8b9Okqx1SzH5Lcc
3AKNPmWZoUnUQ8Yz8H/HcXOz31+Xl4vNvwuX7a/sTDt9j33vNv8Xhd3+icI3QHqnLiC6XitRH8gM
6EHkHrDWNdS7PH0MoBAH9qCV+x6zC5DFdZYD4heBB7cnl8BnRm145sDEBJYchc9wza2WhQj4RVpN
OGWK43xlP2ziNRhvpfr+lKl5x8BkqhjC6N+WbZNqhFNdGMUIAmhIZPmwFDwmxrc/UEACbYjHmrRR
h5myf7Qyf/SpCWEI4MZ4NgUT5I984Knuff38e/odXmgPW/v5UBCdx0Npv59aOVgkPrLRXngMjbJ0
rR9VhJIOfrEGWLv/+vvt8hKCxdbWGecuXY1YBotl/RgjKdmCXbzzMYFw1aGxHFoxnlsH6aqBR8kN
VWcAocPYPySaoPMGSSpj83sfeMVwRkj61HJdepDR9tBMQWbHa0kmv3T+xX+sqtzUBbDt73H6I/Yf
Jz1vm0k5kZedO25eAX73NbOmHwKHcSNq9TyK95AIu/6sh9gwwePhhgJDulKZJsn91r46Q0N2RKOr
j/WWy6zVOcKKLn3azUoQw67NYXOfJhsmSKIKYCpBaBM8nmRM8JhtfWsz+GS/turHJOgdWm3YXioa
W1J10/PWeSGnZWs+J0jpfclnP9yP7DJGgwnaa0JoaDXFnsmJ3GIAVUhiQTuk+YOQ5ZyGYiav+qqN
IQhYy4K8FkynLJmtvQIVAZHSeB7+opPTQTfBNl33EHoe6tMkNenwtOh1/++eCytfpLuAReU9HgDf
gGmOsurmcatChTZng+24DVmQXhqcg581doQMHUgPZ9qy77i8ApKGF3HIpmbVgSw4nEYFCH103OVY
PL0xMLfgqdfL2UOjao9lYTucpxFTuNib48moKyiMtOR8RrqrABLlhFW4k/IVNwDRPaR0IfI6SFbK
J426NkSk4a1n/KkswHhf+QkMLE8415KUdWoTYylFkSk5Zb2GRFRhMvYLDc/bdWslHsZ0OTFNUWEY
Hsnd8KU8fha3h5R7JgxahB+QgLxEC9hrpJrAYcI/51OP30xhWwzrb0Ej1KTsfqxxXB0rQIO+ui5g
Jhx09K+LGT2jTaTMYBCgLeFw0+GAEqJx4CjDa01c+tSFSTfB551atNA+aeo3m/w7/hExOaWiPij4
D6I0lTu1D5px26ToJXXQes8wk7+rNkS6fuo+aIRYinAuTrSn1+MoRfxyWdyKAwZTHNh35vGa6b0/
eXqbMii/XwpN5hF7BuMQDXkZ0pbAtzbVnsbgCVWyAh6QsZQsdTuDRyJOCfl+Ebt07Itp2WVi9alB
u805t7FYts5tVPAOBvygT0J7Lc54a9r8D4roBxJouKLHa8TMOmYLKDp+p5dJVXBuJrLlNfrMVMq7
WKiqgC8hl6CiT0BXPf7fExtWgT5KlKrG9Xm2bJEDq5XVot/DVhBTex00I6bH3IbXjmKMdLBnO6eJ
ptbhxK8xboeIVuyDMn+jeVt0JMGd42ai+1GUu1zTRVI6GZyFPdKVUM//dBhQ7GX5WMsg7324b2IW
qejSW1M5N+IrAHL1jPGPRaS6tLZsCwYyTDY+m5M03NCTIke2tvQcpGhjyxtPwueKUAksBqCCQ08Z
kvy5wAZbidiFbUTD2IIcdoTlXP8AfyuawdPqkX87n0GZBO8W+R40oRNrjYTLeDktJnPG6itC3Rry
Z9voG4zC7BiuoJdoh9xMDPnbTn8mSgw4ElUK61kq1r9ZG5tTbG1+UXIJemvne2WK/qzi+zgKINVD
6vJoIHOInIRLXnSkC/gYkUgttbcrip8yr/DSB4LkgT9BXWCwGbIoppUMSZXJ/gxi2JGoRY/HNZp9
uU8i4BY6MpIbOskS3j2EzKjB5U/5Qi7MQsbu/mAxrDzNZQBwv3IQCOHWvZT6VeajfWFbC9tMIDjv
7aRiUsUj37bYp100CZSrfj+fAWdG8dnF7yWJb59f5b0Dy8KH6cqDwhYZoN93E8B+n79ofuXn5M75
P47IgsWxBf+4RL+Kin7D5yoMervM9raesn3aLwmtYP/y1/HDACqdeJnCM2zbOFmB2De0AQD2qY55
RPmujf6iHZkiCnDPQHJiIkldkz01cwYSNzfQKamMe1FEIh2C9FWNW/YCNvk1nddimdjn4i2dQhaA
/ET/0tN54s809r513oH515iG9LSC/SFm4DhWNi9NOJCtkoo5KITE5bEk2qOG6rJNL48LTW/uC3P+
L9dz3zquOrgYj0Byv+2T6I4S8cidppahHn3HcmGEIc8LQZhaKHN9fuMjzZXrEfNuyFPM08TiucYe
N7maGRlVeBW/fduZC2yiOmAheVlSbg8Ltq4hIPc4mgqPd47OFxShK7JYmTUqLRcWQ+r4UWQQPWDt
CCNx6cUBhfcjFAQvm62X7Fbt0ypklFL/5eMzgIvdubxlBfMI9S4Mr4Zvq3WCVGXQLLT/sfqRTuKl
WtwGWQI1058BZqgniEWfIx6q35uOpstekDoi4LC543uohGbH7ej6MMrCAHoBDo++0Zq2xowyclf2
s9Z0poLT9zT6ohWYL577yhCF1AaYq+5BpCxgTu0NT9CSoazgjxmsyl8XpdAh+r4tKBuh9W/E84mW
yJAwh2+8JljPiKjmLM/jlhrtC8jNqRkkYz7/3UWE40FXvbEOUk1XV4j4HP1EqRvWkrRV0pP6M19e
ARPte8XH693wgTdCUjoiJl0KGCm3080WZXtrhzKXDos37kdOhf3cWpsvLO3GHrrSFPGteZ9FXDTi
O/cwXh3gHq5xNEWT+wJ2c8Wb2v0UMbwyfSW76O+Xr5LaB0e0875ryhMU8XruMHU/muuqWy3BsM0T
47Gt5S2UA+bR8VkPz4jLYe0VEn59rmEUXKlmYaRwQSotVXI9LemOiHsty3R24TzJhtA1gTuEC3ih
ipaxT6FFQpQOGGQvjshctrV7Srqlxo+uPUsEJUDYk2SaGWNiKGS2nRxAhksoXWIpKHfDwx3ziww8
lm+QbqMcMRrQW4XyGk2ViDnrng+XzrxfqtSA0leyF/oUyVB/Gbj+MMf4CwHVxzEz/NXnbC5s5jCi
x+/77m80wqcJGHNO6hiX75Fu35TVbOhCtHxdH3QAAq+YQnaEkpH1Dwxk2c1CcvJ5DLUBSDcUNmO/
Oxuf9xKUU8ELvc3dSDpxmLCzL3FFiCd9MxgL29YnZ01wzCIYAESqcHQNlNa3+z1QzSq9D/qOR1Oy
4a6EKdtqtOnS+DHm/E5S4c6ELsXBeF7pjKXTkF9zAKNhW8DtlYqMDRHWihj2fTvUE8OaBRtlPHbx
I/ogbaze8V0czJBv7d3lZ2uMoZ9uBnqXguidNxOGHLhyHMNG+4uLKOeRLS065dBCOX9ZQMeYs134
LkZYvJxDhovhOzBT2bgBNLjWjvy69Ys1i+v/XLGPvaItytbXrrI/WLyqzrTYWZu7qBS/hF6jQ4Nv
2EcZbbaJ3inZ5050KyU/lGdA7+0pkrY0q+2VbWgSCPuH9ujMU50BNAHz8vxakUUA/kTESN3ZFf1I
A2/HmN2/Psb7HIsbRsp0agWWX1Tq7S1CZQhehGxDERQyVrc7Ar8XdoqNruFSWMgg+wtXG5SGP+Cd
Q9mAo4QP4YMseeY7S7RFrtq0p6ZwikFkYUdBEyteYtaTX8HG4TxMNwFkbKXCqZxVnAGvPUFAspkr
5g65U7Bkb3jqqEIuyFnDI4q5nGIdAEK8XInFWabt0nsYhbTlTE9KYGNUbW2JFBJRq5cX0V8LwkM5
uZiUzD+VPSWPw82QNhKkuEOD1/3yu6m8UwtBjgF+r44197jWrwA2yA9cR9P4cCj5UXa7RwTu6e8r
HGYuos4QW1NFSiObkYIu5eFQ+YQuviZBnUSw3BO3kBffEOW/O2fOHmffK6GvN7CpeCFY9vnPH9cZ
j5Sc0Zcx8CtxsiiHnQ0ObxOFiPECkvM28qFWR++YZ8e/hAb4NDiYQz/Cy2N6BSirdyvFKGSrnL9E
jAOfs0wWkW8FUpIQSyK/q7FQQRK/UO6Bm5h02gcAmbLIwouyUURRkUWxCFvNzeMJz3eM3hI/ZXry
SykwI/0JtJHBbwmwJwd7y2K1XFt+o+WyEcXdGJ82VXm+qdKG4jenFP7KFh6C/ZV2Y9EXs7tZfMK9
CsRjgXYRlklbT4drYX4RJoZXznep9iqJ2ZC1o0t4CyVE/mXsvvdntmHOs/0EtUIs9l+a+BjToGAr
uoduDsTw7Uq8L0A6D8mBWr8Hxq8xOF9bJLJc52LGD68nM6PBZo11vmG6yhwxgPb85oFCNj5tat4D
cBqSDgcM+OaDtekBd0H1PFVctqWc5lDUDFg5LxNsfL05OVK87dvssFazDoPhPaR0sQFpvyzidzZi
mN+HEyF35kiFj3K870srHUuuOpelXzb9VwSgKN0Itk6VEr5Ju3xT0mPm+54FBZoqiran6glDGVII
YSxeVA+n7ayTURlPVgFmXHdDezouDXCgWNnhPr3cgXGk2QAYcjJd9o2bWiQVj+XzV1HiLfaLLqar
yy40g6JOVU/5LUeNNyrxddZhnZEFcCXWjui77nY7aXcJbUIBNrhMIiSe5QvaI8Lz3ZamQB2LbtXs
tTU3LJ/sCrgCXhhUSL3r912xOlHcJsEO4uMeNNijzwubPj8kC0r87mCS72kng+aj1U8cF/1SKIfZ
vXV7JCpXCOIpPhVIeQwZ0fF6Ke/qYx9fcIdZKqFuQ6fXTIB2BHc0g3q/CPqqsHQyYFD6GqMaY2oV
NCFu4kdXvdrLYL0PaCJmzbZBmfJ2/tQO5ChHdDCfLw0GvP20i/bhfqHJVyJUeqnias0UUI2LhjvK
1Ytl8sDZ/SYUyxWOEWBGoN/6CswJCR6qzwlX9zECpCdUTTZmrG4XxNraug9hPQmYwpNuAUxbr5BP
E63p6IGQn7uwxEwm+67TXI8Fth/gAbyL9vSLJ5tcJFfjWPxSL68o6Dd9w+IHLNJZlrD+Bfi4u1G5
0Q9PyaJZh1Ex5idlwNREWGGqiTV4nIE5yPGNDD+2ebEG39kKUQAXd6FjpQ/tD9Q2ZhpaUHGdjiD3
L0Bj2c+28CDsQ8FwbIIWtt75uC35TqPGKqdI23f8RUvOvyu2A2d4QTuZ0Q2od+pzIHbJxDTguJ8+
erTEI1uAvoSvJGctjsuounkOnyNb/syv8UNzlHQZENNg/SS+qZTfFg7r/TvEuQEae20Bhoo7HSN/
A5KCugLvlUwaKux5ZxHVPJJT3LBoDInjFxIjiGTv9CuaDawQZmSiPF4e3cyDtADzlDUrHN2+okDh
nhaIuTAafrCm3qWUPbtMSZf8Z28JY36XuqqvbvskmJBKjFS0RC4e/9lFxwn/PRvFQXAdm0GX900t
XjcQBEKNx02eNFZ1zMdjcEvUoSUKfM4ZvI/8CDnTkORMRcjPW/jW7nxQJwT1et59NuHe74s6z9tS
NWEHzik8vf74ZMtwSS+Z0WGUvoE3EsFATLzA/8qeuPNXLzkXpvoFZKO21o2/+xjNWoUWoGI1sS7e
c/NrHFoGckuOCtMTw9w9pRKdgZPSBsPvGJ/sHLNEimo/jgujhrt4AKsCODDf7Q+Qi/tSAIHMINfl
MHtfDsdAObpmjsaJ3WZZsZup9mZH3hZkf7tvoXOJkGpayeRmmXgJzirxIm3i/tirLc5AoDo+16qf
dHsihSbOPJIgLTG6R2qvKxzOru2qYOqyvKAmuLpT+ki+jtWiBPITB6+qA5CThOiZeqBzrkvRc3kz
IyonSn65SP9vgn2yFrIb1Cpbjj5HMOqK5Pm7xT91WaP/a1rd5LvfXyu3fPFvTe8uYQu0D0UkBPiz
12X62rLr4XPbLVykMEr6XfTDe7W5PINJhofq9jV8TiMdORM+LlYO/9QPO58I8SEklFkzDA7/7HYH
X/XtBxTDbna6oQWwM8XFtjsGVx8IHuntHBENWfSszAJVPVlKZsU7JPfCEJn/zpvTaDBbIioBiSma
4w3Yh207iA/VdtCU9SPcFOwrfCNO+kEPTluWqF83BapXYaKIYt75ebFirOhV0emmxLAzLG3Zi3w0
MII3WCLZgkPM6iCrcxrrt/jUinRq2BEw3ZGb3qk4QnfuAUZffCvdG3WbIHC81ShUtrCtEAiZz24t
H/e6CSLEQWACPOoKFUhArP/pwJtz4D0GBMOKfVCB9qVa23OzHPjLtTOqehJ2xYqj6raFDnjI6CO7
S9D/g1Djxjni3ySjK4s1DQS4rEZ8Ya8akIwIgXNzp0oIETo4PV4xYfLiXAaSfV/6oudcy379412l
JtxFpeGgVi0PFSog4GUdUCGProlDkhzjewL3Sc4t6cIG0e4SE1m5vJRZzColAh07dNeJLUZmiP6g
7qshnR7EkLpPGwIHokvijA+jKDd67vv7ZE7q3ptaO/+6vRcnuyfEMWynB6XiRGdzFE7AyBGnSZlK
psYnnr/TgcUjLPBxMdPIbLfWmifwI8X7elIP1XDASJNKp+wPm5hEQ9RBDi93iBI3sDIU5DciePE2
7wbnVz1cwe2JIhYg5UAthQpynN/xE2gnjf60P36IMn1/wH9P/lzv6nFMab0BwC4qfb2foq3ZGKEv
+mHGIW1zrqC5FbsFw4G9NYHEmr+GEdskSo0gwoGbKVZXcqo+FC1sXwG3dZ9B6nDGYzBTGJS3Ptht
FL7U3PjIher6mWA370lEgF5Va8MSoix34FKLEnfCrptVpp470t2GQdsd1GfMsz5bKrcrQSyQrD6p
pTWuOE0jmkh3AvpnyL6K4JTnKvSPGtjtxOjz90EfkcATY0X3GNddl/IZ2H9xIiIVLgSJhtCfYkLf
PGLxJiDz+Isx4YQ3EoyQ05orOdE8RJ06kPntP2lMYRgQnPBwUQ3vVXOY4nvJxVy4q7GPbIQ/Tcyw
TQ0mg4u1OHzIpXlEGc4xqTCHjefLc0pg9pnSQcUQmWsjOBSAS4P0tFWS8esH783KTrbXUToKLapb
f4QVXFbSlh9rE4G7SiK4fsl8Eb6QNPkuyTBr7iCic7qkSfet7rjcJZBBj0QdUFsISZjNQMn/r6GX
OGzYcFOVwzsu9BUS+019z2QmZHlS1NLzckuPZvF6E5fVkwdaQI0O4Sz7GsM9zmruBPy6J/1254Pf
EbEDxLlqiaDzz0+hDl/6FF5lKQZHggYdcFg+Iu00QzJpn0UxV6FlC+hC7bDXB60ev3yAEnuIGgfB
gRVF3SSawY6ak8947PpGTRdkJzaJt0HgSrPX8EvxpXKNXRu1hBhA5K4SLTrrI9/XscVSaMZ09y1S
i5HebXOGWx5d3QpkgQkSUjNU/qgse0ic8OQNqmLkd32kUGWlWI2pDGdC1hh2Jys8keLqasl7fqPC
rD2esXq8UZIeUoklM5ecy1VC+EMadEl1VpuiJWvLXeGhbXTIsOg/+3ZlMd/+Ic7fTlIeF5cayqcW
DadARowMzZp2OjOlIpAr02jRN6XXNDSqrHVP8EP+NuVY2OomqXJjiEd6heHr0mBY1XrfKJLLyjy2
Aq7Qj8WJrKLbvAP3hVZ3cntfKiFmfVdxDqtd65oVC0AMO9KdMf9IqOUO84yLblmKKlgPUt8SEXKZ
0/rlFEakENeynfsJ2Ct5mf+Mh15pzkcCb/2V5VmCRgpbw4sKwwlTX9KwPTo30Y/nWVf/XTZEwdN+
gj9uQmU/o1+uenV9UaM9bijyWy/FUhqsMTcuWRsknVpOAv+7wuk0Ia3dDQ/Ofa7qY4PNO5hJisFN
m2r1g5dI9fZb84it5zZGxMaJGgOAL371BmOKdE1adDUxOoT1YgHypdICoTjWFbZp6IFqY9vL4I3I
3tNO7OiKvEB6I0KW6zAudInzO43ene+xMb4H/866v3EDTtfKnLVY0bKaQYUwsEcg+gsXt+PI1177
V23NylKQO3n/s+sPyXQs/fR02dBByguU2C2hjV8r5AZd5wHYan3feDgj9m4gpfkQbtseJgHXE49Q
kYvtV9xRs4uPpHjjkkvNjrbMGj3PCAM863NkbR251HzIgDiT0cTgyrB627SZKEpMPkN8LM4z1aex
+jJSn7gwIbNKVfxKsgJfIM/I4Lhf9xJGWRMjY2EfqX1BDA5jIzm2X9bKdo7AC3mqjxSwrCvk1Os3
WtEqH345xFx5FWETFkaoBXEgsAsrevbr5DpX671R4OJY/2VWX8xfYbeOOu3qo5e8v2CliXkDpzla
/g7H/mz3kc9Quo2aUyJgDqDL/DZUjHYba4Ulygpw9KrPFCgi+BH9g4RPHTimVPww/qvtvlCbnQIR
rwtYyk/E1gEMJpejiKrZyng2ds+u9RxWRj3JaCG4fGwduzX66xEvGpaiKrXjhBfRH2DWAcK58okA
uIB93WLoWGATYyd+9xHinWpcr7Tr0J4qvKJgobGyy3NfMt3TauPcye2mYQzUUO1LQnj/+xPzVnmH
JYLFzZeRqeTEbrckE2tL0jYL6YUM2Stceinb6Ch/hAtpp90oxMVZHlA0NbSeudT+Y4HPlOA9k52b
+bv2aZ1PW3cmk082jwMGsSW5x3U/3O2DwLHqfKY2/K/y4cM+fCU1DS7cnV4PpMMN49tUtB9D7RRk
nzhHgCpUXSg0QSRnqtmOoQII/BMB3Q9Z8dER3RhFMLSvSlPdrE5/9LYe3qpA7Bq3IDBKPPYe/HAa
2xorKBy9wgbQ1OS/0Ss4wGjU6uRz2v2MdQM6TtCYXkfTS3aA0+SfPDUuolm9OKfvWlWnDFWEqpr1
CX/1zvdDgSUfYknp+LP6c7YHERtj7wUtEG+mZ+QvcDTbB8K5LNNnT2xUT+rgFndlfNanEL97Yy0w
cA0DQuud0UA/KLIfhWk47zgQlgSIxGWgn6h9jrO+j7/ZzzKnp+T5ZEMpvzGgVSBqUWflGza9pk4D
xIPPhMUwJL8PwWEfaEZeOYTuMqJiJAfYF9oysTeP7xo+JqoDm6fPOrk6sJn/XMbqBMNDLJQ3aNxx
KDCcSMTsfiKHu3CE4NiW2agJiDCZFVYuQCh3f8lJuXbbUdQeTSEaV84NGGdrJ72FFYFY9F5vts+q
/xid2FvkwC+FADNvBNVkGqsvRLUXViy1OlqPTcM5+Kf79+eo3eRtBwx3wUiqRn/CR03WS19uHNUx
eP6jH5CdQebO5CZR1tGoOhwcREXyUC0LDdjTumCgjiVvJiGX+DwsiQas7nUTA2cFnSbx2Af4pQgJ
mgoSghW4Zp8Ve7w3otQfu/vOjjTR6/DQbg1ceJxeR1U72+ivH0Rji7FVzIeOF2UGu7ZKIPMPd03j
8d7IkJFgddOuJUMVbHBTAdXGHcI+E1kMN5daK6xu8ju4FyHnY9OmzSwMtvSiSQ/agzaCpmo4z8S/
KV9EC4uaQwFLBlSp9+iX+v/F7DTS/pd+K55Xq/pumqus/+Cc/cCCMxwpbDWTwlg2m/Gf6iSKm227
Ai7QRCK4MGbclZMl/E74QjemrRo+j6lqu+uZFxWik2Ae1rkudtq3TaDSYbLm9zNhh/b8C/Ju4ru7
ebD/PvI7UcIl0khrN/ThKPRnqFXHbUurCAgWczLzlOHB3iuce7F9WpzSj00Y8+Na6ms2azJY8A6e
XdWp3Z2izgA9LKEz4VYzAAwu7l+QiuYnLhsPKq6plj0H0kNPqA+Gj9PYyN5YSl6AF+8XMASp1YpA
O3Z2MgzUKa81h/U3X/HdxXmu2lFP0YRshMyGlghd0UOpVSC7iwajrHs4kJzH3hV/pGyHJYFV5pzy
Aclt12p/MGfEDRvJpFGWCqDqrUcEuOBpMm0S76Gp62SWhacJCVRlyDkpJyupH8ouxzxf7SNQHoT/
Kc+08flBbUoMMq6Ln5iVJQ7qbDxq83hENvKI6LvxkFCcJNIpzR2hYt7w7k3zzVtIpzpK1xtB0GTU
NCnYp6X/V8aOThn5ViRFecF4NqBthhGsGwYaD7Z7le1/VU8Ime56prdAiQxECbmKum8Syc7e3RWF
6L7UyPk7JsqU88WAW/t8ueRIsFevzfGYcLxuMOX5IRZx9mG0bjL9nTknJlWTTJaGTKoFA8o8nBEN
DHH8lngydBpSxM+eYSHCnfCNP/rRseNrjEZ12MmNDlQKZFGEUWwpjkjnAcrKNWemiD5giXnOILT6
lAAJ0P2rUaOyVj3c63fJow6ArvwuBaivLDRVyF5MN1wB/7V8lNbHGprBDCFV2EZKcGiAGXWv9mFl
o4lyL+xxzWRoeqJWdOk5auKk7nIdz4VquwJdgdJgHZ1cgWNU9DA36qPCdU47HhMa6xxsDabdixZ4
Fs1W/vqOa3KOPO9NdjDeqGQai8QnytDjtYVZTjkLkUF+7xfXd/k2kiAArY5hDuPAKHetBgs/qYR0
mngHtEkSY771Ei7vapjozR95v86v+7mw07sOMao9a8EzY0k4yJyOxrFKQwIHvUT7wnbOc/WPp7pS
jGZhppunrFOXZtm9GKsXx0/b9toSIzaPDOk12ARLFQksGeIfZtAWXpQzbtX/csPlRcdegmKuiuvE
DhHJmt5xe19zdGVLvzUojpUqiZ4PYt4dTA3WnROxOd66jPGNJBYfqziXtT8ZCN9zisCiFb15RUNn
W6kHrLSwsZaBrbBWvSWwrSzBveRosQSbmIGjC9apQRxX3OKeJaa5MdOniHVQwwFPEKJ2pTZ/xa3O
s8PFkjISpqYnvrWTqJby0iG4QbblsUxbQCs5Qugl+IquYN17kJSahHIpG5Q4KytKekTYhwKXcalH
SPZyiY4sq064qcZ399hSkcY3MwlJ+tgUHvm8MvIkq0TkAllV31v0UFTnVM9KX67wlspmndph2Feh
J7Ww3cIEkLJqCLs3jPfOotC/dAi3hwm8mZsMF/aAGV+yDZjSxaTvbMBUi+d2H4jw6tPkKEXDnjvZ
Wc4QyJkF9nTVUWWdRpUZHM0Xtyn94+Fvjola0jhf3gFxIXlZgWQ9vBs6Wb6OyZcP8s3NnOGjSfJp
D/CO15ye7gmfH6wPVoP7nuHfa32qIEh1fPW8KKrFf0yq7f9kF39NEYEVA3eP78/oGFmdsdtXY7eN
ANoSGbLZviSxU1WNJKa3jaRyq0tW59jP7wnM4gtAXQsrsZ/rl/dKjzW/2hkv/whWzGy8zIIAZHxI
K32iYO9ETiT6jCSCI9p2LSS5oh9dhn+s3R+uaFd5nnfD5pxGB+jYVZIwGiOTqLpduotZQj0P5ANU
DuOx6B0q/ZP+V2xT7E52eCA9YvILDt9NKIXY/G6iBOOK6KpT7vtabyv+93YkOT4Q3DkimufR9xva
wQYqtNYIrX6Ds2u6LA+IVsUvOAmBFmXpArfEvZ22GjMfbXUleEZGnQU8q4jOKto3IW9oep/wrSdZ
kCgphho61cNWNkHnNGSm8a/Oy2fk5xtbit9cjul1ONCYtAuF6tY4zIbP9JjH19+FKc9hgiynXc5W
qob6is9G7aOXRHUx1E9APpjQp3XY0+X9hHhhQOblUgeDl5bGi46nu55eXHnPxA3fV56V1ZVzhMqc
e4qsKT/Op+xH/PzKylcWsPNlz4T9qmzehTxzKkY3qBUcNwYM1Hvhr47KD2JAVdIu/Zgr0Gvm8iGi
hYbLkwJ9MQ3odjy33ju+Y26URyyOibCSHfDrRYUDg/ZJwXxwwZHhLu/0xD6vWEVzbaStXal5JpQc
Q3UW5GoZZ9Tk6EJ94Pb0GlCooFuPWM0hVc51zniJknxmWubTb4UzqrKC3q/W8cTNPLnAQisYB+TI
C0qABTGO/WQdixWadIWJ5EFfIs23Kikv00FUsGi/aaif9fSAnGrIq2WQW7yXvMUyY48XMlhQvSBA
w/GSBRypTGDYkvEPVQyfETBNHhUqBy+OIE2+ghYVnVU0S1H0QvQRA4Vx/yH7NZ/TH7wVcETUnI5x
kf1Zpevwa2/EX4o+y+OHeaE2+DcmQhyco+3aavU1JByaqKRU2nY5SLnngog2WrDx/59fWLUpisfT
RRWSgK9CT6/7Kv2iDdXwPZ4sSyN4ihFPx4K0zkSrKE/r9YWq9OKSjqu+CzmEB2dDwwKChu4DD04P
QIPipdhc7baWZkKGf1oeck41hSDo5l12hhcZRjen/lJ6eHJirpho2JccPt6xcy7BVVY5yFiaF8b4
hsAiXC17zSGkdu8Au6Z13x5oXG0ddPHz/fCwvyP0/mXjh5al9FLeemMVSL6a5r23sf7lQPC1WOEg
Zygz4z+XGFzCEPtK3mOfpFOcI2zCh3/SyyUdEi6WeK4jN7yyh6bsr5tRVwlgzKs36wcwjaQsixUr
QXDUcLy4q15n1s8qh4lgGAXD+u6UR1DeB2se9rkHu6Hs0uShbFssxAOrycq3UJVx9UxO4/AJfVBb
GNAX1+6O94m7rEWfTu0+dqEUgF81ajs1LqsQ4fgY6eN6nmF9eMonHaFjfayK+J9N2aoDxqtARTDq
Tw21nwYP0dbXqPIU6qtEvdSRQp1JLIgKsGDY7/5j1RMImlwzYZ42676UzBOFazT5ixM4K37NWNhS
Wyp38TzjmgG/TRTgfMfZGlwvSpY3I1gOvNftn9fI8L1N61HHO8ipneRfaAam2jyIqnWkVdUto4au
KWQjOadKhk5CmQphNTDvKfG7gN/PlZkI68LWvRfmm1UE7/D6e1IRQfdm94ygOScxx1wj74a76faj
UHvjpwkTaYEkl2RTyDU1nraS+byv7yioU88vtVxkzxzES82JEy9gYfE79JmILGppK41ams24dBFx
ejExoI9idq9jwh0OV9gR7Vo29XK/Z7DAPTUaivdlwaENAkRodW5rERyZxCkI0bJNUitxjU2p7BuD
9z0aIw4OXw2oYfGZy6UaDJiVR2cFZbzeqQABH86eKKH1BhYKwnkvDfzYwfpE9vSb1MlCG9zSZJTT
YItwV/ql/JTxyZyPtABZwNEMGytzwm4htiMu1RjvZd55J+6NSfh+xVYqVsD4vS5D+xu97xo58caA
FM5l8P+7mZ9YwozFfA9Sl2pv0YEUl9WDdprw1seMTLfI0atGUxpz1zX9AU5pMdJ2XbxNbD4YMHXF
1S2aelzwb4/lfQfyn+tPS4MGmG6+pBPvR6Nwb1xTxPdR0yHGNgkufjc8nXXqpQLNDmNkJLLdrmzX
t3O+T94SR3w0TkXsZ1ynEZEpzdtFFKtH/F1za2xTZAXcGl2VoFA15u2v9jKVD6ry7SXhw7jyLISR
ucJqLf+Akc8mWGpVQXM1WP4LdgCUWeX2Kd8x3ZWwzelsmnKvx8xRq8OXDC+tidiAqev1Aam6DSa9
IJmor8IQDsCc8KUEab92KTixygBrjElg+cwGQ/90bgucQzSBbrADjpSM80/F3x/o3IOKGc6danZ+
Mwx6ni+iHrzWYGiKZgQmTCxtWftmAKVgKBVyvo9TmjjBvjLQ+TaaNhs80GxNI+pQNJmU3RZ0WZqi
aNuB6ibQQY0WQRHfhGLFSNhy9OJiPK+exz40gS8uy7IdoMPpOi6+XI+AkFWwxjgnTi9JLzoaTBBh
LUpBf/DwUOq7qxltZ69oSwNzBPpFuhFgT7W6dan4Yjl4SeOx+H8dyJM9un/tBdP2HdkCpd8L4qX9
y1vhZnkFOF9X0pkHwof4W0+CFc50ZgoIW5KsF5dpFRyq8b5E9p9pxrMJbMJPj0ozJfiDwBEB8ylh
ZgABP6sAANxrNli8hBEDWzkDfM8aRj/5EpTW3fEGVl62uxrATO9tL2twsffWJV6T+9abvGUZRQrE
dleAvytYXF/HJyfA2gvh9ZboXU8Shp2g6NUyB2LLKeYhh81wevs86N9ClWTDjkpTrembIuuL7jyc
YvvckEnzpCG72blRDewNoG+EMznMCr0ecC1BvU7CByzSAyF3xrd1/ueTpvDckIZphp2ApVHA1NZn
e7+ak+/FSg0gsyLCmR3aKcVmcnBlxHEy0jiSWo0vWcc/oIDLkFweA1IeEDLot7zi2UIyO387YUIZ
19XkPOnURx4BbHWiGemeyOts8ZxAWynhCbfV61ayGy5GdPeV7FC5e1+Tr94BMW70BtI96XNCp0ru
1Kana/J33HDwENeAukKpaYblMDpOmrOicUKFfuehy6Miwm+G61DrTVgTkwDyYriSJsOU86Mr065l
iMJTaPpBL574w6StD6JaIM72ZjDtCWArFxRl2GZHgo2YeHz0u9FfBMzJ79r0QnBp+76fUzvaY5Lg
WQQG8L+DJfw6GLkaOPN++FlD8FU9W6aTpyP9XeFPxrThUQNM9BgSp+Ucs+QwLa9kkIMEPsv74y8x
73dwnkEH8efMh+YvCalR137vp1HqABssaT1JvNkevTtv92PJ5kQPnTqRJXCe4mqX0ItSl5H6nvVT
tyDWUarZCqg6/f3KxxyVGV/eiQxKcFAy2Nj3UVYNwQ71xCbUDv6TtvlRwuk+24Nu6wUmXUqKqcMr
mE7ls6W708tT80dWj3lxMn5cDtAQRDP7yFWkhrDQTGCFEVGsKiJvRfoiP5fPU8bQ3hbIt+3+hDc2
rIOA94mlPsajQbm8V/sINbkfMv6UUPJXjmUhC29BlUIrKkkhvNN/0LxsUSrjlHCp/6xro0Yaa3dx
MALHnPV/UQDeYKAyeMUhCXzol/nUdeYA9SqdjrqjyA3MH+bI5+TypCOKnv82qs0YKoC5gHakh3SB
f13FnNx8KxPeqCPmsmRP6aP3FqYod5GzEImaTfNnjyDbm91QGMtZeTA4r5YkqlZJ5ZiKmrsXnN3k
p1rOPZtwPC8zB0aGubkmkJ29f5jVfITPhEFfO0uTbpn8zb9zaoogpq2zPIz5a3YuivxOVgkfbEOG
tFeKOVvPvFkBQnW2QK7dUTP5zel4IsUi5kOrT+3cW72Ybb7oXZK2uVTcAcGjswFVi7MbzMlrdNTZ
F80x9GAlEExy8NLL6SZKlLFfmpkpzcptk3aazI9a3N+pf63jjurwngJSF2B/3RS0iIAGHNEPN2WV
zvz6b4qjXNIRumjqxKpiyAKSTqjzw5iKvJggiNfGXjgQfHCouOxE1TqD4nLcw/Z2OlMoZOYdxv5P
VIqvouWSeM8HbUuOk1Ns+MZ/KeKkTi04Ck3Yu7QTUystN/WGViEKlQXiADWMi9OXTiSYS021MdVj
+9cytxQW49k6GLbfBxdWi/JEnKEnmPKZeN5e0ntnBmw3RMyJJYKY0DJTJZ8ppVHVuw4PNLFtoiY2
T4VPTQ9OUXgY8JMjJFp6/GrLp1pbGPTdCT72tlnHhL+ENm1QdBGSjaVvR0UjzZjTm2Ke4eYRcqxJ
odhtQ5vq64s8p7yIERM1eKhtIv26IdxHrmtlxEHpW6g0E4ZfcfU5SrdgKFwBeQ4ClfWsR0uE/8jD
TDNhCtXth/bwPzC/DMi8xKoSeVissm5AaUT/7Gu+wYCoNP/rgJKj7zkPwhS/R9zSDnooMt+PHS9v
1hMfuJb0dUic0W9J3dyPPTVkeW7MFtqS+WeUzdsKCAT909bkKmu2SdpNo8n2PGkxiVZuycm2jkvz
p16j9OrpnlVudnJDshwQNXXuv0QRb2vOlp1KrfkDnONvjSIGn6yXgKM6VTQMNuZmwMOZYEV90Q/o
+V1NITy2FBH/uVDbXd1zJ/aRKOtiwHvsX8Hx9Rl1Xu7z2ERBjWeVmm3WxdNDKSgyz4BkRaDo3FVg
WI+9X8Mwd9dYgI9Zbr1x6fmTRVZChLF0QKnCtDuSpJjM8651PLznobdo5x59/wA7vPQGD83nRiYl
oMlePZfqeOif+EzxOXpcrkHg+0NhUx2gv3YFp85x9TPj/ptu3gCiDh5DEKQ8UQm2DkC00g31RgY4
J3MmLo528tJYwL9XclT7NqdePobg0JenOaxRaXnORUSrIb+GzEWyC/wcdNXWLBLpi1sGgvK47Uik
iLZfWYP00x9pDdF9vq7vz5ur7hO06QHE6xlPFU4GQ9bbtCZTry3CAx7tI5IN8scjr0sRGb3sLtj4
yK2A4M6DvkztUpeZEfMRF9XH83lQlNPuibuwo6SJyxxOoNR6wib0oMhW8TUQAcjDYOs5pgwDwHDs
GPxBiz9OFoN8Uc0WBs/yuZCT5LOOUH1ytOKfjK0jFsR4bmQRpT7YmgrLibevaMhNHBXDRJg9KTM9
dN5iwEspLVzTuG4uaozEI/AuahrluajGvpevfTYffvuf3sT27bSq36fUlvr0487ZKoDs1G47qlCY
PH91HvBMJLHzOZL4GDz3+QYxy9dujlIScptxhvX5u7xdMJnZEVlbl9nqwEBTAC2CSJ2skXzZlrd+
/3Fhu8BRGwftyzlWCw0xC0IzvDxlIY7Z4T9wW2sYoxPAd1TG9Z0vBif/pwdfCaBS5Jb27vwUR5xB
u0yZmjCciaZWv2JntDAxb82PCRGQs+YMDdVFCBBMC1V2tn7+Zw3GvQYefAUuRKP9iFIpuVUmDksC
OCNZCbR1IMcQh8EUJk9h9IGAG5iq62TwFt8y/m15XpJLLPNN9GSDTxZoaGCBb+pPIdn853Q0AEcg
Rxm5YMI2R5eFIGOHt+5+K7OmglTEkTvMAshR+gP+w0bAdWm2jPggv8QtXsKF42RkNfSc3Mm2YrRM
DK8NIQ3gJsah+teobADpW3ZdZmDzt5JLsPmIP/vem/bQclVMqUfY0+plv045yH269NVT9k6U6qGv
JVPhGd/ndiKLHdQCqwPF5kHcP11HMqYLOOMsFYXr0QR/+D4gM3rhRpPsoIVgwcE7qI62Bi7YGppg
Pt5u+7GkaLNnptAuENRZpU0r6iKO2wa1TVxaeh5hfww7fwVXNXur1OyaCyy7UWakR5eQt9HKpR26
iemktJ6p3wl8Q6kkU5fkwwVnkxASLFkgM9LUrSBnOJH9wHlhHLMiyTy15Mbdi3Yo4fyP5/K8t0la
c5voNKPhs0NuY9GBhQo59kQ5TqsyMd5IncIXh6EgP10Le0mozSDSwp7y1lOXfa4bw1Uqfyv5aDbe
IrQUlgQtHwDoGVNr+8/nKBT0IdUDum99PF3gBg+nG/NqzdoRSeWG0lEdZTzeb377kz7YmJ3pRYkR
q1uiqfkCTOiOyO8X1Jv+CWAomLEM4Ix2K3T4mcw/fIqTGrfIHE+n8j2Zt+bwwNN0ia3rvKn3XD/7
cWicS6y9Kv0NFpATJSaO+pS50j0F4hHD5XXOzexzu6jIzcaIr+zeeqVigWKT7rDXDRR7gTbh4u0R
i9CIaOA/TFplBig2jvjBp6Id79KtnIx2NiwvRklT9c5jNr940YFZqoiWCk7x84l+Z912NxHD7F4w
eo9YEynvNUmwOm/7q9KcX6eSbD+b/EUqmNzK9eeC+KMV2YQsBL4DZ3ILVv4mVymCHtc7JUEHpyDm
TD+NtHLlRHA5Asdc2pJ+MKl/jhmuSoM/xHmv9iJmbgDazVoVV2N98sVI6Md+Z2l/abNaIy8SXAUw
XlTPkKO5ZQG3d74o/VbFVp/IOa6eWI682MB/8fTD+aBbqgYiUzgurF5qA+/opUTR5AdCAhWNDBfV
rfn7h4AnjxfyKYpQPdig/eBqnNvjT4/7sEiYxro7wLEsn+v5bf+zkcZYsJb4HaB69RsEmziFDaRa
nh6Fe+qWPhE2CtqhxoZksACWbH3nhOrw5GF6F5FGYC13EkDosGNpabRI7NECioaWHXpRbV7tbDmZ
h7+sKKqalEsEBKPHU7s0sAEdqp5BxU4o8wtwLgF7Qg0hPSDr0An5fS2ajLyhKouIh06BTROQQm6y
2ycZ5/pkEKEV+raHM50pdAHDUq7TTTv1vGXp9+TgMKVHJ9Cw+lI/mfVTPoQG8jhXCCu9xM0l2Au5
MGyGAgEbWm/CikrXqYxzeGGCi0QA27L2MzgdkTMBh70oY/prdE8fN39e9Wv+Ni9fS1BdUDB2++gU
BECal9Q3wFQakIJnJn/BRXQ/IYMfPsCam0Pd1c/CfV2taZlTdcyRqcQoeVNu4VWJqskBW3LtEqyD
iZJRym6BUFt1wZI8jlbnX15d+TnPJEc9sa6hByE2fQOgsYbAnoe+Q4/tH4YmSLsXod26iQdQ5Rd6
Q2uEtKZgbQL4tpiJzRHyr6Fl+2+9PVmMWqxQnO4muXwlUtYakEf4Eguo7ni5BBVfJXpgK6Bxzoo3
LIWlLicQ0Unh63saNaH84M4nQXnSlWVlXOmUaAj+9gCB3Uo5eRWXVae0kI7L+2BXpHVtpI6OMRqg
+OpLfQJhr8r8JToSu0wJFUuUtI/RBrgNqA2oe2S9NdIPzu39J9oQXCoLHhcB2WG5D/ofuHw5dYxX
z72uZ5ywbsQY2KlJoOlUUFjsX9uX+PysWFZLCm3D+dikZqrrJRMnWX1E63FVuvytpzX2XjYtldxC
xOmFBgzRIfrksIdkBecqOOXeIM8VoIsUXleqX0/Cx/upMWeFz3wBq6GuggutUozk9Ri4T0K8FPjy
5aU0SisCdvYE+p99WBj54jrCJVHcfKp1sUr+FISor929MwvTpvbblU06RIgjT55cxUQxZGymeQa4
7Z3SifDRSLkl44unq5sfTvSPGkAyoHEHKmTzomFJPKbelx0lrQl5gt0ONMx2a1GA52zAeW3PxIYh
wgL23jdVWjjqjim8ax+oVajA6+WtnUHNKyERXeW3pIoRMI1cLD6dNYivzkz7ZMsWcd3Zr0xOVVum
78SJiWVCF8kg4ZJue1b0aC2rTyfJruJ/Tm3sxjCs8tFfqyuMLiITqYrwajYVy6g8TpWb/ZHhNIpO
tkm9kjItiXpTONqyc9Go3+w2NLWINm259CM2pnPstFdlOuueWTIcW0bcWJ5ci+m078kr1RPq+jru
shE9vGW6NEqQnS8RiBm0ThlHwEz36CtQFuC17qlpiTns27+bClDr9OEFgYK9TTfQ2Lm+MOoOtqpi
YqZARuLFxaoqUJpCKQfdpgVHECevsD3BqcDbwjuL/Y3qiBln0TckqVH/6qimV6i6Ctm76S4Pz+Qp
7RH1iNUvwYL2nlU+Z4sTq3X+T+Op2HDPQkz558M5jPpMH6Ls20fmLD+jD+CrcRnZncSOh6PDCxuJ
WptUcOuQSw7blod/FIrRUvYhE439TvAYxfHpVX3VvfrywBwfNptnDs8DSyyszVNvIwE3wgTxCqv+
zxkcMoIikEMSALoHWCaI3UV9N7iWDkZ7soOmiQiyr6hxnyAfoUdjsJH8bdmZeex06Yo7SL7rtPxQ
aw9YpA2WtcMDw9udmtt0ugsz6rAmBRRvN8YwhnWgUBaex30ZJa5M4P5HCmo/En6dvglGMS4tnsVB
+ucZdpyhnKzls/LifGOqZLcZwRSYNZtpRCNl+C79qwK6BrldPoHAQfTTJjBS1juaddDORRqHKs1r
e+VA1LZZhZXZ8tvfaAWkdOLUpndSkSyK7EBTQdLWXg9bk5+vlaUWOjVdzjt+euJvRVAzepSMFfuk
shBzBOqpvLAc/3QOTGcAVrl5EIL2lFff3mGev2WBi/A6Jx780F5EgYYqTbg9Kl+iIyWvUo+l0R58
Pbwws61+fNKVVBI4zQZzOWf5y4aeJtUN9INH4J2BRt8Bg2MoFstvejQoyB9NGsbzgiSMXiEk6K+0
ZhU2PL5pCsfMZgEFRZpvtvsS6jWzXSdSmiPMzU1z9yixPab0gBM66CD7nO+QYXlhN6ioY/R7Xte2
NPvfys30v41CYFnsFO5W665VaIiTeVptsv/+5ocBLlkFkvxBGU3LoTodXRGY/qkJTbdnPuLh6/X6
Nv7dUjPmri19sd59/Bo/xkB2Lql11b9yiEtt2FfvKa8I6fMYo63bWbrRNOOesfmBV1dPnaT1Tw36
bvZSRvspGb4tSdIgEcyKgFAK8rpCrbATdx8tdsYuX6u+QXhQSX64aOkypVqSlKkgWSffGo8JIbGB
mOloG033U/Z2mKlyg6w3GHAF96JiJB3pymMA1tCPjUwtVK4zpq+Xu55x8J0QNS14xIkN0dt6EyP2
ZfYiNF4RiD8TgHCasmU3WweGxSC0jlLXuAZyW7U89R/jq1SrH9G3rxpp1jeE96Hg1PFZQ1PlnDi7
cEvmz/zZo1ASKQ6Qicj4dpwOsRSC2kkaFK/3qHq1V0/n+DMpOAgAt4KAIu9smVCianqTUG3cYJK0
r0tmaBKiNSNSpkYDLxbcETAaFaQQ132FYTo/E9qfsjd0cPPud1AwXvRky/pT3qhQmz0e/2iM+Ec3
Y5rMtf9L4O9DjDWEeKaZ5acr5Q61jFGErEHMdIZgcZc/4V0msZI4QW5QHJYPbK3yr85s9PiWKOLf
rBLGIsxIJ0JYjxUvJQqlso85gWOQ6y5Pjcxq4V+km7TkUe+PKK+d2ZGQYUFP7i0Dhh8IqLqp6asA
9w5b98v+gPfcfjDASZwG8f+pCt311+RmanHNdW5UTpDOACxrlkCWssInsjKKVBPbaUD4oUrAXH9m
ejD3ofdMF2cuYkfNt8VDfVo8eSqwF5U6JMYFoH5UyfU6Zdqv19gGCI6wZoau1D6ohuljEzdca+R4
3La/MhBHCI3ENB5VJ7VGdSrFoSYuEferj4g3Z64dWGV0MR86Io1Qv3NAwbpFuUtM1/wWv5jjVmSL
WroepF5ymPjNXjhCOhSkg/frHsskpXkqDbaTDuj62hWJ+WAc6MPs8rff33M6Lj3fEoNLupuSaQG/
ruxLVN6YJsdN1bsRga4wSsKArzCCleIf631nEaS9psGHUkSuVSqlbDhzS8zSJVnHrYMe9msAQe/r
B7PP32oVnq1/7pxgE9/BS7sDdMSTWL2hHSVPU6N7PtT+RbsGXlS9qujnsGJG/3aILx94KlgFoZic
ciDLcXPPzrE3PGa210HwX8X6/PKBN60ZFTgUqHekldLIfKb3/per4H+84C+yR7FHlM6HlN1Z2LtF
eeOa3HQ5tJDId4sQKllwZuE9FIyPaoefF9PbNYi1U1uCiFvYFHSwYzVacAtktlSHzS4IlfMnl/aS
1WtaUH6+zeRBGCiO1BEGnsxK8ksOwl+DNZZNtLbD1rWSgNdHYquPDLDQxLI0E/qyW6JusaU+yf7+
QhHWagrVy5jlgnivJKA14q9b46gzmRNTp7tKVQkGeTOyvZWohtwHrR7mdnn/VpXOTMIL6ycMwqiN
+eMYbes4tadEEFYFuHyUkRP+myjcDOKxz9t8ChDNuDTm1RHtX2SeMqYBkxcnIpe4n4T0orETa16+
i+5ho+FxfVkTtB43vUqsF2xpd0EUZB7WRA0sky8MZdSZ9RZG+n1X3gAi07MLgzh0kLRq4wst9F3N
MecqmUMvafSf3hye3VmhLk+RjpTuch+ry7BSF0mDPU2kdhKuUpeOo1Udaa0weBbe9Uy64Xuab2SW
sgnIAVx/iGHS0DXdj6Vwr9GL3lFPKv6QxqE679izOFl7KPWxCatgUZ0St+wiyMzyR5buz6d1O8jg
ScihOAxaast0tqTD4mb5W3McbYTeQNR9MoA1l7ElNKtw+qFhi8/QQMF8UQoq2Oce7r24f6AyI5a8
9ndEuiQas9XTZZLRC5lalWdp+dTncyidBF9AQ4BReldjiROR+dPbm5jDpy3+BsjwDnK1+BYwguaj
lqpknBUEsRKb8VC89/XpV4IwDWLnXzAiWiZhXi8oMgqlDA/svlOk3M0wolMoAW6c6i//adzbDfDo
xEtirT1KYCj5UU7S7vRVGdr2sD5tbNOe8q6jlpphx3aSGHZ2h+kE4QWOoMfuet1CyJN5V53cPBNG
WafvMOScYJzFIBqRujVTm5gdQk2OOBUy+nVc8kas9r0x6J0/1eNQGr2e/NDhoqWlOiDw8Cq6ngz8
d1B98bA7+xnmHiZrS8utKpjoZgCSByPE0z425Jget0rK/QXMZm4zNli/XlzRiD4P6yXuMKDYZZeD
f3qgjEwsHrl4st0JaQKIejWrKXK4kObuWf4RbVZ6jTLPPZ6XrQm3rOTdWU24asHcsesjYCm1o8QB
mq6coCuQZthRt+LUcJMI1ZHJofs88hLptt4+iq+zQwpF8F4embvqWK2TW28FEKDJe3/ZBBpOrSjK
0wciiURhcmoquyDZtD4hNEwquZpNKYO/fNBqZF1JOIPAzmUkEWe31tWvD00lF5nFNsmdERnNirMQ
kjLfF6AacfvfGD3syasIZbABoglW9pVOar5Psdzs6wokhvzLnfpjiRVHSxxKYeuHDRGMNWdN6dxN
ZSX/6JCwTpil1GUPWJXJznhg9O2Lg0yChUUtvK7Z2V+s0Ng1mDBWjlA3/685vS+xHE7kJW1Jga8v
+b6oNerl8uPFinYbFq6WOZeugv1qG+fSaRVJ6qOByIifqWjOm35UDZ8k6HTXC9GuJ7u9OGNvMdqL
q0NHP/PFpswKUW2hWdXrL/Ueaf6AST3H9xtWL4gZoLT1ZEzrHcnbr3IGD//7MZpvlD2607kgXSJc
foO72B6Q/z6WNfu2cndVCJ6fUh5Bpngze3KB9HRwb0MzlcU8dGo0FDo03yCkw9M0mRLkf2IkW0NY
fuYUQqnB4jFSBgdLv30OHu/Cto0pWQa+Ge5YsvxydhUi7A2SzwpM/FHXqN+9aPDU94+MD20hpQto
zcgAp1l3Y8/ZuyGnXGU8cRTQCQeCJfsNYZkzsl4fxxJpZuo0PYA5hGioytSMZE+bOGGiULQ8cdj1
FpXhh5jnOkU+9GsvkJu4jzz0pC5/6IPQcHO/y6CM5vFMoepSzr7YuoTss+SWwlfuNUYj6ELPkiTD
xS45gWakpKnxIpW8kAzWkodhwNorFv5AsVg2o+nYdX5yDNbtLu5tb1v6HzFK+0NyUHmR82IN6Vm5
nGtp1Cbhg0G1/fdArAuaCulmVgXsd714PwPxJAe64ZiAc4VSZijrw/MHz+gmxcrVWhtwoJV4/olb
DMVuzlFBkypZgvQrddGownpLm/OV6+pu3Rpa+hnwMKZ7koZq7+DECmetUmUa9uKwFEW3cL+Y8QM7
tr/xAMOHu7U27DWhR0Ww47DLA9OcXPBMb9rZ4R+BFKCLvKw9G883VqCwIl8KGM7WN9NfQx41fJnw
t3VgL9fM46iz+KiHTacLtDKgnUBkLTUe2kKt2qh0J66OnJL82cZ8cUYNRfwTAzoh06Rd3Gx9qkpA
cSCu+5KtRD79qHUnN1ndp27btBlaTbpG2UPgutEwFCj0TcvNfeYjaTWJQ78Dt4GKmgwmcaaya18J
QC4h+vVisYollwJX6L3rgnYyCgw2DdxRemS7/pl/CAqMlDK6qZDSk0P6jntfda+YcOdDnwPabfdS
6/ubG+3uqUJiaNAirSQvGKQeVIM68lQ9uToerWn+cUD05nz88KYtu8v46t4LJHgsYYK+bph7amIr
aWFkltHAApWIr03qlaBB6tHJ3OyJl0aVy3+l9QtJRS2BeB+H+WeOC7UJng0N7WaxQ8VSWlIg4Y1Q
fwdHVWvaLDhKZklzhuPQFslHURai1jyLMd2f432wRSJWojePNCTEHxEWly7iOlSEt+kBw0BV3RTi
wMSTYay7Y8+6k/iNzdZZ3ZKehxaKbA1UibjAVr5vrZkdvp/rBGjFdmYA6c2EuDocKO/UCA5lx/rZ
R7cX3MJdJRHCzvaSknx7aI8xZmLlM0T1M/7NSKxz/huhrf9b6YbkEYFX2lKGvQTHcG8HCoZGcaHP
r/4dInURHTGgzcOpgwM+2E/y/G63hTXK92ExBMm+B9zjfr8f6OqYAdBglH8AmYOUvpfSkuk4huqo
ZY/Jtj5jKsRWFHqGMSu46GBppiD072y1xLsdySKYb2yehD1uTSF+cXwlCZLKJti1dncNanBE5PsD
f4Ej0+QbPvtc9tppvcZfq7cjQLBW3bjDdZc+vR9FejPt0rG/dkNckn0Iaos3uj62QEZPX6Rgng7P
LhhQzzmScc80Az+tayT2lqeXQNez47Guoxy3aIZn/mkO7GOC1EoELYtLYDnoyC1NzQU7JmTggG89
tZ7bT0BFyhR8g/egE+5+V8a2nz2LJgI69o+njzKat3us0/TPT9p/crCGqckejPs3HIA7+AlXh3fc
0q7qxMB8LTJHn9Lp/fKfO5VdDivF5wsdWrc+GnuWBGUdhPs+fxP1VoxZCnLBYOTtG/O65tmQojar
3tQJBjYY4tF6TwPmruXXeBU3PM4wGYcWGtF1XVukFb19xouS4Y1zELUGQNZGT+T4pRPvUEPqz6fI
6YzTTtYUZVnstCKCylcuSBbqSnBAo0/4GBD11y3FZSBvS7YQRh0Y6Qipusqu+0LN4rECcxOUiS+l
pXyoo7+hiwjGKRllAQ8rz59gUZ+sLp9BSGh5J37aITn8Oo2SK8XkYsXXhx9Eg9hTV7/xJGsPAhIW
dlBHCiEzWze2f1ANKU8SJLiemmzhXx0RTDPq2MWn5RGYsbJqo8Ajbbo2VZbGnhBDo3OQsTCQ3fgz
u8DyILJ+ObWSgLacD1W94ub7BA4p72Pj2GL+bXKfQ9rc+SkQ2MGMox9hwG3Wuyz2nOkEpWRd67br
4T2IuEWK407dEkH9/fbNqFmSzgnTIxVv10E6fBMSaniFlWX4gCVrZKV85cimOdmT0HmFywwY92Vd
6NSCTvUhwsHVR749vzllPT9DAuwVhUAe3XUlr9FcywONIwmZLRkVwJs3kWG0q6ZF8CkZwxZ3YpKf
cUJHCbFyIqfPAzZL65iEgNpH//FJ4rTaPUwuo1OLKX4IBOm2pHL0ltyYO4Z9RETqbrPgugfjxoZq
67ghqSwV/iAv6hD84URwSFUZ/N2Uedy/wLco/WFOkXbP8a18QQ710M97gvvxrAkRYTWX43d50d0c
BgerbwRLk10vmF68/6aGcmcvnbwtkkJ4RDyBES09ggT6Euqwa8o7ZOFs2mBfNw5rGTI6zr7DNmp8
vHpU3ZeInK8JxHbn2NFWdWOiyfTqhxczzkyox5iusndIGm4BwUMcwRs+XO7D4ST7FGTg32TO/WcN
N5dO2yf19Krd3WLyE+iOnHPXwVaF9QUUWh8wcnsFvYZb6omDruZlGYpNJvKYwVMvNkDIV8DFx452
LCbikF5Sfnzp6D1YlkRIiNiO90rUOMEPaeW9rOYU0iITne576nl9XTeDXpeGaKpZPW8uMDmNLNwV
hC7ZACFDptdZE63SLwx5gSTuAU3Ku0PMNHB0zlLUqO2usODPuzARL1GI9NKz4wWP9bMctMlbNc3U
/0MKrOhyOcRUiEBd+1Vn29OMVGdVNri9/PjgqUFXJVS9nUyjm8Z+VXaASSmUFd3MdTih6eL3b/yZ
xYVQSkOs9WI2DL9YB8YombZoDoeKflsJ2MXrfFczSN8b8tRUX87mvRzKtSPKfCXccy9peNLm8lqp
ofkPM+R7pI2kVUX/7iSmNueJiNhsSqEP2FTKyDwdq93MM9gjgXnvDFFuhY5Sx1951+Tg+sAGJOon
HGbKOEb+DqHmuFcYrYsIuo8v+sa5jUTwVrKpK7zaiaJQXOHHHgZSXaucer0CW0mWCIMz7InB5qYb
7aJ3nlwv44Zi/Q9o+3ujQdlA2ltVSeX0BsfDCuTG1+u2APx3cbvBOeg//OtZXjQfBDIA/inR0o4T
tzs2v+EZ2JJxeifnPIE1GjslgTjuemLFMXJYtNXuuvjwyTdSP8D6jqV3QPpDxDPgiGpyY+5FvlH0
kmmmHaIj/k1vNDOZXYus9ig3nze6OD8RiBqceZq4akAppNvui0np1+f/6CErhHp5W7Mtl6B/Wiea
VJjyzz0M57/9ESsMTWUYsuIWZKDvKTQW7LZDevNT5g5TLPPBpPxv/Pm8n80SFfGP9EKxB83GusaF
fAtBdvD/1I4/IOh9ZqXcn96w8gCkliY1f1eknpmv6ehPC+UqrVGKWjCHw8kriMnPSR/8Z5ttKnyJ
3ZvEePAX/Vxi0ZVzMrxN4xcuwWdAeKXCt9jc663yMMd7osPBIvRfJ2HTK1aTLh+qzpth4DicndD1
F5qKHWraPxQX6em/T8Cj+Qul7G3dOwIg2hcPnV/9BfkyQZkGPUPh6C9B4ZY8W/lob5VR4l2EE24p
Gzlu5yvxQ0hp+4Y7iu8ZuJEVIvAMLPLwVfhEho0VV2cWXoTsZXUkTT1WbfYMrP2ZcKRtk5KDB6yg
sSWtXbEXkUWzfeJYQ1veacPAfmBMMo5HTF1j5spVDNbswaAYVCIx3dg7HsCdYKovyyfHtYxFGI5P
ZjgiXwWaqRckljbSeRr6kci9Difgit8wR+xW0sWsziILFmKUifaXO4ret0iJjbyTzHaKHdD7RBVL
AnVxj8CXXB79NUDcAcgsJRzJNvhthZbIBpA6Fihtm2i7ldrpA41pBk4WQXMr1HdMb4bo1qmj/vgO
p6kj3VWIQzpHwra57/2VBKo4U/wNfkh1yysxh/S4NydE8Ic4w/Blz6IVK+fCLoDO3SfO+vMsLxRp
LsdHCTkkTatjwVKtAbCiTc8haeQoSizfyvVdGsBv72N4DHbh6Upr340NfVhZA6rmSFE4zgSSYVX8
vl4CTQTdbMMzNseSiE3ag8+FeR2T+U64ddYNy2h8kqPiMLuIQjzedKnaCYx3DdFoVNvmq5k9/dZM
xGtjmiSPTcg6Km7E3/KY03/7TXxaXeM2CmjiehxaalgkomMFJXOajcaDk/IoDRYECOy6gtRrw5CR
81Ki4NFIzhnBaSzBO+349RFB8Yz3Gjt6HeK5infnVrAyK3BNUABg64cXLSqCjTBWVz6ZDGQfM1R5
EZiI/WmALLCbkTbrahwt3/KrbLU/Tbb6b2ZwNo8hx3OMQh5eCQLaBu3NHVxvL8Dmqbq7buhhSbAz
Sd5C5u/I9nhvkOWC07iQF9/CVwRwZcfLsSQlPHnPO7hKn+Ug3hYwqKeNgM8jk2YLnLMJ7j6CPUWq
oR8RtQaGfkQ/CLvPmjr4Du1PLObIoB9ZClzZLj1SCUCr0nZbPm37UYu/pIW4+aQaHRCjexi65fhF
B3IPl2luUTd3VoUai7v19eNSYYXiqSbHMriWVPBjubw4s5HWzs1QiQLrd8uErku8qWCcqQXl5w6j
iQTyorhjOgVHClVtO3yTciw9Uxlax+hOWlIgN8ehmQRdyMmCVkXOwrXg2ff5Rxwpd8iiHc3eDXp9
XYM6xzFxeNZxh8GcNCQfmSAyBhoaPK6L9WqkLV8elBVbUr8Sk/XfzZB7Jvet0ostIsKMgmNc3MeI
Olu18v7tL0rz8qgDdldn3OZM8/NybsVF8/D8rh69BatGb9B6PXQ16OvEJzp3kSVFY5MSeiid6doB
nEOu8tehqqAzWayQYGBayEqDPePgRO48pPLBh5ODnjLMYenneH9SvJM9QPWLWw7q2iM79Gvc0xQX
e6+xL8AP6Szq5NVH83gaQZwdXP4fHVhPuHgub8ic39TJKKChi2Pp+XaNvOrLlM768O+LNhh+F74o
GhfWpOMKePQo3ALqRndF4Zmmaj3rBOINlTggVhsiV9axKS5QctJTHsp8CO5wgmEQHCteRizu/ZYQ
a9nl5iWv6Vz3Qthfthw9Cfnj0na+qLSkJkvc2LdHDdnSQ7M9eC4Xz56UhJdOZ3lHdl3fEY6YRBXf
eCAF+PTnl+lu0l2cmRgv9Wo82Z97rV106N1b+9iSxVCF0+N2eu0lmCaBWEvpz+HskLNO51IbNviy
zH7xq/aPiq6HIjt5w4vk95PAJLR0KqBLTS/3MYlPsnFZWQW2FWbZBtQNUcFZxGFuLJ/daIh+8kpE
l47hiTqAZMqtmHsqNw6vExEPkEkk/i7mjnA7F7TziVvH5X1ujFFUcw/TaERihpcBtw3AVmejS+dT
ouyBWnWeGILTuOemBx3fTuUfR2lH/DWz3snuQbNVqBF9ypV6rIgNA/ujRX6QU67DEHt10NbYuD4R
sg7MDELhzjnRRL/TjPudVlQ0D+RoY6GqIBozoes3QuAWdWOFAZSiRwPlRhviOGFCpE8khtZr4CRb
iKC75qc+oTmKOkiTC+sViNd1v8T3b8CWvqpLrIkmWIY0Z3ttXAG4esGkktIcivp+aHZdThTgjzE5
S8qeb0qj7BKIsv2rq/0FMNMB2GSauwjy1K6zlAZe8KPzE7oTwKX3XCBCJckKXrcgSIOexFKlA/Vq
2M4/k3X6++pkfZ25cAUT3v9ucRCZ7eW7WkJL/IZSe6iAYlJQnv9e0Zg/CvXat4FtjAHH1jf7ntzs
ZM8VXZNIOScVQrke1EuVUGi3ICBfX6ObyHawSfB1I2udLWd4Hb7DaAwiKSB+SkVQj4GMnZvYp9Iz
kTtOtHN0Pzy/yyoHWou9F2dAdr1uS4G8vW8NhA3v64xEpQoXE8sBOJnG3Wr+hjJHSmOSeh6SJHK1
YWb0/j/osCfBz/EFh7+VDk2fQ5inwUFu4krC6ho9EBoE4o1OlVimAd59jwQrb8OOabOKG4fRXHK1
B2E1sKDEY+qssYwR6Z2JYjulE8tSp4jcuiI38kSiEUk/bxGIKS1/WBvRvzhZuscsgce6bAYtkbT4
hGowm2kvQWKYbNGmcuOAddAvcEMEF9vV9Xwv/0Tpgw724r6Z8DZWbWiB45GJWnDS+fV6bw7LKAuU
kYN7Sg/bBbSqwUTiBXX2XBHM2od1HHDxvCUb7gLj4mpP/byrKr3IztIEzlJDYjBxVWlOrOdQguNT
gyqlCvbWPl1YmeRG4UTJdMn9kOL1qHAhuJlZ4V54BtlrvAi6MCIinB5PPXAsUKrDm93dGK9ZLBu/
DPtnK9Nv7OWpStkqYLhD7GXR5CuJ74FUcrlqaC8XgujImzgonb4QEwT9KK8Hb/DO1rP+GfiGzj3Q
O0TwpACPIRgNCjovfWsDHZCNIy40TGsMRSa6ABlyNimdga30A2RoCcDOHOrnTPWUObmnP4BuV6I8
C86yIPIoaVd3/oOgjP330iqHDhuKxo/NwZfISFYD1rxUZp6otF0MVy7LWb98bzCtydxJhm795HMI
60TFdDwQsJYZY391iEVWC5Hnl5QDv9oOclQXgcck9l4ARYKNAA9+jCHqmmyPpRQLr4bokqrAPhEW
iKUvT8NGP2XmiC4g3Z26m+qfzwfp2IRHKvqvvYZh1k7kNcfXeFhQn/9cencTSzsxlFAGoO4oRx8J
DySt0k2wjTb0zcNLOLAkdGKTYMpEeH/I2FEFnEZlRG+JKgxc9a4LEwZ3nmhLHQC76uXvX1ZUTiP/
vO5V7vSz2osMo2+zw6vTDGaHesCL5o/NWpMmzjkZpuzjH8O/qD/y13bzByW6j7CzPGT4BSjclqlE
JKBrWn8o4U2rTFQjKWTPgi7i1Kn7iGR/aV4um7EDNb3vOpvrgeXWuo97c8b+X/8pfYoqwUGeM2WC
4nEyAJ2HzsHhX2GpcRJbr9/+QSlHXDgKc2/cBJzpb6m9oq1tu05se5hC2FZ6cMMq3Z6Vq1gqOn3i
S8QCISZPs3XRY6D7jmuF7xT2UqBz3OAstwo6yZBvB+F2GXre7ejUml56FHp4Fj5aykjIjIQtjXwe
mgG1zFMayGIoxo67ewBrFGNcK9CXiYsHV+lQEkKvfhrNmThX8nG4/D7aJBr0vEh2OaxM6PNB2kFv
kKsqs92bfMceNrEWfP10yWP7u4fDdYwOu69VJI8F7vXX7CVMDSFjhaTbzc3bBr5zmanoJmaVJEDO
G+nzYfN5/f9q/pvAgXqMVeLADT5t83zS3ZbxrLth3bsCRleAVofKYdfO/Hirl1Lt74UMXhb4TnsI
ttmr08fO/q0dDOzBhC+jt2xe4pIOLmmmREqF50BIkKQ6f/j8ligzy+nuTz7Ut6d8lmLUMqS/bo3R
2vQJhf4yUQP5nn0PtKAJVjkg671PRJFRHe4pZyfeyQhuiIyvZ7+SdVPtX6/10pCAxVy+90fGdAjC
yG8idBKQfkpgDWVtFzlMLxumwrnTyv4gtsFZq3fBeW/ZKacvWrOMMivBuJsnGX1btB3LoWKizm36
PQPWkJgx3+hC51rSBR0WPufaod0Tva4dHpUvXzR+WXGS3bLiNMO29lRsIhQ37BFKvUcKeyoDvtI3
digYvP2Qqig+CBVXJa2I00oVwF10W3652NkCqcJO5Si53zqxKOnScbZgYmo/Ik5MocQf7LoeFjrk
tEjwihlfiBXiKj2psj9/FdWAYxkDOJN/r9p7+c1/So3+TCSyt/Z88sKlp9kM6ZOYRD9DTHykd4OQ
oe3A49ZlIbP9LYc42Y7L+tWLWVqIOTZ0LzEvXui2JZv+Br75CJRburIKFhhCbW/r03F/RAFjf4nJ
C446nSEaz8LVE3kwdGsruIPuuhgHqH9X0GmOSCzv8yU++jVgPcsDsYn1td/yFiL8iQ1sJuwMeVOG
FNqKVo+wPKT1C/lok2fwSifNRfrOKA91IVgdyJN23te8a7w3rJokNWTYMCrGU1ovX074yE6pI8Nv
PCbL48tirPm3q+NkjNl20vnBgRlAB7+BolY29FWvaNbbj39xvFBocy4zvEleO36ZUsQTpOU3rOxQ
pF07jGd42BzaRmpirmD+1BBlM0w7Ke59wPEvSXbmgWGXLz+iAgj6yI/eUB0o5DF93p0nVlyApChx
oXsnh61jmouAQvBxh43cu5hVbSjxClMo5EmZ9P4WWV7tkzeGgkLKjZiUDcDt2G8NjF0su75oSHE3
KKXMrtBS8lUS8cwbkUKLjJ03+cZlqbQLtE41A870VJlNKw+lQ/H8U2Mwy21/w9rXVjTSWFp5RXSR
uhfvEQ16MFrkb6i63BvS6RcrMrRZ1xL9OpLscL3Kdv54/p93Rb43c/0wYM1wrdv/ShYlboGXgEKY
d+CxW3oyJfZsOSk5Q7lV2FgIC0f8hZwJcNrOaFrnhA3hsBbAKam8av1WXLjhOPycUa0s2Lsc7+JB
ACNyVoGhpKtshDm6fgphnkr4l3a8MYANP9ccI7EvTV4FPMn/wQydGvleAw8XNe4bNv6a/5s/splS
2kHUqB6HpEn5lm6Tccr+WFfEsCFFXSkdIok6qjTUck01mSW6qdgwTmWF8C9fTGmQdYPPklHNDpxC
Pxk5A1KTIp4DVTw9uX8VkCvoBuFDJPBnhaV05QBM+owEldHNK1CDDKD/hfdvipreVv2ETP3EEzEh
WvlltxyG5Mjbq3aonNd2URM8mo/viOTun1q9MaJsUhsgSj3JKe706XcP/oI2UZ/OteAoINIgE15B
4IDyBw+MFrjz3fg8nSbV0aUHbdyRLbc802EDIDDvi2szUwoXtH7XU5scjd5keAeHaK0jh2hrjMzy
o3eminUkAiQzKEUumFLYgU2m9kdh7pwvL/igXud1L3V9RWfVXPeLjhXoTPaN5vGW6BDskF/fOvZ/
Q+XP8PJQfGywC5WwVfp3kNvmr8ueVzuv7hvUWhgpyo96TEdC3ptC78yFEYODFt9b66BxZBWpzkSg
WvlePKhL1z2k5jcJTmIqVZBo8KUnF5+r1TI/LMV9oi++HdCu4lPF+ztvilqex1kg9tZJZaKfW86a
f8VNxGhOwiezL7mVsua4Fv9uw6U+dANTg5Get4l7DYUGOK+OhcUQeukDVEtYdB+mCO2DIGmMg/Pi
2/9cLsvqrd1gyTcLqPYEiAPAJyjbwuztoRhcwAsW1Xfhqsfb4R0hK5AT3bqcl99/ZeZRar2QXOEM
4p1CO1CDNQTdOtXUqRb9w7I1cvAJ/SR8K/7NEUdH08ApV2mB2vFmTleG0R2Bl0uaGJRoKyKTd0B/
uV60FXwfcojU/fwoYQswmOTzyMyIOsBHFBAiw2xxeRItfKJcoaxFAnsfjeFGr7vsODgk1Ns2O/WQ
oPoiY3kmz/+DQZKX9JLNr4kNDvSbgbEVjt9r04dmvFL9L5kP+u+4OPfBgyyuheHu70IpuwKB9RIH
IFTcye1d592xL3szsqsIGHWCjt0dyqo4/3d9mwQumQafDmgc/r6uq8bDdSCVylPxls18qBu/UO3g
LkaMJL+x5TUI85VAKg5+25VAyGqWjtsV3wrbTKS+jlEO01aCCfugozWtiDYYQyENH6Ns5O0dGWKN
LCACCx7d7OBiPjKTmGqonpqM5Nr3a3v0kVmM+hDXdERfbtIVLnGHbfNzkzBxDgM8HtwiHnXcSIC8
Lvhr87E+UU9IITzdfJ8GI1fm+fhJ5Hj+o8BjFpyDKcyd7yT529R8NybL4NVlVZHevXeaGIUaVSyk
Pj4FF5PAx6RYj+HCyOuiYu4JdZMFQZr0uGZCKT79hWdZGM19LxpLzma5VDjBcey8GLwnanARs+dD
3bhO5YJK+z6ZaMgDAoR6PFDMV2TjHBbqSW+CUJd2v1Eh52OiMGsvexT8HIAY6sGFFVXBXFesZtbn
4Mnto2nPu3F1Mq28LfGH0y/RWpW/2/teJdLe1N24PXO8wFtqZC4S18hKo+anDypqHFeBb5w/iylO
L5KI7OfabH3u37avafiL826sFT2kOQRW4xrXvAWuUYOXd4AFA2iFaOdxMjiHEisAN9LWCO2HY8Uk
SRoLD85kW5MjdcTFIyP6Zc7XOIqnL9iWyWWTj52PxKfYMWMXhIHakV/grMhwWRFYrpvUqN4ya7/R
68ebCmvdMVeDaS5pxFvKT+fgWX3uhHsF2qMv+inkuxhUn4BlXQkr7eA7TSGX1agZ0j+px0pkjsfM
dcpD2GAUvxyjiC7s4dVTR82Os76F62bwoLu5Nsmp8uAdcIaB8vwZApq25I5F6ATyjgwq2aZCj4HH
S2UOTLf4phbSJ/2gdNdLVssXcMLxd3TZcT8qWA55W6QQza+t12P0Rv4WMc0gBVFS5E6qtfOXYkaV
JwtP/I4pUJKaLjn6/DOVjXqerySgM9pL9T5a+5hScA3Oa+FhmQfgZshZA803k08sTYrDsp110z6p
oSAshcLXUaEQuFaQcF3Ej0X0f5tS8m3davDp5R375OddlWoD02t083B4fLclS7tt1Tp5Gi8aUpts
Rwyu389vsJ8wkAneaB/deoY/hRboVg0a1Jb7dzJcmlc2oYN+HrfKvCHpxdvGU9unLR+OZVVNc9o5
Z2yo/0K/TW/lUrSIDJVWAtN5m2Tt18Vooe6UKsi7uFmLB1/lF58vaJ/5PCReRTTbSjHcL1vIshNG
nLBwx3uw0rYI0od8tqvre4CjvWbE1CT97EEFwQEkD6kkcMwZPClvSr3FxJZAs0dwYDCpKOg7ssyB
F9R13UjqxzGRgXbh2yUPwHSIT/Q4QRJZMMtOuRZ5jHm6y+8Vi9SmSdGvzsoTdUgKY6lReeYo/plM
CQ971ES9NSemXQ3B8pB/XAGMkk8o8+ito4I9jgbGVOW4i8Esb42lw9fMwSiEcOvTrPOezU2Ps83l
Ldwo9x6Vdc/xTa37z8QELeT1McUpS/YNuAI4JD4VJjDmDiWxpkqbKI6hphn7dfVG+W5jTgsJDsdr
xtvSZR2kq2l37hWz2r7YSK4y7anfzh/6i7fgvrdeqX6RfmhAoJm86slZmXkyq2AzH8wx3vyZ5mqG
TS9HrpQH+ykYNjM/+1dqAVFO6LRP8VkeU9vm5hO5co6XBXoZs2QjKk1Uaanmfyh2EW1UoZbtAMkI
TVtc6VcuiJyuFX2aMJqQN/5YL6VvSC8Or3ntOjpf/pApO8seI5B5YVi6S3ofC1IJoY0qBjAbgetS
6BxdmSATV9gwaXc7nsNL143R0vMJgAT0IssIfJaJRHPR+c6GtaSMS3sTrmS2aUCWKaYGmZzloD5C
bczlGPxrzwWL+BdO6pMyG7PA5hmMGHPpATPVivPbOtrb1IFbgvtCqh8+Ybp/iWcaMQXv/OmPxQd0
+wWI45xIvVK7tThjcfvt5kDdvfc2/7Sq4ok49R71s/MyvTVqMajzszITpUI15jhm+7o6QqcZsPeZ
UJmYKAfjAfmsE7coGomgJ5c+eVkYh+lN0z08hA/R84CkKDauGdfRUVJtBC5y9ktybvY6j90KZw6R
GYcYSxyJWxRJTO3J0mIflRa7RAY34JcppNGDFCkZZ/baj4GvGYNi2zMXH4NE1Gl5tZ+WnSUY+DQj
z1+LJm01yNiMNO8jb2tO6+xerap5VZTme2z8+X5OyE35XYZd6ZbN+IgOf+pWwBchWxNWoRTy0dO6
cmu2fpEp4nH4bPDNYvqMKHAl0HDy8DD4JpEFIYAhYQxdewzrAHzwWCb2+oK24c8UalqmVckNr53O
ljpU4mWfvl8hoUKiQSd9wS8z1EwQeYSdffanxuf9KvPYuX4ptDlIJxx2cU+tgQ0sNUmrOdwfSvpF
IJYqnqbhozkHjFBDZQr6pLGtMJKom4pk77qtf4ToZEX7ZNAO5pYTOLOwR49cqHEnHwCkDNsU/noi
mGT8iQU9SjlpKRHVu1O/mN6PbY7DM7roZ3dAF/ykUB7G2tGUmNg/YbA45HUNTA4C4i6XRLtoZXsK
xkxjQvlMzBB+h/B5Mu378MBMcWBIkTNpKN4n0agV3NAN+aUU3kJqW61OqgX1JtjKd+rhX3iVUjtN
xBRTP4Je/mkzNEJTC60OIOb+PqkpG2+cqWAC0D+SwjwCksZ8drBKbub3kKQBQQDHmHgd0vbTSoPd
HlVeSILxf/ZMQzyDQGUG6g+9+xh5oywKQcjo3p6uTQbIR3c+3m/1hvjoFqhy84wFfeoA/nsjLIMp
2eb68Bql31C9Sm+t9+ug3PtCkmdrGkFeTllLe16Hbk7GClpncAnTE7EUusmYkvgnEyNHuJXDPr8R
LEX+iqpB/DHFZi+UaotCH7HHwqPByHwxiXV3sseMBwSS1s0RRieAeV1SHqXwU4lqNYEy1B+iuwdb
sTqme3qYNQ+Oy0BQ5dQpmxCS9EOoXbstElEc4kOQDMReWCQj/zyRvhZo146WaCTg8UceSgoJbQiV
ES/K5CMbHhrXQ8ItQqVmV/fDQOZzuyTgw07yTebiR8RE4VR4AbRtfNUqrVid/4ry6XoSMqrnOLQH
IJklRWAq71nPFiiLPhcm5vALtNIl86AHsJ8JdeCpHvlK2bw0kvpE3gDeVXty4RibzyPxKIUhd0qj
iy185kkIIRxJmghFznvU/9s9QOAym13wbkYd4CVULn0OlQGrbvn6468oFbBpA8zsy1lBPRQ2rh93
cIt/JO9X5ipNGGaTrkqX38i7icdF5wa5ilFz7Twmo/AK3Pn1mOuH4dRZbHSLoGNQ3GbRT4/RGaFZ
3LxiCm2gHG3cqC+WjRLsy1dLZJfD3LKv7mLAiydwIvq9Che19GU8STKnlcrIJahLMKkgDnfTcg2L
dafADBYsELtYxD9pOMaNGNBIzcyfxmRToN8TBEofpVuJyja6FTD6aUM7gP53ecMTjzcJZyJGiumF
InBTVIBOPsABP/obvQ8osRExCjv6hIdVnGGZtnVIK+rgAgHUh6Xk4kO5eyKmLF3jXF2t0Yvxe/6d
HOjCKesGwy+DG7Vw2Mh7FHzGmqcxbddiwmM6+tSdPPn9Rq3pJEzyqzqREJr8myDA/H9w1KQTv9eb
Zp+XesrXQvx4uUIfyS2JxrQplPeyPeY84U7oN7QYM4Xpl0eY4tw9s/MAbtbPL0ChNUMCrqMYBV5x
mdDtV+zAFHl3OuTGYbXHyhCseiZXtr97ApibUz4dw5DKBboEMP9xOhBfLxTMA0BkqEygiY/ha/hZ
eoxNGbNWTiTFvumMBEJMiy/FIYJpA/M0gbNUBtxXMiP71XgFRyajpVyinusuWgKztY0zP/xVRjIt
POLo+7cZscQsxVm9tP+AwtyA6ULe0xQLOMkUPnKSFnOlKdpoaAqYRvjNaftfKURn9gfWHRtHUdz9
i8iUcVCpNOmvhbdDqRGOljpGFO0BfHXSM5+krhH8qrnDydLzJJMR4uBDzn6JMvZE+5llP/19BRcH
YgP0NRjSeebkOmqp93BsTolcWtWbmXT6EK8bRU286HijAG4/tElkDxydAmTawatCEXvzUqMS5jYT
LjaCLY/9CwZ3rN6MyjbihbSjTYaseRKYy8mFKORqwiY9RIsi/rBRwaVsdXwdc4PwsXTzNiC7ZEez
oVT/mnvr35GKQUJ6+JnRvETnTeU0FhMBduMWGoi0Tu2qig/ztOM/d9HsJyT9idj9q3sy7ReYxrZm
zEjQyMdBUKDAmI9GqSxrnoGQ1pBNnf2+Y106F3bdU/bgPV/GBmxpCA2xuYpavhzIypvGEBUiVkxt
q8K8i9lNsXqQ2O+rQO6bntN14k4w7cAAgLHe9n9cZiFb8vsqXUm1ydlz3QKwEmgDMfOvFlfC5BGy
S9Ic3XVRDiU8+ze1yJLotnSfBtBqV26ncq1xUg+bZlBCI7qHvGn8V+GawIGPKELSbLP4xlmhD54h
QwITIDUX6KrCjOwReq0M3NB8KITk1h+gyAHhC3UD5MZx9wzw4j4tA8g8E0NssE6H3tMdt9uRoBqg
qpWYDPh+akKFbayJCb0HBuqOjyhEZO8OBxaaoHb5JlPgzoBCG/1AE4ZcOxBpucnpHqoVXcYmOfHC
zinHbsWr6uNpYpQ0LGpyJ7ziu7zYS0UCVEWQdCNYPpoliJfZ+CjH+mck85qDnIQ7JuYA0GCIwESI
vuvsx2w5+/l4EfG6Vxp6S5LmQngI9h2BUHVSDsuo44r402SJSnU8rmGJ9Voi+UXvVp7FXL25tDUG
qfmnRH+hq/9kAns6hDSHcSZKZnQfcHdrnJOK2yjclaJU0E8gIvDauIQnuiAKnkADj2cGfLXLsrAu
6V6IdoiWvgtATIHbGS3LnnPn2QmaQlwV1QNBpmLnQkpXjIyazBUpNy8JK+adK3hzjMUeSsf2tWCH
m3EKjE5yPF3jZK/nPVKX5uqKTrvIAJ+tGKwyc+PPCYybyEtwVpPq2r0buhOOrtkbEr6fgd8zDu+f
94PBs9xFmK69wNfH46YjopaHxVr4JpW4eyUiaFyjgzoQb5VGWJQBO/sv+hpMbb4NUUQbSa+SgE1n
8nk7qEBh1sg0CMFHdlcHmg+4e4XMDqkW5aTu1w7dW3urmhP4jJK02PzDhNBzCu+P+Hc6uzZrFZ9Z
Kmg3CHKrG5b/cpgR15SHxw/h6VmHCkH4bvbYPEfjwhv8LAP0YjSMrMDvaUbFuzCZsSG6WB9lUlIs
uNoytX/qkv//44dfSWlCrkyGPuTo+YLH9iAD7lVnB5A5OcHQu4IinufoRjOSP6bYVcyrfPauLR9a
b6dlCacnNKgfXH2ScbVn2C3foHq2pKlPXzj2sl+sHIwZBsP4kaqlJ+a0X9iPsO0+Xirg1zqMGlPg
y839XoRl+/RZwZp9GU/NDYNY6x9BLsCwP2czrR4PjatfLBaxTecTcMvxeSBTV/HVxYgWAdJYddlL
25fXUV0KR+1wWFyM3/vw5cpPMdebhRO8UpLh+ZbIBLlXmgTHO9GHvvtPreujfFX+yvFKi3V2bZqM
bEvJ4a07AVQ04jxFDli1KHmSbutBcBXkCvM375vO3w1WjHJTm+8EchuDyaWk1iBIr6I0W5czkvr2
f4EtxK2guGmTipYCLPJ0tdVMLr8oysQEvTYEN7k0+tgVcO5J8fuqUV56Fj4bO3ekdofz1AD5I1AE
kz+NszMTDF5U6watYb2Ce3HCqej3frngx+XiUH8cEUCDAOWM2cF0FCXDifRfjpwxyC5q6dvIMzUp
Ua5BALmn/gLKIGub3EeXSSSMUSNBs2XuJBriOA8SapfT2qsnqL4feE+K86oS/LqhsDJZV0ZFbV9U
jTwR2YA2779EKtMJuNfUomlpmzRjst6eEURTkk80p+LT+4+RVgBnnLfCwa6SEJHIEqf42GYqmpnG
E1UZVmnwMiY2GQYCGPgbxuLtV3e8ICBDOzEP3eeoUnkK3XBTGgVYSRuO7Kymk4rwubsPY9ED/rZc
x/iS/ngn6b37JzEQNAWeZh21XX7ahfAd/Cz6gWYWegW+D2Cynp58m6JiFWEE48dnunhQcgtrbCxt
AGsWYZ5vCbeUq+lZ2iHHryB3ZEUUNAid6jDJs8hTIvJALOO+aKzYvujVSvpWFBm3bDAGfdkyJK9a
Og7m2/GCb3IMrxtz1xXHjU5cj9hP02t7XpmtMi8+eMGVrw5tOQxQpt1E78MpTqP8EEPuoanFZ3uT
5A+EfuXd37kZpoaqa1xLnU9jYRJVPwdVEiOpUB9QKFzuvRexl0j5BVal+6iYr+/mYO4oMGFYR706
/tU9qDyREDHRnQi5s6OP+67KJbIk7NkPfQed3dAebbUImn/+pBLIll6bVO64+AWJeIPMPNLyJjUC
sA10qbYkpNF9BsJ1jag0dtxKfiqdcuz7+lzS3GXEF5RjO2JBazvfEs5W+VEQBm03vt64GpLxIclN
ndHKqitN6BL4MLtJWrvZiP/lDi3TYJcHcfiuAyyj7w/TXnC1f6NjIKZRoJU3vJ7fgxO4pQ2a3ngg
xh8heOM3J38fmQfFcpL/cLHHsy1p1M+WcN1ZUNxDdBYt0hXwwjfibHNqSlOSM4HgMgnZvOilgRZq
nnmDFqvy35NnMCNUZkPjjW80aEkJuQbiRq9ctCyIHUgBrMxQ5q4lFs0odWLkDV6CgQ8l0oi3fy+n
hLeIVlo359HvMzLiiQ6R2h4oAvLfOYEtI3a4f5+VYbsY14dCUm8/LVtvnxiFxpVQ9HqBggc/qXwb
IvBRqZxs//Vg41lsD8yAcKR2+PDzEt6ng6kokj36nsE96ryz806lVGPaPr5/EDs9nLTTgoja/Opo
RVreL+/7B1YBhSwXCggUzT8hKjEMOAjfk5sq0mHPlwlAmmAe25Ji1dzSn6DrH12lBeZnY1IRnBDk
71AsgxkQg3IkBHQVPmw6Zma8f71D48m+rHYObfYgsFiiSTLlUYYJEXiuL+jGmXJBnsrFxjxTodVY
NwQC7faLLu7S4q2rG3QbNr7dG0WFUPzIMBQkafxBJvyIiMRop852h7MdxLT9h4waVjnZYpVtqGtt
ZUALCtPxGbyXMK2wtQfLE15F+qr4lFoLm8ch0umiGzajHBYNX2r7wRpraop7HdnLwWOUWrolCrxG
dYC9ltlZ6hLLs4XTkbG42IxX20nK1D50lkrWUXK7WjNoGBJ2gANfKzbP85nNXfDBcSyhZWDpKqQD
MBINjkbz8camscHWG9saARPaSymA1OlMshK8Y3AuPgELkuuPVp9W07++6YLTUl2fLuwMlWd/kQ2V
HIrxpZQHfeapPAQ3ykc5sE7NnW+cCWunBayLEHdSctGcOvm7TWgP7yExzUABGrx8Zd1cB3j8kckx
IdE2sY979XbAAgm1yklH4/UQm0+43BsFcbI2FTwm1BqmKbzuPg0RiXHL5N9qO7uQMXZntGNKHhKU
VsYMHXgp0O41V3JIdI783JZ/DRSIK7heAw83uWbLxBVXoEPxsmIOYjxK3HcNidAOVNJhbCuiSSUm
ByA5NSuMzCmC6z5hf2HtI24Oao8v2IB+iczY29w6um37I+jj4ABcYhLrLdDT0yaFyTdm4UTI3HYe
gak/LUvdIsRui2zcB7VjzSqWCly3yrutA2bMR5wkX4Awu6MSJoj6yXlG1mlW8Cc62ZX6if8an06k
d6Hi6Bg962W6oWyyfNkm0HqY/YevPLVY2XvUuJGqx9ydQ4V8sHLBEBWr7CcW8qgrjw7o9OAqQO1r
MZ8HjfX3XRebq3Q8qm23l/IfM+BzjOAoXVLltdx5XiJ8A6evin7FNd9qgxOSMpBcniKoiv2gw1pd
eyy4zYs9Sh00YkNGvak4pvOxdJu+GOlYJmzRiF8nQhXifbgCA8YqzNfF6iLzigoRfu4F5xihQi9O
BGu0CC/r/LkuKwM4KJyHQRm2XdBVC3EPJ05/MM5aMPYx6SWojktcZMlvaWuGObbSyW61xHvMw6P9
gj3Kyv0nSGWUUcd3ApIcqHn4zBlyEcX0V0t+MLRvNZmPsz4+sIWLqKmxqpC+zu7HvzcwLrc9jJSI
dht8LeMDTMM/FF8wNefqJwdSdDAg5P4TLZyN5Eu9yDM5MQ4nZw8+MGllsJybXK/ow8hJ44rsINSn
zeRA2UEDDk7XJfnc+V3qeN8SyR0GIP+KdC7iNiV0FtPpZKYJtyMB3UzXumqpFZRBzs/6KCsqXWn/
sAtK/7E2nCoA7DGHL1wSsPYa0jcRnbEpIv2rXoIzq9FMMrK3PjHqzjgDfp6fyTjUy7zk84L3Tfcv
agNgbitg85SjuluTg285urAuELXvmd8wZnVwtTOtOnsmbRen3piJ4B4QtaMELj+wfyCyjG0DLIxL
jKzw/C8kxqI1uFq2NhkV9cLDwxqPCvMsR8OrBQDA5dUI3CLldMi+N+S778oFVAqwTgCjT/n+Pm+x
46xObkpz4fAMS4gfIQ1YEhszzEMjaNfieA8eUp6CgAAq+QZTwS3oKzu2ZoTjRX52Iy9bUuFBXCkh
D6o8pgOawAfefdnQKqxjm6DU8vNT3iMNQG3BHJaiQLfv0vsWHUqmbGNu3+KthPmjYhnQomCA/k4x
KsnvCIPQ+2TNCM+ux4PPwT8v2V4LcXO3QMx+hEe0DrJpxHz81LKcBKoVoVN7g0D4bXte3ZZ7XOWH
m0bZ0OpRNuDvTlVn3ZAm/6P86LtCQGrgEO2OG8E5wbwfaoyaUEpamIawlDqrZwlsRZZs1HRuOeUu
LhdHb4XrXnyPP0FOvcKbl50DiER9YJYQL/RIF7H/Ihmv/tzepWDvMikxxT7TI99/M9FDsZjLJvWx
O/nWC/5hoHzRj/uMBTHSkZqpQ4tzg37wOPMv1IKV0t0AoPu6OpS3/cCmN2CpCLjdwsJGEAOlxyf+
nJeSdWxml2WN6br3PxLIHSHI9/zNI+61rO4XEPlQ3/s2k5UTn1hj8btuo27jguWmysk1PbE9QhFH
E3PuqWhV22BRDbvuUmp/iLp37BIDx+Hlm9coIxuo+GwBxq6lk/4nyJ5Ha7+ZU8s7o8E8o8PIH2vh
TE5hgqF0gmm4rySrbhKrb3pTyxLn3irQrYxSnNAvH8Pl3EPRJOqZqtv8xv4leSMI1Z5oLkDR06rk
UV1TwHpdVhLbAwfoyHYpK4dhP658FRpsIf9d5O3W3uj3u85iYJjfc9Syq44hrB8POBgG8ZLwtToI
kh1njBWLx6NvNwtvMbOUEqPsb8Ly1B67jOaWkVHX/+8e0DG9hl/tqp/lBUuXFw0i8wnCdkv1pD2/
KI0esdhRsVqkHu2ftJCzPCILs/HLupZ5a7kvEF7M4HiHxYXltqUDD+KC/hTkWeHsfXIT9VOLVe0c
u3UYiztj6+xgLCoQHK8b4FB5njW+GjBVJeIllpe0wVZQYC+iPkz4FT8QL++OG3LkbVbpe5PUNGBS
mTE/Ykqhv42A8fBydn8RftNjWufD98+UHGuvazoE5iW/IOVB4Um8cK2eDr50jNmB0Sp8U953JU1k
SFrLuUkl0rBN8CYKQbJF1rvB0H99BpeFgHmkYeVQXnHTFmN5Ag7anx3bR6UXr06D5BiMs/Fm0rXK
7061uSftOzr84JEaXt+KXg0NR6E3rWs08e8jHhQW9Fb4RF9NDwsTVoGtM9mAjAjMIJQuni2VASHe
1ekrm2MBH4kB3kIOXeiaXMKSWI5VBnAkyd6lICVxyysF9/GZBPXOa7ZA6/wUEHrL6a/R5vnhm7mV
TnF9HRGCM1BQtUuf3i1ABGO8OpAWopNMimp1SELQPCXMwZBb6uoAtMmewXVbYJ4KvIPt2tXlkW/l
ZETRwQyftjLIoIKM2u60D80sX1CWeSY+50AX1ZCvtOOjoTFaFEoBdCAMgmJSeoll44lsBEkLS+Fi
Wlpho//1QUqLZb9vY+0UfDI830hYmHw/+2tdT7HE5zjvfVHH+Zmjj/bxv2ImGgWfGfAGgG5QfKx9
O8ZAOr2IDdybXaitsu0TxJaxmobnKEu9Ue2WdKABqY12JKFxpf4pwjCT4T+WONE9bZHlzgYiV0YC
P27Oge86dOrIkqyCeQ3IfvCRSieIuZpta5u7F+GqLhb5K2NNWBImYFAKO1UBfWRoPDzyDUZEQvlh
ayP57/veOPr1Uili43PjaKicFsiWd1Z6GHQHX1dyy3hmZMrual4a93S0h1lkwrNekamtPl5yqdKt
UArG/MuLL2qmEC/TB8L2iOjUWa87YTY5lH10B6eXOfQoc58M1i9zntgtbmJGOJwwCpxeXpmeUd4V
QK2KTbaqO/u72cMtd86N8QgV6sX5eD5dyyDJ50fvPnTBYS2sYj2Ue+3r5hazvd7sm7otvS/BYI2e
fv20DboTzucN97Yii+hhTRK8xXpITO7jobP5ptyvOnCHpb9jgANFJuCo4wV+yGjwF7m+sLa3UXfh
xDkP2gm+5fX+79gAKZYMVd0PeL3qytMsdCWx+E0jAlyppY/yhwr0BQW3b66JZWXSXutTpxX+TNFI
ohjNr7+wNLZjVvMS9uLt4cI6+ULtJku/67LDE4sT2gp/6wn/7RAb2msac6llJBLN5/On7WQ0XUT/
hQs2uc/z5vQdDjjvAhdXe4W7+oWq7UnurJUO637IrbwVOOY6N1uf2nr/kLgkEsLUMnD+F59cZZgV
X93KiX9HJvj+p7NMWU9Seu6MogTbpajt5uevqeTzQHXuMFHUymOQHkVcgE1S/P2JFv2pmhHcFX3w
TE9h1xKAAEOA4bgPclW+q6FYsUhuoUSjKM3XTg9VnUTKPvwqh3YMwhlDi4GsL6d/Ja5KDmm720E2
ctmySaW5+fl4Z8OEwN0PY3b3sIIannlB3r+Y21LUzkLkymlYH3Q0lJ5eWfAv8PTFWgmN/pQJq6si
klf7hDxs/sVR8iV6Orw5kbhj1r8fdlM+E8QZ/NgQiKZRvqR7UlY1CUYJ4FFlUOkfoq9+sEnD58Ny
Dx+AQ0C7ucrZZhXeGSoA7QHYQjYbEKAF13DbDGr4yndRf/NBgkKIR0AneszpE/09718CKnQsrEEf
oC5xPgXW66l+eXR+ahSJpgD0NXteoXeLmCOcSNnzxcQek+RApzopCB05PfUjiF5ztZGYxYU8QrpU
rqH9R9XRX3vlRiBSRwdOgf8DnXLQAEHsr4KrFWiscIYTUmY5mjhWRMulUGvjvFpj4eGQ8v2Q2ZWt
UWW47fxun+XdksbbgV81ovjMsNaqMg6XVCG77fygIyin56G7Eqq6jJz3nfzJhejhSVPsH/JSDFbr
cZ1RCo9fFn52iiZ4m3oh7UN8XE1AJgR4Xt5iyDrJqV0H9EKHxa7nuqb6sV/ws9IBhxE47lZT038t
tIHKj3BieYswYKmUFoBJIY1+8Z4oQ66g5gEqm0o4ha80pB5OGtAu19SdOOxiWJeWWZn0UITzvOLE
7Y4f/Mr6HKBDGHJM1EBFydRjEKpWMrhMR8zVn7rz0bwYJj/nKZqVCbMB2lvzTNo2+6jFRHv9kERD
HQgVh9PB8qdVyckeJktjD/rj66EfeXXX47VlTCIHIqSnksxriA/3f3vQTRDOAn5+fo7831KJF1lg
A+Gy6aN5SrI3b0pKcc4KVjU43jsBue0fy0qehN3pZcKuFrjXn68+o+ye1YG0J0BLTAzfhYAtG0wG
tJfxN2k0uwXtBc1Rwlch6YM7r84HSK9ylhFgvkPxsdsyMVle/KA0fUNuXBFePndCOzGpNBCrH0C8
obBA5y125c3GuR9Gw2F+wT+Dn30Czrkry3ZGZl5gXUh68H0E/gm+PkSMU6V92ts6mwB7RusHqOnT
+Q6pfL+Uzo3hEN7Xz/UY4L2nj055QoIhkzomef2DRAEoObHgiUcgFrMWquSj0kqa918uaB7EwFOw
DllGd0nMHAXm45HUjTDnYMCf5epUfrEmekYIQOBXnQJKTKISEFKg2kWZDIpVJbHdpf4bSDTq39wf
K/Za/9g38Tkt3RYA6YnJnF9pe//kYmJTVr4NBlO0jtFDpLy0ACIIP4U2vnowivNyCXKpceacj4gI
pic9GU1SnTVOseqxJf0DmYz+jRXT5WlfErF3K0LNHqdgbjfbj1aWkEh7+zZ6kVX8cXnR/lcNtKW9
W4X5Z1KFC/s/QLvW/FQ2HSX8dtGxbFsDwK9N1h/uJhdCHspiYnHUp1ITpav8TEPWcvyDovCrVHiE
TRHABbq/F73ag4GjYOQTyrEvR/1RKycrAB2AnPTkrwxHshXeJXzg/nG1sd/E1p/F9NB/ERO7Mhlf
XsDBQBzZSFVUxK5TRgxSkSi+wg7W3oFgGB4dIdFffVpwSUqaJ5yhK8tbHfPcSLQWW/ZoACjy+UWF
vTDWBqVs+M6jzRUUZuzeST36Hl+Y99ca0tDf8en7wKxBIpXJV9P7SZmnZvE8J4WVXZ40P9OmZkxU
aZDjH36FTY5TFelwI2Y/3VSHXE6IcNSZ5kUAaEyhYJCUmvED26NuKEGSOisz17p/CgjY+4qbdqDj
UvsSxdqBzTyxxBlRmmLawnji2IR2Tmr+/dLLT6TdriHrFCG3WCo0AQNHjSBk/Zhgx1LDkYK1QRTH
3pOwGYu2WF21p7Bsm1Rjz4vUToqUBNwXolT3ubH3R0MwlvamATcaS5I+mruW6n+Db2w5KGuEzMoj
LGpjv7GKvTcw71KVjEm5Sckj378gr1Q/usm9bOgjTahIWcT86+JDhOvTpYUPjeqkiRBqEYWLJKHg
8VbSx1oL35XxDTBP1RVGuKJF+aHAEWef6s+CuWAvzw3oxRx5sbWFApNG+uGiJ2QxUDm9FRUAbeFw
IunaBIq8s7xqSAbY2eetHi05W/xjJ6/SVfZFe1KTC1idBDCxCOEZVgsWtKb/SZWk3UShW6gIivkM
TAm7uNkUM2Z0gR/ZFABM8pG+GnBtLqhqCS+BqgDdj0wwLOfx34yoGm+0Bfk6EFQtdZ+Bn6ZSmVyo
Tvoty7TbPobrJO1mBDioT3oyzqkNfNTMb95rspOXaBbY0X5x/B9f2y7sf9nU7XjTSe3p/gc7OY3W
eX6iIMc1P0v5Ok5ZdU10dpDudCFuffiCZsmOs1p5330uh4yiETyhA0OIgSOXW1YAtNQS+WUYJczw
VH/+KxJbnqvuaZj6z+2CFMp8I4FxqkxuaDOYUpc6Pq7ztKZYoQsNg3y4ZLIxCmU75yCQlABGX7Fp
ZO+2UhwsBALavRqYC+P/dKzYHZiJBb5MNyrMbZWDSKnQJHs6VkPY7kCugA+E7hIza9SE+K9mBwSr
XxTHG7Agl+sGm2hvW1Wv4OhMPHjMilQkDlgpB0SSwf2/eqsuW+HBSTjubm3+A7xbzpHW91h1Atyr
Rj0Hz1cLLXw4p2zZFzwk1XgpvvLPvZzAmQQ8PnNCOrSEtNXksB7YfDs3NM4qaig90265yo8wCi4u
ziWdT2NHqiRuyd5SBPoOWXij2BchlLSfm4sM4QjSneJuIwxozFbfeyTzh8nydRMnzUszfvvIKX3Y
+S5xWVwDGrlkcjPBysK5g2ASZ8jgXVxIEPRFzsNrcxu5jIDZLcFP24tT83eQekXFAlXYVycU4qJq
B52DIcFVCVMw7jcatV0hWeN9d6197cxUkpsCCZI+6nbr8uJBtg2a3rpzv+Fh/Av4L6QLZZLusthP
3zZ4URQ0avRugvcuk0zCqqKqQd88phgRybXJOjoukrEQ2Zb77h7YkqlU8mG9awsQEqhhRaYLfwxr
beImLn3azRlMQRwYsSyos5GStrWEVsnz2Ez+uHOvScFId07Hlnc37oNNFdgFJkH4PH5xgvEfgkql
KxU1z3FmHU6W3oDdmIbXvgCTPd4TnB8sBlWjhWLeiqiaxC6UMcBxcYJX3ZVivJl/GDHSKoNnrIeI
HlY6OxHzcUN8PK41mTFO+gkleCHkrMhAiVUjntg4Ry9TRov+roBtJAL/g+zdiKSblzBXZ2/Wp3sM
zFhM/bNqqrsEDULE0OKjcXdcxPlnWbE+QRlj42ZOvTRV7KcpOKOx9WH1g2ohmTELn1JkudcPRKhL
07Y0l8fmGo0e+TBeq9CY4SUTIAXuRxyRkS7Dwv4+Z7rV1txtdt2cyM38orWBhfVoWzmxSEzxFkN6
jbXiIYZKy5+fUcUEIgxaNC8EdhweFYr8BVb6RJcaR5dF6BW0VlSswA+xFA2IZSTV79ecpxahyNVI
3ZDrlezdzJyhrk5hGju37HoC5RFTkFMoexaiB+/j2sWuFR+SVUbD0MvNNTSbk45P2y7iuqWxnXiD
JXQWS07u36KTGa9pAyCY8YuTsKd3idmE/Bt365Kh+zNMdt7jQ/jVrjwYYSH9wIBVmKy/8j9oTzc2
EnV68jQ9IG5S6uWDDXsJURZivJpVQQdakJDFXEY8R/XU0FtUcrY8g+vgmhftdEqErV1gQ4WFdDyQ
PQS2GGCiUIVBpZRIju67IXGbVFg5w0oCb0RfLnj5dvadTYhGiWD4zBprAPl/mVbf3DG4csWdGyky
f6hvOyw8R83IaWUZgWv/wqoqjgjcfz4/G1A/8tD9BcJ6fookFvW31EZif3wZ2h2HeDW9Mzdpn9uh
HAZylmhkFwvHceMRtfKSQBWzwr3cVDOEIpfECLxy1N+fBwmAoqEU5vRdX6jSGEZRqUC7Qel9a7JX
zzg9HpT00agxBEKgXB2+rNh/oiAHrt476ySU4BwPqWj/G9SYFMDp4cE5ciGCAH7TTNxCQ/41nbUf
MIWRNMUu0wBAt2hTMUa6zcJZ5mMGA/rTRQeZ0+5wAdBJTcVxsGBmNjlKxX6LGpRXkrXNP6UrBF84
i+0dm0uoVS2dGSSPLCveBcDo14AN2bXPixLaDR2HoRB/ZW5kZbsJIC8Yf81kSFu+jWCps2wWeDW/
1jTTSoDMywrWCRtnIfiXmPu/mTVfcP2uIUljJ9yP7KsZ2sRc2y4+Z/jUo8It5YbzuyAOlSidfeaG
UIgDZ4ABQk8b0BJTBqNGoR6YBVg1XxAqj8ud+7gK2ArH2K79cXj71BLj3wYfhM8stIy9e0/NU6j9
UdaCYt8oC5Zh0aZt265xzmHfGL7BIzdtkfkxZt9LHljjv/J9U/PBJFihvo4r8oVbTy2NdEwouCvt
ayPHSeNBNqn+W3TmfBtUPjiw2pavffl9ZX/asmtc/GHY1cAFrZMZ86uII7yvcIy4KPgYMh7hVPT+
XopPG6x+HLB3U+lNa0nYx9mmzE9LkFmgzBZDN0DWm2Dwjd+E71pEIJgxFstw7D1tc67rXF7XY5Bm
zvTqF5Kx/16oSMHTPJOrpfaUyx1wWX2LvH3QQas/EvhGcWOirTwqeehqoApqNT0lvsBuKyKfd9EB
8Ekvtj9zUsKoF5E37fbnmswmsAQbuIsk2IxXa3seEdSGkMbMXgob+GMSocmdDqYJCcqp+jNskNZR
IvqOrR/zPiN3kSG7HvNNrlcJogpL+mxX3onA3ixp51wfJYTG2fMUa0rc5pkZc3LEpTVsLmBHnY6N
hOmD8xHlW6KsbZuaQNrYYl/ODNRB9Y0tTvMScNXIg2aOh14izuw/KjUE4MBZL7bUFX2WjPmj7kAb
oFOheMC0BLQQtv2JjFGpB7JGzN5PVohb3v8vw34dDSboGoBzFidXUsE422zTqWFFH8Y3AmEpmaV8
f4rEGsrb7ZGD8lpuNqT5nuDvQNOdjjwezHDWD3R3iyQT3ZHoIW2iAFw6Gga1vdneQ1tRqM476LXu
xV5T/FJ8Wy/XbbB51uQRkk6wusbfufr28vYz4OpcGwxpN4I55HurJRmDYAwZe+KZwA8V+WT7qF1V
xiIEcTQsys0jb41skY9yRIiC/uhyoSPj/VyWfT76P6GP1YdlA/avFqZ6/acXUqfvym7QVb7+S3w4
ltX5EnlAvMvGFLmBGy7081vMv4sWSsedXgToURZ6ciNAp/ZhAgVmXvyVgF1FsjHS1BgugXRZhXH4
31t8FoG6uiTQ0bWXV76kZb0lFCjWqzsNr/3GqhDWblEH0T5k2Tbj+31u0nkOvYcqlsPPZGu8KiMP
mZ4Ls8iYt0Tyq+70iGswMOzRv3rkjkVqhnS+RmH6nIQzMPcEqcW20M4egXEGzTFxHM7oQWjzTY3M
0vez5x4XE+dhB5hyLf4l4J75A6DA0ZPUO+5h84S2mU3MTI65MUaozGyd1EWvMjyujfvA0Op0dFFK
XiZa5pAWsV9SEyzAPplHUlg9hUKBibsVRdVHPkJTjyxYSunPgif2o9a5nvrTbqhFJXACEdNRSPTI
xhb4nU7Fkiyx0fg9yiryr3M89kQXCjHhWz+6fiWl/35BckrJ6VjwZpcMWJ5ypTcndIqgGjOWOdVp
X3SpO9qzMcOBPOqGkBTUobYmnEswvWEtmmRLgg4jp9Bibok0ErjivtGE4BQzHrF9nrAvtNMXtjNV
JroauUFVJciWfCxVFwi/70hA/6U8M8hWqDLuwSsRoet/cCPAXxGWDQnreGbOBwFoN1JVKt0n2eGp
K3cVIJyK7rLlbgM1ER92ZwXRE1DLOLuB6vaTrCRob3XbmNLpHzrfoIe424nBO1GN68Wvrd7ibsbU
LeFdCNdZglf8hJH3/jaosEJrgZ+YxEUg52OOyseFQvdxEcXcuIhjqOwCWwCLEcEa7XsCcVg0LewD
naev4QW52GvAICfXVY3sE5MSkH25+U16MFyw8MOA7RB6c4Y9J3Bl11nSGBdvmAD9QKThpNkTAtCT
sfG/S9rkV/FLJZnu2pBKA77TK4YH2Sx5RgkO2cexKTRbxNHWwdwYThRH/luYYBvEG+jGOU8iUzcT
HH0yoFPoIu3/eTE3V+/WPfuCqzeD2x2BJtkoX7Uzep47Dqdh/O3715DPNvmF6QldIIb26DNiIz5O
NB+LTJ5VUBiJLMthM7Q1lXoP0uRLcX1CT2KfwJTJaWc/MDzUtBDzbXPQvdmFFXn+vRIC4PTpR+1N
IozZU57jZ2Z0qgcVs5Pn7agPZKDcyesl4hCP5SovQaNoumZcpE1at6vak69yPpHI+3JK9pqSKa3k
3GE/Uj5fZpIlC1gW2XJdzBdDYMlz/9YX9NLyKDcvbVulcDVMQV5dqqPVXJv/XJ6iwgpPZTw5UaUx
4TlxkCkd9u8xyyV6Ivd88evMxoAdaLeTJemrLp4RMGjgB3eXifYhbFUq7sW99IvuYTTSFxbgCR2d
cp1T5c6dG5797KGKIsM5VJfR1+/3tyc+vmyWMeQFMHJmBleviQ1Xxqq3Zz16kfx/Zm5vVXaP+Cml
qGFS0HfanY5G3G9ojd9nhIk6ThpGmKh5t0kBsdh/Q7UVt/NoIp2COVOLlbRBtuonAuCugulyGFiu
f5ggKbUJXLqIf7CnrK5ZkX6g0nvIlZ7dcmE84yC2fCRhc7fSYUpx/aWQimYaq7Y3RNrFwvynTdsZ
yPQ1Dm81a5L47ZdPqzq+/08ENUa7x+GwXLVMbMfzob2wnFIqzcdcbgj/mKr2MWIqVbaeemCwn/u9
R2HFutc9G6og7bGjR9VuR9Aemfkh/hzby+an9XKW6NVKx57LMfXnEI/jHL62iQnxV0Qh1exSTj/a
tD/QgdYXEs+P3XR/FazS+WUf664zoM7DlqcZyCQYtNpBi0oKhzTV1ddpyePxlNpt4aYH8LhQkcVu
0DE5EenvzHUb31je6xuOlzwJ/rKmOzB740CBCFBWizM+5GpyTdWYJ+uXvnD6h3cPM+D/JwFPHCAS
2M19EI66Bo8PGCBeDT9/K388jKZY7zHrjQ9K7xa2GdkX/LLPkBMQYPrSGvm2NqV1b8/KVNXCBZMq
CsjKVP+hqxKlPky6d6a/ulSDGq0pzVlJqoY5IoHEmvnRabcnnS5gbMGtyKGMWMx+pGjt6tfMJLOn
szHcH65QplwB6gHeiKaEj8U/Oz5YvEuU6txCMJvUQuJ3/QpVpf3m9xsL9MynBzlhN44Wrc1Atulp
Xep0aRN13k6D/MNFX8ykNzVUCCmnAWFxhx/i+B7BJNztY4q+IXBvlNvbDVIyvSHkZkEtmk08P++X
i07IjxUuqfd2hnxNGnmqkkds3H6bnA4WHJs9buso2tXco00dirRnLS5AW3u8b1Qkp8xL8i+tGafZ
vQIENa04eIUjTB7W1cLjx9+IvMY7OIjIbmA/V8WhsmiO98jzhiZXTw0H7fMQr4AYHDOoeI+/FMUE
LeQLojIDhoEda6mtr5Zn42D9RGyNjQBX80VuwYiU/6xkpOvAVpN9PTMqR2Ui85DemUb9hluqteZy
VP0fMrkPVMdj0M/fnbHYysBXfz4eUbigZ4xKiIj+5WMoKT7QLm5WZ6ETaX9KD5JDV8MwUwEIe1S4
E0+0o25eSbJwu0we3byPa3RAgmBb34LOH9Uyzw35mH6qPooTIqnebUEoAkNHozWo74GmImD55rzT
s52wSp5t72VMXx0NzG3k0ySgekBW+DCQ+KWDVn6EAJ20sz+Y8G6yMBgwBS4stKRBt4AFryHBQ5oc
f6PT0o0d/qLiukgmcle0gj201g7eSc6GA0eWAWMDSCgzmOn7nCfJC+tjGVvf0EsslARmVjbMaJhi
CfojiaAjNsYdULNo58zchy57VjorSKK7BoM2Xvjv3eyh6fPAZ1lDZd8ZypsgW59Sd+V1aylSqNiB
AFJHYGTjQarnCAosOfE5ibWc1Xufw6/0eOjd76HDJCdTl9aVGsIkQu9deIYj0m0sFl64sE+Ug5BV
wojHpYbb8r8b8czKOmBHudbM/5WQVfCBABOxRHAWVLLpCcjJxluxqr/TMJVR4XVaT3NikVsIVg+e
/kG0Kqgb5ltH5Ey6zR1FRQVtxT8IwloZXlUCFFHQN+zbWpGyAcO5XYvCXYJkygkLL0+gO6XD9KIc
l9zVAYF2LYCHJk81tBlnqgLSX+NbC1YjcWqwYtiY4Tuen+LhRcH46DN26Znaxxr/3RN7dptozYA3
3EdagwX+Dvzwp8F1qRlWPekPN6Wwpg31YTwS5Lh/re4JiRnYgCwt5qSj5J+7u3MLJxx+Qhnwdskt
j3FCzhwEFCl8WzBro/pSJ9ilmn4OhY6g/j3swVlNWpXzIm7fx61MMKxZl0DY9fJ09w7FLoMIFKdz
Ov1ayUQw7AQ+J5EiYAiGENaLh0GV0lCw5tjC64g1Zm5GeHtwd6DfozyFLGH/e2r5bMaWTeke7wI3
m97kd/QVuoooDTKLdqkrzEVzAkU8IBBygUB73Xh46t18Tv4iCGLXC07d6OF987FtVke7qPPwD0pX
9qs9K3SF79D00gHXBGQV/6DjMruQHHrPSD8E5DUPoQr1jfTU9iYlo0dmOprMhOU79dzr7GNygS/Y
zdkZRpu89POmjsnM1AetRfoByGY/tYAmcuKDaeD58jEv7X2eUZfAFF5Eudx2a+DemPgDbgCvk4wt
TTTVhexsYUvpb6t4ZBCajpwuWb8XD7Jks8iypnxk5qSFHUMn2hNTb2cNaoidJ37KzffIt3q9J3+W
LOk3JnxaMdNzNnAngSumpTSPoL/eErRiBJkXFGUrbDNuCNzFH06xCpNIdnwzQHg9a8RfIF2zTJ7j
gbNWQbsx4KXj/42dLXYmlaeE8YChsOghGooIJBR17I42HH5mUj4Pw7TC7MRi3CDu+m08JM0vG6BJ
gln2SHXIQ8RQ0NsOMn59/io5d/AwJYlnqgg6rpKBbgUGNdaCXPGRuppnDLx1MVTQnTHQH5HWbnAH
CYHpWXJO6j/gJrfCiHZMQdi5Sp38uwhIfIrXoflSKHc34HOHy8xxMX/YvUPfG5Gq6njRRHaajmLe
SOT4yUJQ7zWSxJHEMNR+neHJXRIfsk8fw5DremAjwMhu45VsIffPHbSAz/QnHUzjDLSDbVPBo8B9
nkDFFjqH8ZvTl79kn94SlbbpOM935dp1E3moGptKHs/U8ghIVNsM9Dvc7gTUAfJ2hGjzXyBIVLAr
SbxnZBBcpnoeaG8to1sC6KpwsiSgKgkJDMlgeVKcBUiS8aglsUkCMDPoR8w+RrfhLhO26MPMCciO
XMoOsDvPv2QoGolMKJuZM3Z05/93ROhCtPju85rtyHocKaV/XfAoo6IRipwtshXeJDb+l4ZNDom9
Wr+FWhqK9V5ejhGmbiTgHakjPHdFFjBnAJfHKH7J7d5DeSZwBOH+Yp+BydJMDAouv1GTNv2GNaIU
7/UQhpbIIuOlXcOX5AOPUCDhQFDggEch9mBwHXHyLFxE6kHZVLPmAnxKVvwoX84Cgtp2NtrWPyXK
EKqwYm0uIHuhGv5+GqUaoXob4KczQ3pPYIsRLKG6v8lfQ+Dwlm00pQIQoPMRDB2QpcQjtZTcYnP3
GBm7/QSEr6zqxhZ7G9h4iqyONPyA6z9GLgUJWrjGbpITdV7MNWkLs7u21xp4Fvy3hVOWeHC/7MkA
NCw6gZ8G0LbJWcO3Xi6ohtoBV6BhJlJP8pARstIR6HZ+v0ONx28bromfbuoKxJib4RLtXEb5M0jk
dQXDdWO6yEeN/aQePF0xzA2QeS+QJ204dyu0jijwTTFBNcNG+0fmvWvgjSmF9yfFMnKLi4kB0Tcn
zOyIo7Oe4yo+6YsPaYTe4SRJosksv/XOicfiHXuv543HZxfVEsaMQckut8bOO4ZpKy20TLfXzPOX
nBiZWcWbMUkFZHzci29M1ShTwGRnxDkJRGKnwPV9NXKgYDUPI2VhuGK6vKi47c58BCbL4QY+tzfR
paJ7e02wmYVQFHfgE4/+i8/1Rtqm4wUg6vskRx3RJnVbxMHPTTzBCdk2UpsfYk6uRp+3N7Y0BQrC
hjoQ44qfog9s9pzEooyzbMMQBI96LzB6WIqxrs+vPivRsxSGX8AoD/UMBi18zSPVhJejggu0DG3x
wey/TBlfVDum8e7X6OFaX/vFmA5eqWeVa+PKK6qLq/DPcCiGrtrpTmT4syi1ZeautgQdHCl9ylyZ
J7r7CGlaQxkRH4H6I5QE1P9KDD/22ZfHonQ+lRrNSx+Eqb3Cn/9bR3PknEhWt0AKg3mV/Qaa2I+E
B+XfjqUGE3/rEbjTDdHfuanNM4/k2cXte5BUctT+4jPZ6sIcPwfVBDq+yzzwhzCgkNVGaaviBZOZ
FLuWR05gpJ/91MV1slFipopXjrP+XpFnBv5PTTTMTqiOUcuS7aE2D7zKDBXP5VYdYVyHWah+098e
zf4M3hGqcyI8N6k4unfBzlcljVEnS6Nfh8o8H+CUGs4HvXiqe/dcb2KsfAgB3u/L8G3pVtTJMg6G
XyPyJLq1bbVGBuQJipdGfk7fKADEw8JsRsiK+e8SWUa2jRf3cu0MgQIBlzYMEjMUL85F/lDLobeb
G5gxSlWS6KYcf6BbXzOo9VCbVddFS8JZGvtZ24KBRSyVu+CUjLplo19Tb6MJf3Tv9xtpRcwt4ZMa
E2fzRKVkRgiKmOkNtprej75IPwe+B3BjSqykVnf8iJJmEeBN9hGeWPyzNIjFFBwFNLBL1F+j5Ymk
J5N1vwzyxXcm8tVfDyn0ZJRj6ppR/+Oz88S8MLG7iXBJo1vR6rpBrHi7vpdmrs7ybK86IVnXf80d
qAK6MT3UWeEsBtv2x4a+vReQyUgUPYlSeaY6tk1Wc0xtg/L3yOaynxq/yhMcEhlKJ7oxKmV6oCSE
UiKc0ITY8tnBNfqyOPDgewRCDr5k7daNCYIn808E49zAHqa4KVaEyl9EtMI5HMmpOJ+HavZNI2Fm
d2vFSFxSoPWpV+wDDaO1eqK7NQBk+EHxja6bp0wtS4VcxSQgxAEKzLZatS5uUoAka6GMJApzPlVd
BKDXBdYprU45y+CIhya1uygrIV1pyjKJOB8rEpfMwmfxnI2YAOOUKv9NNiqQfDrpvHAqdBdpaRdJ
8Ghf155E+qRigOvYJsv553juKjX/IiiW/i3ZFl0jRjSS3R6HSfNwJjjnb0l3L7s5Sw9y08VWX4Gn
QM+Be4X4hYuLPH0pLhVRFs2CzP/wCAIwyDArS4T3CSYjOUZDkon25X3sliNT33pQQxZ7vyX5hvr/
lRHdNmlhO1PAQOrC6TPsDiu1O5+PgTUuRWlofYHVZF1fwPVvBVktf1WdHT0UTysmPqTQ/fdkvPHP
SQUSG4Ba2Uq2iMROlyaP0DClnSvJnkD0X3uC/buFSELqNc0xfjJywNnRXZh1uVUNA4XvJndSb87z
M0Hqx6kyyYf7aMvuPYN9QFt2g4urk/M5i60FcevUtPdNuAJIEYfDETip+N1pDmI7+/xWa1GtNtyG
Yw2RZoyN0BbItrU+phm57C8V03jVkKqAh9agetspCWOCK8gBoMyAzMlxJO+f9j/Yf/aKrJVIPFDd
Wm9kuYlHqzNoQt/AZvaTcB7kcE8yD+mmgaup+nJZTZnpTWtOP48EF1iIAI18l0XXqmFbKzyEk2x5
VLwS1ES0AXhxQJAT7fYCL+FkBL3rJ3Ni6/Dq4OpFVR7+XZlF55NVMHphSubPMX0rB0KEV0K7jNti
lBHEFCXjpubI4hjCacMSipdN8sNGN1NxqndOMPKuYffxMtmwrr0hq/XmLFnykUcoh//IGmoLMyj1
9Eq+1FktLVF05EzLexWPNQGEfIQg1p3/uLzf2V99OzMCHN1x7eYl5oJq/4bzj2rkZ1S26BVL4Rl6
WhU426LnbGrWDrX1iyM2vM4EFv8vXbJGJ9ZYJms5HKiS3suAetVhIFzip/rsZ+ufBlIAC8WaETar
1Vmf1SvpaAGwEolIm+YNult9gbGSC8ZHENbZCqE+qPhX/VG2wdddZ3FpRiXRWNljbMdGj+QVPwdH
P4brtfd5Sow70qJ/P4xsTRJuBODta482yKsggGjV3trSn19u9mdrDVkKtnIV+lVA7naKi8xPhYtQ
OJJ6nM5bz3xbg3lqF9yaakKPuPWzhmRgt1UqLcNQm5pLkrFRqqG7OTC9BOr33im62m+b493PLJDt
tJhd/z8RMHcN4C4IaB0kkiGLh172mgpHJXRMRJ8BTdAPF9MxOayNzgSsg/WWP0kt3ysRsEcfAqJM
f7B8vuaNbvUVZOPoXvTXjj+vuk3NC/+8S8ylG2VkV0/GHPJBRrKKfJzvH6gp1u3QN/791pnhKVoi
H5NON3AZMKJKrny5eAgy10iaytc28sapFW6lObQiCAPj0YpcAKo9lmMsaCO195tXEW9YbmQZKi6B
/Xdxq61haShBKc82pWAits/q3M9BJwtke4sj0GG8z46O1zebiNFxOmqE0yCSHzMI+eM+foXmFElo
cxDK9x7J16UjTJuiP0SlnrVshDhBi8QIRFiihKUzbh73p1Nrth2D7x4h6+6uGGvqk5fl61lCkU9f
iEXowg1V8D1soH2FUQjcQzT6G5BSnJadMZ5ZiSra1UCXYLbIbnnvCZVBv70eJ/OMCk0Rp4qnNmOC
rmaBMdkvT5YUHp7TrG34ZMCW0g7t3GJc5agjuQgDT1lh48kR7uoC0WEmyrts6ajPIyz/PdxWgW9q
+5FvYoaDm75S8BrKyeFpojDTHtBvvIVJS0P3HJTCzUXy/avXK4UFZJVBHBf+76cYxfjw0/15TpvS
UZ8/w0iKRmXU9cAk72y76lNpTozi1sWmAXKEeDxg8NWYazg/G3NmS3bbrL45UpMuFaq+eHN+CJOs
cLccuw+02UH8YhaO3kDu0ckkQye4XVWfyrUUkfyYEah0kdLMMno+i4FJxKi0peMF7Gsv9SfmjIOV
/fqWHtIK0ycBkJX6nXEgaWiyX+Lf9929CDixIancX2wFos9T4Ds8Bz4HYux9Xk1MsKfkMAQTJAGS
ofnbcRybl9322BYDPqm2Lp17r0oP5dHs4G9jf0kHD0nU5iO3JVaybjIjqJFlUWq2RecPUoNhhwHB
DS0TTXOkFEw03mfPybpe4lr9dRySLIIfL/Lajea/ZpxfkQDzUckKla8hmV5n0mEjmvUMXEhWSjLt
i64dEkJDujL7WNN/4dyHGG0N82zc5kQX1yHh0WrMZBfJpkN4dOKiXRHeMp9E5UuD1O6JYEGqwRON
ZgIR7rJ8KJEq0gUPrcrbPKw6b6rAb3+BUhEb2zPufETlRFLrP0+TZGsp/DSY2XKyK/mWXu0CikzT
8C9Yc3CW/VsO1hhaDCYMZOoCc2m3asNxohycU+y/hYRyPdOKZPYRzCbHYPrPOEZFZD0mAvxVAwxN
JBXJlT03WgwnxNhSOlXtcsmwXgZRp1wKmJSxhulB7sZQ15AYAYm4/BCov/AE2ZOgIl8napzyFeEv
BsdKC/qbm4JVbO7cmAWB+z+x7/3ofkwCQs5L+8i5S3AwRQpQ3eW0d/fo+c0QlLG9Ln+Os3Mq9/rk
9ovx9yORbG97P29Z2LcqHWLlZFqByjutkptTwL6PBoKcy/ZQbwOzU4qJuHoZNguNcXEtdAL1epAc
UaYf3vhAKc+a8OWgEzYOIIEu7xg1L+odjvcHtsGwFozRKyKebSqzNF16IMNOs4uUYjDyndHI5VA3
dvhFUjoedN49mz2BYt6Leq7SDg0L5KOfV/kg/Ls/grMQwsISppcDhIVCxATQd/btSSK6j/TKLS22
tOvWYlLdKtGvCguWbYzuAJ1ey2ype92BVAtVQQi0QfGMwjHBYVJFjN3ppQUjc6r7HbpuAotWliCW
PuVQFDjeOrlfRNvWDbGLX7lfhcNjkdrZP0W4ONGxRocFac70juzrTWBanyih/DlMzslX0XChnByB
Vwi1bRsaS/R46wXN27E4N+/Dl7vnPSyhONJaCMIIbY1/VcBcdPIVICTdg6n7BcsXodi7XcRHFFeV
j07t+7pkiuTJUigRr25GZ+iQyHBBBEkS1DIjd7xgeiZYDXSw4rWNMHh8rxfGjoFGjaQMBA+jgwa7
z027GaKb2CXpTFwae7+wPTTLFoexYtom07/GFPrWt04Hu57IxyrJsBYwf383HGFb5PdN+jzKTEtS
JQjLDB1LDFRtSubCobNMlhsZtEbaFBji8PXkqG9NhWGz7JRgfyWVuAbfTfvt5R/kC6PaC2iXcXZw
Db/nV3PSju/4fSTuyU/ZbBFx4hHnAzonaQVEbPk8YNetF3XjigRD0H1Ofop+A3Y4K8SlPtKy1PBU
3iFbi/hl0Yu42arDRv+hsnxwlsIdV8rw78YjCK939BCnpVxpu8fx0rQlwptNaAMcyWyuRYNaUGb8
/yQGEr9b4Y8o7diitDyzcG5QfKpLRJc0wPYMnhoN26Tfsq3bezVQTqIR1VS/DBIbWRehuQ/Ke3Ua
Jjv3Gt7jiuHtDewkbOmGDUywcc2c3C8WNSOlPfPtwQnr0HDcvEV9WmJ7kfgfAWjRNVajVmUxZqqv
ySe6CYtBpzEeUk2h24GsRFhKlWmjEQpEofbA1XBesY7BWQILWVsDdydyXTsIimhLdzrHNGFXAbje
0uHawf3zdsT6YfBEa1AwxEXxuH+sWo/5eReuoPYfZLgOc5WmYqfxlWLNlRMCTfAsdyquu56RWEXb
3QwvtjCDDAV5CrI5GLhB8pLnPSzg+G5fonFXudm4lLrr/q10Nh0swOjwOjFrQvK9Z2qhgdK9tKie
bnkSKaFPbjyYDZL27HqafhZ/0Q3CXEIV1sISDenak15LeHRXYN0Nebfxcphk8GsL/ZfU7t5F/lL8
X9df+eBmNTZE9TCnXuup3W8S7FnLdkpg13rOWtNuoFZMkv3hy4w3k2b+Po0dOlOmN76k0tK0RDRX
h5dI+WBeFhjoQX5V3qOHeb935jxhg2ly12IowuAN7HWlrQgzC7qSP9lAAhGq05H6QS5w0ilI9sGj
eogMYXHa9s9C3aw5+7tf/nYTkGzdGw56z2BSsspUtrZZ4qAhUVrJC1MKc19k7GQ4pGLcJLTe/Jvb
zM0ydRB34QIYudq55EpkwySD57kksCj3J7VhAlkZK0FV/Fj+g3fK7LXJ645AVlzoakFDQcxycVb5
baJiyghJjJvAbgpURgC1QBgfJu29pAipdPEGZWGysQIFACYZKRoZZGJHz5RLQtOL6W2YyOP25M4u
KwwoQ5iyy6ftXstjNP1lDe8LlypXDvCPCUX/TMuWYoMh2OYnnRyZWVK9ss5grXNvualZ+jSaCXxW
Yu7y4uVqdcVPDB5B515hWGlg9dJa5298oWW/6DcSgTZhlUf4szyLIVWzVM4VJWBFkNtci5DqzRJg
8G3cWi4bhAUiqAzVc3FsS5vuZ6Dj/BCu2Ie96Y4+5fi9nI0jsKJwNLXrLQPivN3mQ2MuW7XCFWrE
f8zhZlpK563Ko3V7+mtBnP1nrgHD9Jb5OgTCgYQE5J3mT+6i0hfs4rrpDbeP/YNiSli+N55AJEaf
C7SMQ957RJCLevC3JoSCFYf7rqo+zORG4d2vBqg+NYMdptK/MWK7Jzl0OdCzgLEBZa1vHIx4/GSm
BCkdt0sVa0WcOs2eBQSQ8DfbwqKbVyj7n1s0O4kUcptPq8C4n+7p6DEdrOIFogsubxdLJz+OIBB7
icjvMoWP36Z6zjy+xc1bPI9vop8RMffmZOnzE+MmsxxaBNxUxUGKWvdcjssGB2V/Kg22VnWNebEb
sjSnxwFp7BnTH7ne1tEqDSFuqHF0p9U4pVaedEJBSR8TVXRI0sEcTDVkFwgTluysAZtoZh4K7Rah
KnvKTVF9Xin0spd0OJrXojNeCPoq4hnx0kAx9uM0VjiYBZdF5ctdcpc4MvXxWa75SWagL3g/rP2v
dftQ/o7KkyPLYKg8RhAOuC9EceWU/irqUsLKuK/CEwoidOfafxI1JmPO3PW9cfc/DAn7pG+xP4Mb
mYAtHHw24vWynPownEYb/xyPUtHSnXWsrWKk+J96M+53fR40ULB1yIACqc61Fenzi8uceSgod266
Ymnk+2MHK9fVDGgGUlr9zU18K8sdhPSoky2FKNQa7TnuPA31/U4QylSfQ2Q9y43DxZrjYiWaRdHp
dmCMINOgCqnIBCy9A7pvmnoE9FijAigxFEURupdOE1es5c/MHLekXejiK2TBedFFsW1Zihj0P+eV
c7e8fdx26w81QI/0wiOEVaFzmg1AvvjnujOK7qTgbCtVtn8/0QPTGqlpGKMffO6JZYTSER/oGOZO
CrQuyL4p6OFZIUjtqu1k8Chx6BaOrok6kbwm7IqioUzz/eHfv7oTIp+5foJwwl92TsymYU++NbVu
iRgcBtc6TWq81re2OfvEmoFotC1ab0xkPGSaGCZUSTFE5SL4vtjCIBdlqF+FVyDrCNZxL6YWZmpJ
gtW5fG2htzbRcN8kbd+d6D5u/G+JkpGXYRyX7iSstpSZttRKJ2SFhv/X7dBO7Edgm7xuTsHqAsQX
Nr9kRb1vjqNfjvSEBUlMrlTgl3V6p253WzznF0cTe7h8LLXVisBPNM09wqK7TEQDdp2epTstOHWf
yfWclThhKZJp/VN+htrBjwu4zh/WuKEbnHpdDAv0CgbmGcvi/VbqHgx3hoYlLGn6JGWeThLbzgmt
8z/xr58f4EMCzZ5cxC+IfdHEDJI0qAqosoKsMZQ1I9Pb/jL4IP8yEvbV/HpyXZld/pkc8LtJe9RP
RwtmvzqUTGYGyX1glnX9W48BGKDnHyloo5daPEkNI13jKtnrjJRFzeXUZ0fIIrWU3w9RWZImSqtF
rIuGlKV75GHHPztuMNdPF2IQUVyrzXPD7rtnc7/MO35JYRxeo7IOlhRRWXKAqkPoSBLbmiiafMH7
a/P2jXCxFuGuV+ovaEeqChvc4JLuAvdwogMD0Ge/NOT9PVgWvcoqfc8GtWXI1ALBXl2LQFJZGTLR
r0pPgpBS1/cpFVSNUYBmWwz6yeIw+ax3WqdqS+FlkXzjHXv29EW7R6yTEJwchdjdSxGaccoDPmoq
+4KOg3ubr6i61Mk9XEqPgZXvh7L4fpFGjP9kel5LW5vFBwiCpGj6sB2WK6tNaKJTn2PfaAC2VEZG
vBj9Zqui3Lhlswl75/qgMpch2zedmQ252x9dhOE2zfRcU+TkgfwE94uS7ipp8dwoTdx46dcU4LRB
cLNS7pYMmJueShtSqJAxdgg7/asEXkfYzdAvBNje1i7cs78rZl5s9/y+rh8Qu3dPaB66KYB/hsf2
e9eHN1CIfmKFKAnmI3KZP85a2zYw8qd/RL9OQFmfbZYahX65MmUNKJ6BHW5iN9LZynSCV/BpwRRT
10WERqIJvD+sggRMcnlPY35ylQ47XqW81Vjg1d+Ei/k8kc4F2uwTilUVeMajas+ojejHn7cvZuiP
XFOi3i6fszszLODd85fnTK0LNME5qH4f/VOSRtH/qfU3PHu0lX7H33hYzskJtiYXawJGj2A26MHa
mHdKLQhEy0y5UFqiU9T9A846maL36K9sm0ezOTLxDQNa7DqZm2pYcbu516HUNWMFwtWx7oOC7wSl
Pqmtzo/kbCnSIE2xW6pNL99z35yfOujo28UKpkBBfyrJZOKsMh1jcXJpP6R9nMC55rS3lZmjYcH6
R+l7c0GeuOuyMpo7Pj8cnlem/Rb5luVOV3blV4sU7aRitNNbFEnIPCLsymxFsTHPB9LBLvDrJdXB
XX0WEpdbJdX0c8ShxQW+hPDyYAgYN4Hymo9LCsCn7wmgW0+o+JT2Jw9CBDgDuaEk7/iV1rrEda/s
1Kct5GWzMHx7ax40/HU/vJKOb24eQN7ZkLHrgl2UAt1qDyw1LQU75yjgKKsCV2eY29gRclhLPF9Q
ZkLYypKggloq1Xptp2dKrQOekVNNp68DROHmBVDB2+/0Sexsg2VSh3qUcvb4NXq8vvXGY3uoapvT
fLsk3jds1ncUZLNLXidIWayQE+DsYAMLDxH5HWQVtA+ZpooebxCevAB76SIbYC7rvWxM1hWq6x7d
po9GPqRHa7g4TRcqDIqN1KMdhq8Tf3uyIs0phYpwBI3i/HBU+05U3c8D9aIi9IDQPa09s9QYsxkT
Uw5iSmixk7CJGCEquMyPtjuKnydYMb6gumBPysR/+LknQ+CBRtGvOLVpXnMJoQip1fvZLlEjGJ21
zslDK1BfIYXaxOBAAT8Mnj8op2KltLA6QjoQP7tiFyJlw40In4HtSQyOkvy25nKJRKoobKbosYt3
Kdw4RIAnVCPNnMWZpPpsu9HMbN2Ai6nyydaswrr9BmCb91upkQBvcEb6gsxASF/EZh3QT+54Cywg
TveZRnGWm3V6sACRDhrNaKcJM1/UIjSzvMsxH/ihiRa4m2BUSGEAhZQy4kuIbutkO3a815UGPDKh
81cF6Ouyi4cyNsSir4T86GOfimJpKUymRah+4CeoLBjm5HpT/I6PQ6s+N5TBcFg+yiOzpIqzB1X7
wKYAfDUzn0XHbWcqxbkaEi431NQVhVLdqVSvCg8EmrUhsThjCbsOZ5QQTRXIeY5CUbrcTZOwMUOw
COqDLxA7zg0OXMaN8ENUv4o4JqcPPo8nKW5WRnZ12yjVna0EZCMvncmIAG8gorl/o3EGYMmH+Q/W
FFO6kPHCwzRYWa3RM51prjA5Qz6XI1O9nIjV2MdOtLX6o0XRYdZN2TS17926y5oPzck+kex6h/xk
hbOncxklbt0LGn3v41WlJIhrTp87FV1zy4ofzwgdks0406m/wDWvCpJJhys65fFhw6XSD8sbDGJ7
8Fcnsl0klTzKczLyZKfIlmQd8VLT6kIp8a2WgXUJ0sIbQjO4ZOalZhxOQBDWb86TsjnGQVxnuxT/
Q+uQf6g6MhjuMmZkv9pU1TBHJeaMQIXll7665GlYgJfvlrwms3FVCKR8NoAT1iymW1Cx1p77ijdD
TreSv4lcv3l0bdUY+G1XLmdbvaV9ko450vYqBSpNfsvYTXpdfd/qhaxN6shUI+QyCL4CP9ePcBcT
M8TTvKj1m5ONdpHhc6G5uKN+vrlcgLJ64+wZxXqrlKNHP+PnGuFP5Kq4qn3yqjnCv7Brk2yoAvfq
z/eSihkS5gqZhsqf7hGti+w6A1IUT1JeStS9uggUN9SE19CeuKzzxqVKVAT9FNKkzQAU9e/aYvv+
UJfGIzBh34I7l4+d/trpEe0ovAMAprrkP8Tu5vrIvOP6FXo8kaXNg5xMIjvSpWhZDs9B8Y2kKwry
/ZN6VEQW/sUX84oGEIfLiX7FIfkTvSL8m4S+4pOWjaOUOH3hw1IEhQLLXS8/wh6QEP5iu1qEt3a+
DLfg5/052j4r9vM1BZasQ4dIpcz3zx1y3SEfHAF/dDB2ohBTKhFktmier/vzYF6fjr1mSvg6as4X
cO6y/n3/2nlZjpm6SDaydoSM9IMJUEmcI4utfzxs1QdjIn74A2s5wPq4kbWeowkkmp1Fuc0uerjs
cN6ihmgFcTreDDiBCr5FwOsk6aG5k2y0UyF7KCbCqZaPsXgqE57V+7WN29Onm9/RVCNhdjoxhRsL
VMbSLzgP3XQKLSROPdBxRbHnpMVL3z/rHqOMA2zKO+QxREKEcMtItBmCz50ibuZN5puHjVYhZoYM
EYiD/e6384oP5YGURMdk01jvG72PGR+YksTn+GOohQl5drhER0vvt6yXYMyd1h9c+09QyzolukeD
1sSawm2zbgerbMCSOzdlZI4ldzeTdLE/6C9FwYb6sA5wEwm8LEADiM5mPCfBQ46r93rDizPYGe8Z
ZQtCwi1joE48n9QjGJX/qAYUJKBLtb3JbXGMauvbOyM/1Cvyek7odhtF6ycNrLu2BaQ+eDAF0Dd+
UP3B39etFDYvOKVZGfEI/Q34TN2w60d6LrOB/YTMIuKp3trD/jrbqngZpx7t6ALZ/vqHZjc+YSCC
kGikAB+tMJJ+p4F7KMb7iPdIgooHd8rrdY27YFz+TM6ZaCMG8+b5u1XGLsSJ9RpUQzz4Nrv6O7wO
Lc6Eu89K5aJrASZ4tTDBLSXWdRYTZRaE1g0oTusjtEuzcq3IOmJ5tRLpBdmx7BLwBIFYn5jZJm/J
IYxRoXBccfk/eKE1zqfDwDfezbW8BDIdDZFzeGOkQYqZdJBxmw684cFsmhXSSX75GT68ZpCHMw+e
BGIxLsWY+NryPtedVzctHMI6We9E27ESEZHCBesmdHYyreZFYe2rD0jHkh54mHNAVc9tkQjawZfb
P7OBAwFJOJZEwlor9KvAPPmXYnvF1MLp93CaCFtlU+DAxuxDlniZfTZvR4Qp51RGHcSML9fCf2cV
QbW7qtJQ0oowZ3mpL4f77CLbkavgPV1ktC6H6C2pM7MHd9t7ONBsKCyyWTDpn/vaB3vIkEv+YNCh
M92aBOkzK8HLg58JoSg0bns2dNbcN7QxKX+QwGwvP29XZqpchK0NkAFAiJ3aB/J56c4yKqMahMs7
P5Oc2frFiGxGv3eKYdhlPqa0BmGnWH/jU/xi9Nlt474eZUTFPdnlblYn3cv8m4bYINf1vutJUawi
wpAnjzWYoRe5JlVBOjtczvxd06wIS2CZzkI9K9ssqN9QApjzlm9tHOZwUCXyPTOkeQsA7DWyuAGL
Ok9jSpj9c78Z+TVaXeXrdGdRjUqrtTZfcJckhkJNGgeq+UOp7JhsRp12ZufmlP3Jpqqkt9w2eq09
73l0l5vV2d7e37x18mFtJesSfBecLEyj8f4WquTeOpQ8wcwS+EZwzFXy8RMxQr2OHA6u9zhLIKGd
/8DKY9rghzJ/4hjm6mom7rWsqBMSLgK3jrEizVVwPIGfO0kRCRW8PQTw+O2t34iITRbmd07Kfgqf
g0SJwqk6UUPnjYfpvNC3OQ2MfPL2ZBvD2OYeqcLBp4MdkwnCy+Ee3mdcWx6n9TZnEUNpC0tex5f2
fV6H/IbxP2Xrk7buPlFBmy75wkv6M5Uagm5PGU3YM/O9yo43gKNqeHqODgigHfe7ljMg1MdelQk4
99ISiwlwBVWomxxn/F4EpOxhi1Ibyv4dL2da4lImiam01bdjTlc8nCda3I8lzqwBmpVPb9QRGGa2
+9Lh1BEKyNy5CID3/WYBR0EIG2q6GMHVi6ZG0HL4edhmGRL0kf54uFb0pONauzFPwcm1Lpd4tTB6
LIZXeEa+JTCgpIFElsWFpm5ZhJXVLnEFpgI9GT8UnlhNKIuKPM0SCj17Zy4vVdBy7S1Fa9Xq08kM
7D9zWiN7TVeTbcvDA4V8+BG8JcAfsHWjLt6MJOEl1+eMU1YHOW38MtqGo8KuFDlO1IlWv5GfImZY
YGVg6rVsF1dys0yrJB7nJdG4t76AaXIs9TfJuJD3gqghRaWuPwpJGJ+BHkkPK0WB0PAQRwWygpQe
yg1bUdh/w9HTgygrJujiM9gG8JfGABqIQMBBXBsDK8Xh7/bOiN6gx9dJ0imJyMF8F4hr7oskZfWf
m4G4+WaDRnfzFvKZeflv7s+2GxUBL0Jj5xKfNlq6eYuM8DOfOP27M+By8g6kgVktXayOz38O8w2y
tgLtURheAsxfmVA+BdwUXEIycGXZbCUuCKfQ0xjrMSMyYpVmaLE7RXAiVh0UafAjm3+1PkdsiK+F
7Xtz7Kmm3pU8wulFpWmG0vn4CtO36mkLPtL7/8wtPQETjZP1Ol6WbMfvsvC+8spLUBeRP2U6BC//
RqozODIwjB/V45xgRNRsDprbuAflqwNHdiUR9PXVi9FrHRg1K3Amx9N1DN1shJ7B8qMJwPn57N64
hfS+jdacflLobOcXXDpCmvuyJXLMzCLqMEFq0jkctR5O/NcvOzXuIJTyyTy2v0783nrbqStq9bwl
Q4a07MqpA36A/OsNvdQ9aAxyQS7BkGPII9m1kv0tBnP0as3HCx78KFL9+Po9PQPv99YdDLnP/Hme
v7cyL/tJWcwtAwVrDD2668Ark51vdvovYcQV+FnA5G6PK1IyeNYfdlnLsPcSChNP9EHUoGZwuSfY
Lv7l8l2QDkzJxm47yG/pBoVlAXjgcu7IDuFX21UfBRTtlMHBG22YtMJZsxL8aFKKMOruZRXdAy0d
HcgpQFUZgB6+THXsJ457YLu1XI1dC/hMn8Xacl6lVXZULIVHwYIApfxsvv/oUGNa4oilui5N/t/9
xJteGaMEj0mFuG96l5/ZMt+bnjzvso8za2CiGqlKFqksf6XrkElEU1jiIGCtroQegvhdKsAjgToW
iSEnir8RQjhxdX7iV8CZIBEtkDtoVEAgGn3ia9mk9/+UpqWBY+ExFtqB/3qIsxYn5YpduO86F3CQ
BxAPTuvyyKeoZzaAZJs2NEE6GiDu+t7S6cCagY50jCjGs2hoiXsBfrCKhLvxl/Irch86gEv2EPYd
t+gx6BWUJ5FM9nXYYBrHK8hOOuJlhR7zVxxc0p+aMJ3CM8+Io4d2g4jQMhj5DEeHQdk3FmkQBLc6
0R/mlsKjCEYzhXnojrmC5Uh4VuUDnr/rmOvTxleWHbjLA2ckKWt0zY1+D6KZpu2FGiF6k8uo1xYQ
+yr2q+ZOwu9Hp4t032iVi+mowcGp0TXLJdCkyOItLESfWziZowSGp6/n0rUeptRVDkxQmHjYsC0a
Ez2lxaW2N3VIxoFG5gIs4mZoi3HWR76UTD6xgxS1xqwg6jlbgI6h2oS03iIzX1s5dEtioMvqDTYC
kuwNjy4dLrqdLYhLZzszeBWyV7+jIYTotJ7eL04d3xs3nm9Uv63ggxQtN/4kdXe1wj7b+3pQ2rxr
MeogbTocX8VEAb0/Bk4Au4pdoB14xYnTJbpqj5gW9ocu5S0chRGK830+tmGITY+7y4KyMYo1hx76
QqD07HhyGEQ5dPBZXb8o4yU/qwoWeOcVYeWT0Meihvl9XxBupuRyGVbHYJHDmq2cnmbRpP6+ybTn
8nOXkRsoxFl0gmhC+VUDcnBPDh0F53Lsg/BHo42d6cB7hHJaehaqcGPh2mjHhA+Btk/u0GXnV4qX
yCOY1RAxhJoUepcBcxZiSm+Li1DRp4/G+6ba4qBSmgHe75Dyg5hlDUhHLBySxmARbl1AlwEO1ryh
87ckRRx3YJtBM0hDnOPI7VDc6kjyptJnDC5dCyR2P6rOuBOnEobEK/o3C64dlwkPnkDIX4VTDs+l
t6SqlGNinMWNQO2YEsr0p8kfTvDGL33xD0PPkgOspoZoY09fkfXSOqBTcsPSYmIZI+Hs6J+CCJAQ
duqXrOYhduE59Q/kh4b7ZUuGlpFG8NplQ/NVkew63vdgWa7gQnN6+So4G+bIsl79VEJe78N5Z4GC
O+ap0wBULgEsTptaVM8qpY0m/rSESJPR3MZpSQS+mHPnIBBMxsEU4CJTAsIdry0LEKt12IDCtCVt
JRiso4yoZ7PlkppgP0EkzYgSPPA95Kj/+EAVe3zoCbzl8vvOad+Tq/jg8AvropqK5XTxSO8yYF3g
kAWrjnNDgkl3wHd09RYX7UFesHdrBodlpH9uRcPj0EzaxVTfacHwOv2yvg7QFsoxlNTPqU6re7p1
NmlMd8yhdkdwxw4Ki6HsxWKubU+Hc0KllZIIHWtHTYFKuWWV8zpwkX8Nf7swZCiB93PuKddx4dvi
i1yYjrNtgyfKCI5wl5xAHWaonebnM/RI6Ypcym/M+5Lkuw1aoaUkx8IKMmTLKKpSeDNIUewFdPJy
e0N9PbZxCQdicAHmsPV+TY71qUk7/1lJnGtNjztktxkzqIABHxHa5Jh8KWF7EfcM9FqAy4V9Wza3
xSIR66vGDYk4sLl8ISAX0Mk6Zjh5oeni3jB2kP9EGKIJlVuNt/Ax8Xfb/Vk99+8HsNWHlyQu2L8z
wCYtoGkaxyjbUqow7WneanPEum/ar54ZcntNPUGval4OekRq8Bj9eALJdUX3J7CTwk2jZotMlQxP
WdaLYfzSTckUbr4f5KYhOtvh//3uHZfVOY6TB77Va7yKQeKKyLYbdy5LqqKarn/t1XgOuID1phzV
UFMhHZeDQsNO7kiz/i7eMpYFfOPNHOJz8RcLylt7Mlx+MOhcKYLMKdZnAXY1XY13HaKoJnKQvu73
lfuxWg0/4zr3pGdj7FVY1bpzK7easmszgJIxZ+iLPFgD0mnrhcMM69lpAL43B53avx5TcBBqaWbe
JwnE+mZ9cOb7dXiIS50hRWCF0ensArUJKdZmpfDfucGloihslOp3mWEShZ/dSBx2DXEuLBBteR9v
tsnE7Ex5hvYXhHSCSm3T4BrumSdpKrwqkqXkIZJC7anbcdMLvJH6UPstd7rYKYdmnzrA4ierAxSW
foDLZSD3IycBZvD5/6wDbgEr4tUFhJceOXfkj5iad7mAPxQN9UkiVaGqXBVfyWEptUzlbtO0ZVkM
V/nIiwmJdULr4hIUQ5QOrNbu+ORiOUs6BqBrBsByMSrjyQHlMszIdyrzR7tqx30x+OY/XIfWMKql
E3uiT5nruuBinj30dINQ190b5nn4tbP+vvXbpzKI0o4DX23l2iaunkcM5EbcSmG5DZGX0ueyc+lD
XtgKYVSgQnk6JXi+iv543MX6BjE1I4KfkP5vMJJkCF/EDh/qAWbQ9CdbEnByms1CAOQDWps04Edj
4iILzy8MTGWuug58WJHDn/Psolu/4VTGVmxaS98DLDmJF8M9BTAXgydhVqAW4VT3W5mdiX2Pb1eS
y2mzIQ0/y7HTjELvdo3OVi+fyTDb9KOUqI6l0Guj547K3c+z74M3xWClvGppffiBx0N6AI+ppeqd
emDwwZNI2heI8OcRJh4F0MLpiu212/X4Rl8oEeRDfG7zNN/+e+NRaot/03tpBXcvLjRpmSa77WjI
Wqk+0l8sSm6TrlKei5KVre7vUqtueV7y5/OD4UJhnWwb/YadrLpAD7OT9+f+ZxvUiDCEnT6HtUGr
a0pjLX1ATkIeOmRaNH0qUzRirZ6XF+npKhWgPlF0iMhRjThOfw58go1u/NdLUn1ojG9+bdMYLM/f
PQ9rMYrxtQaKS7BTCActuO2Uq5RXW8bCo5GkMlSLYbmKWONovTTWfu0XY9cdf8rhemS7P2OmidVz
kXyqhqwljF8cz4sHeP7YNmG7vTgrXhGH8r9RLX3HCF9e52r5rNN7ed1/LcLkjWCKYx/TSK9k2uA0
iarFHJj1T2wm07Vf0o1zbBtKv1eUKUO3wp82ou/OUhFQe6n5WI5328zpRqrFCT3SID94QMJapI+N
4Fwor9/LPmclb9wxWrTLqRTbaP5fP3SuJZf+rz7tZHpiYroBw5oqdtWwZgDqMXTwNN6MAs0y1sFW
pGzRGi6TJYFq+bTxYKJXwayoufwcS37e1oTURV7mtOUgRcMR6i+fd1VPcXb1snwOnRe4h6g84Aee
/Z5DqEh2bJSdU9lcxwETu77mEuPx2hAwpuD4DpkCI4diXugYfv6LA6zcsh65eGn6xFgWxfGZ7PPC
KnkQ2yX+AzWYNIPsP2yQTqLqD+ovAulXVF8deVDp0+4XyCVVcR+BBKx3RKkro0DOHk8dcJ1j52PG
fyYpZmMmYDZ0JSBXNd1gkSr4toZH9HaFwVZZvJpryY+3YDE/Iqvy1ZnaVHLkCdERk6WnL0wxUZSs
UW/Y8Hbgig3rIlp4NX/DFsLSFSo2fvvVu5G+DhkCsdlGdw39Usw7UomHPWYJBnB8maaZyXwACKTo
OV7Dh01T/dhy2iLNdHfVWPn1fsJRonV7JHYYdLbzuMAxow/EUUqjgV8IWo7Z/1aXdupES2F5GBOo
tPysuyI6XEgWJ3tzMAB5/0FqXRr9HbAzW0MajUp64eeWUfu/8J6f2MvmT9zUP37mxcmkHodTAR6B
pXzS02ut2iukY6A6wlvbDft0qqOb9KdJctlcyGbO3wsKrM7Yo9gVmV4YiUKyR2ajcc31WOrFDHTA
pRJDe6fNDMJAjJskKSL4BpSmch29OLlJSYsFb5wudMVj5yiZwtQj6UET6SanZLvVZ3Tdl+W+WwJF
MLtTTsC/5RnVrGzyVwDqLA0tRW72R6k0oXpeyg2366+PVrg3jVc2rnxO94YqU5cLBnUz+qtnfaoi
6hcuY0AbF5/Nw7xzCVueHd7Xmr931tFrZOi3wenuiXfoQPKk8+ljg4FAaZN6xVzz+G9u/zL+qOZd
Xno4+V9jk8acp1gLvxcxS8MFy0d5uJED1z+C8WWZg8HAaAqipC6YUDYGYFB6yiWBaqhipzC6BYCG
01FfwUiPYfovTDPrH0MIVpsS+nKoGuieOZ20suhmXajydfS8tU8l16d2YnjZ9JiXyDsEZ9RbmTcL
Pp30+sHdBjcAI2/DkvcG6JL0I54K2ejX4W4YgJAti2qd948FT0kVzOrfiapqa3OM+0v5Ap6skrOt
xpXbu5VRRg5UN2ahgq4CThOh7yUKmCb25aiv9wdXKEvoNfUIMNgn+zOJeJq6yBc0qc/XSy+RcTam
ca4bFwATlf/xMX++pL7/2YgizL6uAe8KHo8h/9mXi9leQ8ZOfgg+7ZKDiXhp5pk0pb8QMx9icFG+
paFdJ8miLzX1itfVdjbAB9ZE+J6q9e/xfhjFYAhCy8up1XEHFbqss0UtuyxixAQf1/uNCREcKtNK
RyMOBil8CjTqkdFRHmBlyKqV4RarCNEn+14L47N0NEecLmHexwlBCqF1Azd1J5F//n6yJ5X+XxY+
EMMzDzEGkciEruDuE6Q7pMDr0Q1oIAV4SC73sBN5k0mIbDcmPxiLOzofHd6X4P0lwyxdY9RsHVnN
ttYHYql+zKJoA5s5w5zUYGoqipI3Mn6SAMrTpWQTMfvS+olEWfhF9CLxvhOzB/B0BLCzj0Ell1jh
U47J25ija/b4dNz6Li+SasTIVVEG61rET6mNib/wWgQyROdvW4CcynQPeo2oDvxPR3gh2ym4CGHG
tWldsg508HVxp1+gQWMAFsIJ3nxT8yDUywJ3KWeyuCMItWHcOXSTbViCZ6mzodcDm1m8f7BxLSSt
eqMACbn5ZUxCraid6mYWkOjEgkoooMqOBrH9m+XR9Jssx7EV2YxhsI5oWiMX32FA+QlzpaiFMDjR
x4pf56692JaKKyC8YP8I4po6/7xlJTK6hR/2CojKyEYHoXwpze922Yrid0NAFC6tGXfr2JHq0Hrt
do+HbvZz6FZosACqporOImgBEwHu6JWfp8jf/WNxwNt71IPi6yCKHJ0P1zq9O8MLB0rA4IrUTB2o
nNuaNU4nP21s5lqR4Lui9UvNI5hB98yk/Zn9Gjo8wGna6OJbQPgUi5uaUbNKY+/6NYRbAojtcPxs
jB1JMxe4HfCP1VN8dfs8SyYnuMOyrZzmNjbF70/gfimMBvDcGFAvfXEK/B9/ciiUGPRWybInKsCX
dFmSUz5xax/4BwjOEiGmSoizYrzA2kT7ZyBl5z7PUrlehJEoz0R5MTbgrdk1gavwuKkddUtWyuN5
jeBvjFtY8Wi5TpKt0Jl0fVbc/AgtuOOk0tGm10btacnY3FS1McYc7rax2MAc/sJ85FLSv/FvZcc6
StCJEtNuPUXLNkjc47IW3CprU/aSB18clMEPokJznnGhG1mR8LAZ8mipj4QvQj6b7ukjx1SfeMgo
84qZeLyEYSR+VVlb/fveXeEOlldCFSMcuDk+jxD6c4ZJuWLiFvPfL9H4Jmd8uhsq4pzT2QepHC4E
X85lPrcSV7BHSlcPPRAr33j0QmKXQQt9IL7GelfMAMBjF6I9iLGra1Tiz1SVtdVGnHHoN1P+UMv5
dx2zN90BEPCb8Lqo/QZO89DXGyoIHoeITsBGqbrpj4Tkga8rVIIJH4vo9kd217eiLppu86qwaa3z
eo4BdCZ+G66N4wmJJ06Zo8Q2uvHGKn6ukAw0fTEZBJR2suVonKll4LhaaGDf7tVsqcQNaSNwY4nM
82ogMqkqZ1d2HKra5L4yYFV13Z0x+LcjZCRc2KA75bO08Q3IoHdDMKSc4VaVVAS2/+3BpochQF5i
iiQnz+maUXh+xnstWLV0NynylcqWn0j8futxzIgM7No372+TnjdtvYiOzWZ5SrEu8orllJixp4WF
VC9FRdjQl4E3i0Oc4I0EdQ1dct+yjK2GZJkR+zOX10DdtBuIP0bIyEzmvEfbymDRuyyJPfiI7HJD
OPR7IZGMSOHiuXUyTwnJUGYA/pvqa7OojBHBSrdJs0E8g7U8pLszL5xYx1CLQvfMVuJCAfxg9ycY
OaKDPGqmgUy4zH5cxjkRm6R0LIhvOl/bfBtp8YY/8gdjugreGnDIRvxzi4uN7E4fN8x/SZzEbkO9
KG7NnZSWSRWNIilkm5beZvjUtkstpss2668VJ59uhn+gBzqWlfe2YHPvoz/aoaX9g38WbTpz4ZSl
81ICWNWpUloBJ6GXQe7mTWg2rvpjs71Ds6vgtsQWDt2f5PB6LpE1MVQbbrgOcF/KiSzclnbKAE1d
Pw1RpIlYm1G+7zDabrr6TDFoRghFVVj6+keeW3xGwOqDILV37JGQi6H1E/TLYBf8CzNa3pZeB244
oUzlw7rSEEG7LAqNzj8qknf2opMf6HN9La/kP+4AKCmCqge9mnf9ajMhAf8jQKdXPaCDHP4CmM23
tzZWhRpMhgfJLdcnepASrlQ3RTBlDi5tXmHBtKfZ33qFS8y0vdEhzd1DdOm9QXEtd0Y9TBzoeLXg
YQJVN6PdjgeYPFrbirqHtA3eKC+PsGydS9PCvTobEFJ+IKa4PiRRG/Dckd6L8nBD9Jti1UvQlKOm
C4u5c5a9P1s4yABHlNX4fb0pLxFXly650W77whKXYe99gQVM2Wl6Bp7bFHMDStDC8RtCdUUEPrrO
EcVR5YmSBYUKs4tyVnh2O4w7GzqjBL8iK9WoD4cVftraND62W3pnwyYT0JhgLBMm2jc/K3O2Wa0b
vPEaFRf7A/9y6Jfo/oJPS2krx732Bfxms61G8Hk/C+WtsB5Tfp1clM3kHs8hlpF4XpV/0wpHK9Zz
PgwPnTBa+f8IME0aUCk6UwQxKO6ZAFt6xGIir1Y9TpCHO5LzoQUZshHmYvtuW7Jj8vCbUAd8TFFf
CCtfe94lovf5HuCfmIjppbyP1FGQ1aC5Q2rVKFg/3syg6wjpJoeW+Lj7gg2K/XYGzwRe5F3Itsk9
pIxBfLYwdCMkMYTWgBYj69ZMxysvJh1Xyp30u1cld9rVhuPrjUkB8cieIkLiB/Vw3zpJ8YfCjDjz
JW8AduchIDieASh+2CcIFEB7TLd0R62IqB7tyCIfNOWrc+lI3YhpthUz50bg+8ERWIwFnropm2Qy
CF/op5Lt8HoxBd1wpS5j/3qNtZeMAtuph/zTGHsWwOCoHIorgd7EsSykOPjFRU0UOQ2ljLi4tOqn
HryFcjMQY8jy6B/3Hbe9a4M1zhimCYTbA5Rh4sLSrJjZTnrGZLgYpYfspt80+iSLnuDyvkaxJ0fx
axKaTPeA3H7u6aNHsSNy/ZMdaD9jInJ9pP/3UQUg2653zs8trffXj4DkzWqt4bq/p2GxlycUWw+j
5io2lsncv6UPAYoJwj9P2YXnTng0ZJH7Twv6YrOLr7OdDb05V1KaZExodPt518Ta6/TOIrxqfdUR
omdgA9h+MRLo7IcFoLo9hMVX+O3kr34LW5orxqiG82Rbp/I9lwfT1GMXZeUWMf1T9D7KJZDmku6C
NXG0ZW8/NDXjD0UAzD7af2vK8Il9LUTldahL6iOVhDaShxbcXKBJ2sRjQEgGk20kU6Uq2gH8Rl7F
yL+g1Bq5DN74ZpQEJBsDtVauovg3r7wA0cSsWQ+SrlQJtXb14AXeRtART7D7BZLX7aqJiA166WHQ
curFvcJjL9qp7kJ1sojE1HYzp/dcFupSo0rirp3guuePoM2DrO/I2Rt4aaxsIM7CR5HnLJGfgXR7
4iUFUuwcLNy7WdqCHGilY+P/1dUwcsXB45CZGI8UnQ4ZgdE6asGBcwJ0t60NWuPftGLNgaN2wISz
Ksd8c479v8inKi5VAuugZsJdt6wFwC3H5pRfS+8NDmvDej+zxkPFOSj/yEFJ6YufK8t/OdZVKKQa
w1s3cMl3ZEhOtDAo3dJ21V4mrO5hg5qJTqU0O/7qP+e9XDSxY6B+aebIUcEtTxg6RgiKSQV5NIA2
5BdiPGmZU4doCZ6ekhzeXTLC4kKl4gaBQJAg6kLwTGKVgyYU53G9jmtleswT9YOD2rf7YCAcMetE
IOkf/11xeiyxMbvgm9E6QYG9t5TrFBytNkedBhIcEYOm0WO6rNfYShFiw+uqvE55ZggLuKfvj7V6
9D0vK20PYGmyEyVhQFKgA7FWsfXRsbyaec2nYShE0mM0XkynCs61FcY8wgSde0rxXY3lwbhZwyNu
g1U4AhA3p3tBZ2Rr3VKgCvBb9uH6fG2svNSUanV3eKeBm8ypmEp+FOzzFfYrh/7YOsfCXRjB/z6V
V4ONjgafjOKgOeBhk3MpqIWIJB1zrCyB0lCj30gP3LubP+7GoDv50L0d5YwcLrGColbPAtBhBhNJ
3zyTir3sSXhAU1bczxMTtOLkPGlv5RAa2SBxZQWZvH8KjxalYnpbtcGKH8mMFaOL1GW2RoW4Pos6
u+epQokSmpov33iRC08GBZjYjO2zLizEd8atBJOSF9eHKxlXWAJrMZnd/L5QEF7l2SCYecG2oRvb
9T4b9sdKfTfJepZnGPajzpF6KciF7c9QVHfGSwd5O32IidZ/g7XNRTwTzuAto6WwZ7yDEHBr68eX
/2BpZtZ/7z0miL+p+0x3ZDCgnuVbTg2G+TSjhACUA8QdyxD4GUJ01jtidrgpIcNnFK31mZmup264
UM7/62sEiwKKn4kWnc/vakpdBT5ZX71UzUCgj+mMlxGnSlw7TvfR3/c47zPRZw5FlPdTbdp9iSjf
2nQy1dJ8cfqVP86PVB+72/IU5R19J0u4sUc2h832F4lYbCtBOTENfmS3fpnco/0UrA57KVj0e9nf
uGWC4o8i7Z9mqDaFsO+UZ+C6HhvzG+BsvOqbaEdv7UkkjUaiEUXDGe9r2P90TtBU7PVUZc2DgmsB
AtjPaUyGW1T9QiNInVKBGHTWS4VSIv3Ozwgrhiz5Ws91dsqnjcUl7DiBmJvS6pXhzPah5Idk+c2c
QzYCsvku+l8Egu4FVsy7EFIXR8LgOXRJSR9xcEBS7TpgFMtLTC9mAFvNdxKE4DOXkMRbXGj//LQ0
C8jS6xSZLfdNoROQBJpdLTVCP6r95uzsk/K3DrtGYYLoNnmjs1VL9FhN9+yKTs/dlNJY/0ef7X4A
BFgkH/cmzFLhtCtiv5uoNsZDp6ib6FgNH8H+I4mWuIKPnC/aSy3dCl01w1mQIhMOJrifyHC+gYU2
otFzBpyppciIPqIMbQXg/Pp8DK6KUucxtvz9K/1BscOslTkal04jUa/x/aeIk7BXZeJ0CnerGCtY
emt8Wn5VyBoS1YXovnKbjraXXDyXFaM66DsimOAaK7xJa6N833sFoQQTWyog2BR4ZUEhKs70jzEX
l5WDF8ClylxE9riVVMPpMrdmtHBftgFORWir2AlM6ngWMoq6uwPcCwpbTWFieOhSXEgaggSuokXd
vVB6CsMm28J68l5YQNlXphpLddpFDUkh6J0juVz3ndkva+oou57M0EDzuitsNmJEIPIJ2oSNqqO8
YtJtfgetI2oWojDF6++DAMOBDR7a7GrEg/oueQdg2+284YBMfW7EgCAh7t8RVMBk2Mclnz3XoymW
I+8tSbmM/EUV+0aRioCMwcZbmC9Dbr86o2GiEk5AXKEzFQY3Jz67VW3FKWa022jA/s+wRvMCs8qb
CwCMwCwPFmQPRLHV42kYX9JbrvaDGSdiadZJPO3Oh24D3lUTDefLQKyjikk0ibxl7+A37DZcZkSR
Jn8ATRm7ciRZh2SaOVJFeE9OKb+3q6dSenPzKlQ+C/ofuuc2UwSnZYRLLYDFxLvf9AN6Pyqx7o2M
tI5w6SQVtgv+QSSWQT4vQ3fwwFfRFiwZ6/kxZ40veVaLwG5jqIJ9KtdDSGkuANb00/oUewm2rKZU
A9aleSVxArji3b86Av2eWHr13BfB7JXzj1b6YPgd9eVkv4+j78wmWOGV1U68a0ZzlSVAqCP3RpsZ
FWiaPpoO70ByQAiV8kxg2pqLP4Ml6nNcW9TKZ8RfmYS1IdOX6p5QiqUnSJXehOcjwEQiB7mh0uhn
Wnas3ua5HL6PFVevB0xyeTfXo8gBV+A5dN9OjcXYsq8T/rxJOgaGecplLIthAAYq0otUBNmm3DEH
nqvuWss9K0MLHSrviCT4DOgBC4JhaJm6gqFOCBX9bIRfexiYulBMXHLx4uT8SbdRYKkaDQcj245s
WOqQhGl034XpiUiud8nNwSToaF+RPDSisO1qgohY9NGeKslG+oWdA3oVYeM7T4nYZCCJ1D3BkLEs
ntA9iWDxLfhpKG6LG56DcvliAkvRovpJ124yKKilPb5GCKRuZRuCpndDVb1hO6iQRLRzOP8iIjo1
B4UHTLWhYNj4IHr6r8BuNyzG/V5L3uXaLURwnDO241DxiNKr3pD+TMx8V9ZrdCgrJIXzDgyyarSY
UavXKQyC8fzy+zPg8bd5pTqKHYRb2d9oYsyo7HDvjPVq1rz2aGZHM0yj7KGJezUgQZokPxvtGv+A
ynp9B3XJ4pZSDN1eVf3VkvgG1nlWRBiuekNGGpwM9dKdeoQ4I0O6ks0dnGxl5yHKlNdLapGQCfRm
uPtJ6k9LR3lf4xjj6361WCV6+612eWKMuK+yzGi+LVASNu4YpxXLXPwD4tVQ9qMADSeYy8fK8qF0
XV3QRbJOla3HblDExe7NmvJMJjsFTaqriTxUnUPP+XQVbmD3yr9G9zokoHfe2vDmqnIpB2L9ONQx
KdNzOUYBb9pg2v6+zpSo3UX15j72OsBn0giKCO6S3+N88bZ/DBoiCyJuAYGHqLFyU8/z/RNkbSD1
4RTTDjJ0ZtQmbuQBd6uEVu3F+qDpfvih9wwz3TxSoFnoJcz1brnFNPvnN60K8/MEHA1+8/5SvZXF
HWvOV8FEjk0Wq/M0vWZ7c7dA/keKASVcr4rfyPlN4IY0LUCDF/kNti5Z9PGRsurryUhTFyiAumLY
PPxg+EM8iRh3/K1BxzZagbJQFDK6M9TMUDx8arRmnJC5kkYPOtIAnStKT6itreCTwaYS7Ofnb85N
nGSQveGMfJyjJEN2jIVJ9Td9J1n8oTodcMdebWfKXns5bwnH0lqs2K/WdHd4HYpqI9FHM157mB3J
dtu/UW7N0OAOs3CCunqfQNLggFS0DIgK6SakyrCnVJUpbs4nGgUPXQBLrOkhaH8W59b91C6ws8Uy
8mFhBRrJI5YttUN9JczH2MfYdozBW5fbZN7VVLZbT5jMvHS8ARL6mO446EWvj7fW9HJIxKe49PEm
zNGFuZYcW20uJ8UWGx5AASUIQYW/KqZDutB7VeiRRI5E4Bz9HruttZGK85sORIqAkm9uwIx0fweX
0GQrc9BJsJvMom2StsV4CioT85YuBEmJe1RsNYTwjhggMbhugoma+l4Zl3YQj5Ff/cTLCaMvkIID
gv65OIRZ3ztM4NvQDS/XY3MNlk7J/NTTBr1WVG8rMEESVMWxt3Kbb6qKnRzaapdvJrSaLZTWMRvJ
OkUO65KY1dGcAuowh/LHRA3/TOcM7Ni8z8uy7KAX5I1RWFogLaVp4kIZD8MBwzWsZzv7FLnKNOcC
fNG0boMsbhX6VbtxZua+19idGvy0dAQCR2x3sZ/V+SC6t/SkaCskOQJx59yPZ58pZpMZNf4LHmCC
iOkslW/ml7flduLrADlmZYEYdu2UN5lX1BHLcKXgdOiv+EqReRKAY6lhHbhpeee+maU9RMDgBlRd
iHOvdQjPcjLrIReYKzQ1zQnIdyY+AQtgbN2D0YHdXheWB3ooZ7+gZ3G2YOO2+xc9O4apCQdT6BHj
kebQDRRntYIvdWLTjjRv0Ry8EornxZdV5XkSbXcKBMMAfu+ZxWTLWqJjAvkIVxTtx85cX3xL6JrK
QSFxwj1SY14Q5/xcbruyrReIWY3HawKxxZUSVMjS0/I0FtpVjuZOq1hvYAZeHJ0u8Osy+nZucyYe
gwdBZvMlMYR70PNd5TLRlfs5YXQcmeEvmdmHUWVCVMZ/d45g3OE51v8k7an9doolOemAYZfO/0sy
j9wwmSvcseGY3jZFy0w8561/kfP5h6hhQfzB9xImx00x1+xn1c+xkspaA/vSCLHhAjk7tt7ofAON
wYObSXbdG0Tx/Uhb5Ih1Jq+3oLgqoKHLNlhy1EGtQpSoXgMlC/nbh7wXV+KvSVBkLPxms+2VGcYe
DbCmBpZ4hDSOy88tOlJKRHlYc7AovA65fpBgniSvA/STcEMzZSgNj1uxBkwx/+OrcBSRefWUokV0
Rtw7a3ZW5nlsqRpz42G4PgmbN904qxOlrsIhLvqMzEm0ZqTpVn6p8FW2O4dQ6uX7K4EX1meR+J6A
8v2NMg2l7kXLRKYb9VOojoBJM6aGG9ro85fDNkCIuiCcdkAKJy27G5Nb0eJfQp57lvUkGiIoWK3Y
xqxG3oaxTa7oargG3vLXolMHBNrgarkREeoSKeTyvcxaes48lkZqE+lTU30wK5eUzQwcb7B68Ub8
TfBLEaWP1cv2WN0f1ahLTalnPdBzwzD8al66kMUtWjIBxSLwKqk84kkK7DaciSzohW2EsEuWxOrc
UHUnMWAMt6Letf4Ed10YoC7zY6wKSGU1VMeWTmH8FS6UXC+fLTBDCQmccmmpoFjTWQ8Lq6wLGg5V
lEku4OwFUzO2AUG3T2A9KnKBdNoaCsGs4Iu2UUzmxvD5Ej2rbd4y87DnlsZDrfb4wu1Nnrxu+yWQ
zrqNc1aXf50FWySNdRylzS1vZUH2gAxOqsLVgBZiguUcLpFmwQXIIU5mQDRTQlCYdZ7MqbFyeugw
PmULw6uc90RGcmRUI4jShaYLfziJZBXGh43HXw76kecael7V10BJb90kTAWwGxqLETzZOVYbGHdx
l25uOOcYTm3d9uJE3E/fxGZFOKZQ/uFBmwrIJU+BwTSJEU7NUDDBUHkAnKgYC882oV7be5Q/azmI
yncht7n7/EcKn/dZ+6mE43Vshvdykh5DAFX+GNBRx/BmOgnU6yaJAx1pGOlsrdvImI6Ws0uqxDmx
hVOLoR9qDvr57ugQPrzujc7/JLU2kQ255+UCrdN9a9PdR3nVOm469ot9acKGKP0y55H6KPyHKHCm
rydmn3JAyy+m1ydTIiSlGMftwnkaJytwz1c6ScNxPcP+L+MN4pjScxTs7xjwK+alYgs+/v7FUV7r
hbHFh3mEByv5b4OZfNdI2Zdrkq7yEg/Z/ayYF9O/n9IJFZ5HX7eUIFDm9UkkeFrlTKKSXTjQdxXZ
qAD4K1t2Y88A9H60A6psvMZMNPsAdbKQlFv+JGFC0UHvx/IYox8y76utRmOS6sp/Y9FaviRhfzXF
w/bHiO2yvtP4Cw6nvhIXW75hNSHMzUrsrmtnjHq6R3C7mxj659pptu4MX5nF8mdtRfJlBv6LhAnd
Qois7/fxiJUCiiYGIggYNv7wKnMTbtCAnPGHNt7E73AiRKmOMGi2u5kDcoahv1v/P9kv1vmGF6n+
bmMYhkNI+vGwT/Q2FYuKWAAUqbHvdq+HOIl+BLpbWRsex2Xp9VeKbOvZVv+pwk7VnghIKZ8qGjdX
YzcxzOpRn/ekxyL5ixWbkDZ8ljdbavgFriRR2lV1bPUgeU2zoRmJGURN7fRLkV35mJ0XpP9BFw0a
1DR1ari5Cmiu9xu7W7o/2ltUlt4Hi1cLb8EO3V87ddVLeo1VwGKaZEmdm3qLF3p+oYobsvUKK7Of
QM9Vp+0ps/SXM2HyoExzS8sP9kOk5dP2ljfb54Tn0vHl2Ag59v7Z+fSZCDaxIBZEagcRFa9TMDWS
arRplIH0CXposEnNluRidnfJty4CJ2+kueB2jHEFrcuRpK/zyGwftJEID1mijKMEDfzDezxzUhzJ
5dcim4aHgZMF4NUj4y/e6FZQuXmoMdQ34K47d1OeHhOaQ2Xp0YYLR/HIZuNEn+pgu26jYa9LuEgv
qFLjNtjgLTJ4ogUYH8tTlXrsXaNVHJrUzqyS9g9Tr2dNYZ3DcdMiFuWC63i3bHlWATvbelwqzupp
Xe3io6B+PmTe3CA2M7efbijBGotxFB+X+WhSqwoUGpoFyYYk9EJlr4TuzUZ9njIDoqt4VlK+sMNX
ivlpvuA4EBIcca7MIcmh1Bf7+klwHfaCO4S9BgQSMB1FZweRPCQmlEiv3Di2pGsPJ7mSRvcf9gwa
YXkSzYwW48O+6vFZeS23D/az/PKrzlioQMtVUlA9tgTNlx4wITiRNvpMgjtxcWLoVi9yLyHmX/lF
TnxhRVAMZ5tCyF/vgMYS78YzD7bwxatYEv/wksjFgxvkzF4oErnuzFDjKBJxXuQM99KOFoK5HbPH
c1xXmucDX8h64HjoI+T9VgMrWPlcHQjrJKZKCnw0z5H4lLhJ0f0xpxoy4kRkFNdL3YnksZ7CiOlB
ffFe357NAPkEdxllzNHV0XbobszIyyh9K9s+XhPbbWURPGACpKed5S5ibiv17WoOYPAEI3tu9no9
APnCBwzC62MCz4GlVOHYzx8kehEyxh9rvRJxNRGDQiZpfQHHtG0LLMFyIxVPzvQPnjduEwFHpMkY
ggMplfK32oSvpC2LEsgQLQXDSy7KtBJaY/xiZBW6q9uANUvUUjityxrQqKKOZritBh0WDHoFrdvJ
8J/v/qQtn1osf7oKNqUw67UZyLpPYDCPWzN+rX//50mV3RbCk3fGRyVqN0xtUVeNOz+xG1A3hAlp
CbeKme7z3FvC3wuYvyRyD8Q2JQyxLSNBY3RX8i3n1tKnOdbFPWFYHIdbxVS2AFASm17PoIIGIsid
35kG8SrM5y59Qy7vAxwX06om9RuffzdLju8QAG+bMEWK1nzODRHNzgXteRmk8gtBrb8KTENJCaHA
WiV8Y0MLj+IlyjoTEP9l+zs5TBaidaNYd2+a0yLzNzON7wL0GbVgPsoX7qk/wyDPS9lQ4F8AysMT
8HDrMtDDOszS4Pr44eT9B1deJJ4hNwLA0C7hWHZyUKnFSfjj/R9vpnYwV8qynvEa6OjObn3pTyrp
Nzfhg/jMMob92GtuDGTMs8BoNV8fzug1W42TZFsF9OWoGZ8N3aVZkL90hSB95yaQEkrR+PZm7KQp
XaExoNs+QjS+PZFtA75ewRi/rVCyeZZUs8qOeqR8vzxId1PUvmZfqs529+qwZiO3HkOBMDjWX/jV
dWhUBZo3EAKxbA611tCw/eA6w4oAuZtIMJkfupgzQy1ZBy45mAvaDUMn/VVrtvYvx863MfKxMRj1
MeReGm+fomZ/PtSv6WmrMldLKtUKUf7wXvDE5g/LzWSL/wTLUXYciXSlA+yokHBFwhGYsL97700J
MNKAXSRiALsnw8RK0aLsXz+tt+RP0RdGQL0HuVR6PRToK5i6TcPEYcPhz+QptcH7wblZFNw83pVm
XJ/WGPqMiepJfhNqxTxwTUzhG7ML1nnHGiYeGBAxv8aQrMY7zgql/9l79B/uqvBpB0PwOmX4X0LR
7/bStvEqBKpaGBha7lhQd1DttiW0AmV/YC+KxKUduvLZRE5p+XmyPYiqzmgJjyTUEhA2APh5ffRd
xermTdeWCZrfnbqJuY3UbjKzrHkuWB1oKPA7rGXRekMJwm5Xbw/wF0E8X4sBbgp8djDAOysZdqbI
du67nHCcLDRJJbc/TH48Gn44D1YuY8m4mOF7hEPlojD4kWwyAevFDAo2TekgsyYMJHPH8v0AN1lm
OU0wEa6f6xm46QiZir27uycIgw8cWzvEbtzS4m+8yUBLpvbimIgD8FS8mVM+xyGViGXMNby3A819
g7bLGjLdhpArXpIc9NhLPGsah6IwW31SY9Zw7mqjjHGogTw8HnX1+a2y/N73LvmEk3Ufys60kRdc
H+4Vk28BlJPq9nDCfl5ConU8d1i2sIYVSaAFmSrd+tuvRwhSGvamXC4SGL/VWZvpgSKFwk4NA7yM
YBY/s1OZzf9HvH774kZjqG8zG9Z0dkcVd2D2k1r7HRTPwK/zGIncOwnGdBp10j/Bg2DgwPtrGdC8
CauoSVTJbHUuSLJQXBZ11Sau1mk7lwujQIFR0ZT29TDAf+YYisFnNk1pnh7I3KuabH80a8XeKBJC
5MUR/2cqcfieisX7Gn3TuykqqqcuvIvwwfOUc/4dZdHAwROfjOWgtOwMf+hWfiqeBBmVyHoEmvNr
oTh9YCHPKX+yIYDkAt0EL2V+38PR3czsVv/oWWgQYTth/ShZ9YM5PnalVs7K+iwCe7vmgT6Zcbxa
uTFjOA46lvNuCiZT/m6C81pCuP97sMfknXGOHRaSC8wnrIMjBWuCeTWLJj39AhPmpkGSWmv2BN0s
FH3fjtktPLNKTzWm359CpEz0R4bzAFziwT4WaEvRJbei2EkrdKHNkbMdxTyvsJDMH9R4riBXqoks
H6V1w7ziw+6oI4e1arpXBOW8+g8TYnEXy+oowI5G1wrtB61Uwra4rlSIh2Dk3ZvZxgjANpRhbdDF
D+9oQry+6Wsh1N1tw0g07eCwYHpc+E+oyAmcheSSO+Ro9vLKZYufkdTXCUZgwtc2WsO82E8IsSV7
cqO3aip/MFhGsdIRUjXQqSL12S7tiIRq/RqXGFvv1Y5zTUYhRsW/LdcjGthHZpBfOHCJ3KJLbeSl
Lk8cVO85bAdKXo6w66N03yrWPMxn2UgR88m9yyrHbPpnCt7S8ED5ZtnOc3DB9cXAq6+iS2adLa0t
UP9YHdfifeaexVcohnMABokDMTkb4mHiIImCSZYrigyKsbTwb18qT0vpumLOSsOU5LL0BA4iwuHM
VtA3C3139ZFulZtLaORPxKNyvof7IxXS28OnvhsN5XQYS3urUuMvM2Vrhe0O+MqBH00pGRWUAdyQ
GRAsL+FSCC2ZnXI9GAhisqhdryn8ZXVUgCkiH89Hy7A/1EMAjYtJbjKf/Qpzx6df+IQFOik2ebzo
XroQlmeolKeSkPqQxf2zR88/m4UQZ9ftXHbsf1HB/rKx/zjt8Z3MKm4s4qu6zhsOJwRbW1ZquCPN
+1Q2KIfVpvYjyxJo8rmHCp9cjk9zyxNZJLWAEokvCOGFkReMs6U+y45lX4BWYiT6tC3RheKoPi8c
vhPpzOhBQ2W9ktPDz+rR3jQ885rYFAuDI1lZYPcUf5a0oJzTH7NnuEHO2wVVxZ0BMmwN2U8qVpnZ
787DIXJiehUlqp+2R5Mqt6cg1DRxzIti7hrrFsmnOyoDZzpRxoGga0GSHSJ1dUTK7Bmf5jP9LT66
/zJQSJ/OBJ9gss+QppV3EF5JFSTal2BaSN4IFo2aY8uR7yoKYRWYy8qVMu9POSTg8XSwLS5yPmlY
3DNsKJlZdkaOeLKSV999XMvWtGTLYCFrPfyAGQrjU/8sq2Vb9f45BmwRlZk8T4yj215CmsmH7ojE
DorNcJ391hJ033NtAknl8TbMOIcAO4I6whfxh1iJTj4g5D9j3Mtl9FDAwLeCW5vZJaIf+8IIySM9
WkyiTLPBxk04L8h7pvwYq6Vu7uKg3KcjQxMuIi37GQDp3omErdkw0rGUnP2xN1aqS5i8vX3mc2iy
gUIHNFqtrHOJa/2dg4M7JRsNJoD4zqlnWF6JWwwlj6h7h27Svt5QqjHQSbYyDf+lh2PcM5daljZ7
86kRpo3o0D3tWPpKSrK/TTThwS4SdYJe530xtlKTBzjE/z3iLiWH/5BNhzRhuGFwm/TDnlUHesUH
gohmUNSJzpnzCQD65fYd5jog0OgPIQRQ/SYfdz4k7la9uixvpjelglTtWAjSSS3jP8nqv9jcyeYr
s99mbwH3VTBgA+g7uVoPb+kWaU5gkZfwPc/h5kLR04IANYGj3DFKUJUXTK3d5VH+xARDaoDLLrVn
KKKbHOfPrPvS6QWxiw43okNzpkClXnG1l3o/0r3DULDRDSQJbutwpg2acb3fXmzF0383QWc9QgD/
c0Kx8Krj2tr4E7H96INSvtIuJO00BJdud9cxmThvmApEIikp30h4jCA5W87GyrJe5c8JQ9WDnEFn
MZNUAX7p1ISHlDexD5vtprySv36ldvpVjlLvafLqczK2b+WvDW69SOn8Do4659Z+6efBDE4q4QNx
C4uRglB9c2Vr4n/rPxf3Nr4+BcPl60sWu0512wUsRhQ9FjdTIl6R26x27zZn1XmG/pCF/Ioovfn9
x6BirSlJo1I6VuG3EG9yFJVYCYFVM+aneca6+jfwZDguCPYWYApnuDzHk6DS5YbGkvTBbxpMDKuC
C5AWksbJc7IjycG3DTTrO+VgbKo4ObhuQSFbaRQ1Z4pyUDsoHwPwjv6XawZH+7Sm62TnkMSkksrI
Cx9gW45XcSTtEp4NQzyKTurCgTeW6+CFDAGQSfgCUxsWKjdckpuzowj0LJv3htgzQgNEIdTYdfma
4HSmA8LHYfFKVFnZwURafPhZShIEba4PtV/JK2Jo0wcs13wZoDzVRG/Pc3CWDaA2CmQTnoaizD7V
WHHGDOI9Hg16GAi5gNTh8+HyzLYNn2YtuYE2lk0buMX/+qYroS/UwtNsNYwT7IqzyKsAnuEwevOM
eCSc5XlhZtyQ2YZDQrllSi7Y9ytFzUUD320DLeZ49n46uBe/RVd37JIqppKQyAvtpu+JItaz2mHO
fh37licQPPC1lN1b7pT/orBz0iZDT/fYXKPO87NecH9YJtSMSKpbx9ZdzLR168vTZqabisq1kImU
oUjNAzA4F9/OXEI+Dq6eYL036PLirCGsbdIzwHF0NxbBvXHSQOLLj2RjYVxfBw6ucymcLZ3W4+8y
Ye/N0lcslgDKBhSaqTYP/0PkWx0qRTqvmyRw7csD++CFaKHZqTqPdqLXY37CoNxSph2H6v0AiZn9
CBPCwWx+l/Cs9glL6LkBsQG4zwAmIeCWTKyGkAcUyaEiVjdi9HwxZRMUUVEmdDyIXFPzkPP6cMOw
yrJbs+AIRpSBTIgAyVD0HrS/sXGtqcRgfYyrBs9UUcPx8yR8xV0kp8RCbZSqe+FqsAVFmkJnKG7z
kWjosOnyapRcJx7mreeP/16X2CWLteP0HHXOOEriyLbo+Iaupe3ZMkYifFVyyjBQkXB7D27HBk+E
Min9FQKkZm9QcerZzyYAAgimKWcc8V6lMZMOHuS87LacEpbVrx5YXybrIrHivgl5sZrxIC/ZAO6k
buebBIa8fcf9EL73fzbW2SHEsDrbfTbzgs0KrPAeksVw8MLByvmvdAzrXp7QZ1kx6+VZ3jIhIlbs
fvtPEl8TOm6qV3voHRXMwARXjgSVyG7rnI2/XMiZ1FtV2aq+Kkll7rRfxWBE6uRhSoSy+ZLfIJ5y
dRPPRFBbKZWEW/3KqSwCG+ga3wtYgy5mvGF90wDdEqZMQ0x2BjXAr+JhwDMxl0Dhrk/AfagpJV3f
UwaLOnyUku0XnhQWSx8xYJEZI+cM6vWLFSCoT2XHWuS0vwWMfUaQFKaU/tIrwfrLUigqRN7QDdWV
tD1WKU4PRWPOAssdgdxPbhp0q1zq32I9QbzFmFUsrHzsrkEZavTyGwBeMKPo1MvGBB6PzXYioQbX
4TdRGzr7dYId/o9yekcrICEcZvcpiD7ekLw6wSKBe3+p4ojmPbgoU9/G1cJnieLy7tkUt4TaW1t2
dICxzAo5H9eDZyu0syc42dDgYNf8RDkPRJ0flGRq1w4noZzi2VuxoWLFBQnARsRvGTxOfMK2SI2k
mx4hX7sv/mmIrr1FumcqT93Wcolj77iSUKO6uANuzXp3M26EGpnPGSjBRkaAILf5bsuq2yiDBSol
U7ZTzCnTPHZbdawbVBOgo8eUFIP3Fbe4FNRo6xW+4+HhHgOdTUUzPB3Z2mQwA29O4V76ZzYz+Npp
/V4tA7CZ/650c8GN547aiOa/BiSoZeiaUlwY+bKncghPtO/BTAnSA/Vc2dZW3/xAGP14+fM5pj0W
CB3Jmm4I+0Tc+k+2zauz5ADNndnT8eYy/rrrqQlJtlkxgZ8dopBdcBstZ2WvJIWuQx0psxEyH0lj
pJGjxeIyuwlg6C3U/t+6ELcppBaS4yQ03xh/87SEsIGCWhJHvAcbIobaRePorHg2EuIPbADkMuIy
Lvz7ayzgZWsIiyHCymAb7mGKP5COFuE3oe+JkkKBjk3QWu+xIzHBmxF/o6gcyDGPO7n7MbsbkJPc
zznZvxA9Z1g8DXmWYVDAGd8NhoV/TH4zecdhRBYqo/wMCzBxUXwKipg63Ea8vDvkprmdRKdKIJ2H
xDH3QaSJvBUvwidk/l2W/ZPX4k0YhwjpjM7/XYuuE/qy6t0oE6vAVPKTIe1IIWYEM5sQ1TAN7sp0
A/n3V1s83HxRN1NDMw5dk9CEyhoQN8as9N3s0+aXRIdF7ei+OeuyLx1TwrEBviaPJOc42QKQZUfg
DfBAuE3KQ+Hj50d7KxwGXKIWJv3MblFXpp/No7SGeRrEeNM2kw3Hq+0bT9ixfedov7DaRXYNJWwa
d0/NzWo6EptYtRtvED9+YfeO+JljpgTxc1Zes9ziaCAqc4YWtCMvkS5Cu9C/zy+29n8Qnaw0/ebU
hOW/kbUFTRTDDflsGJs+0fZpK9dkeEmsxRiMfgfRj/Ta5yZ51QONJNIZh6gH5nbqjvAXKIlg2Ylx
YU2DUQpnmabJXOWwOMWrHKaSDV4HUK3P8GzsQg7/9zsmE984WcpzQaqeotidvBmrlw42js+1Thh5
L+Hfhzxohx7VvJeW4K/jCs7jv3zDt0DDElQVAkIKrzubqIF13paLnO8Ow3dkUdlIUp/ep+jkQy5O
ovcYIq4HLz/kJ9RlP8vjLndAESpuHgr/EMO0aW7v/jdzGp3/nH1PBcf375R6BiiQWgH+MqJdv2sX
kKUU6fHnLirAtmh47ethUGkqubc2QNVuTJzqXCIDFIXxdZ7cZ2uy7S+19464L//3EjUdyP0KnYoU
rDBj7xaMQAoUWupm4jbv5x2rW8KpZOSTQOs+OIY9WeCMOjSzxhKbHCF81yPYOePvN/QrxzOvq4H6
ZzbfCRYxuQUQozCmOR2521mF6KcZPo1WAI5AESaGz7P7CgNDOujK9FGXeMLdadyGoS5PbzsbYcoo
Re74TbzXgB2jFMY2b2I3UpZ9XHWLfvFA5rz7W0qxq5ZcujwKTDk8Dw1aiviBfAQ4VroDb5S7/RV6
7qrXBKS3gEwzPssb9/atUFeRXv+6rQAIWOY7rFbH5UbHE3vaTdSGJtLujDScieZaIs2HRIgpdxH1
O7HzLHeGiOVYu/ykW/QWA7KoWuDYbb0AAVqc6dt21PSZuV7CX6DuCGe+2RKi4XwLbL0Rx5e9bZcP
Q1O1L8BLfJ1CzSzEiURaRnMqdUGqqhKM/3Y6AodDy3u69qQxidNEd8NqvIFeCjkxS3GzZVTV+0B6
0YIrKmtNGk5qgp5Pekgv6wUqSQ46+whhlhqoLp65H5HryfJhsP9EoxaDvFAMHiTda+ScboKjyLVo
yqxOEZxFswPWLgodQ/LWJ5U9I13fuTYDgNgvgcMutwfeZOwChyVSER3/kUteRBAjrqv+Hom5wPCw
ruQ2XdEweO4qxZXm3d9Z4wGANsexE9zpw9ByHm4bdXcpLbXz1ZlO7lVu2zx7OrYFp7axphWHF8/r
QugXOIFQ9x8Q8Yh0qYFGWLALEbFQ1LXvZenu0BtM591MSneX/4Bubj3mZWu9biFOA5A0BsMhqDvw
CtEqFMMlEH7SnurxLfYYQjMwsk1HFei3llXC3VVsGj+uZ8/tu3dNl4k3dGy7PDUhorZq9htEzY8W
FAioxQMSloulNjHjJ77n58D8A/JHiQ4cpbEizB86uz1OMws+gt8uSJq8OwzYHIKHdwDcwTrfc/py
9hD/isYEj8yKiuU6Kwyi5MV13QVEmrdhSnsmi+cavHdCHUQQ08dRbYfPhvlDObfFlJPwOzXVBFJC
r24Xxlr7J0r/lEhJGbvEtRj8YsoOP4j+0XZNNWktNiCUBWQyV9Y7ZEX7BV2O8Qfdc0cuRDTZf0ny
9GJ80WYaGi1zDNi/pTTeyjy2ZhrzjIL1NARrGc/ZjHhGYDjz0PO4TvVs2WUjVlYEG0DtKsUCQEK5
wfv84YeRSY4UXGpIcPK7OdNdiJMVbcrMfHzRLkJtlsfZU4oACW1Np751swZTBOFhah6B2qh7Bs8E
7rNFmVghVkPWzBXC3Y+/AdX9vCy9vjm2n081H1fe8gbD/+YCpzC22kS1CWBM7v/g0zfULHT/oHR4
d+6TQGw64S8ZOZWd8eSWKxzZuDMJok53KFAAmdiizaaop/KY9nTk7lC//iAjAY6GcxT0jbJCzAvq
p0E7njMCu2waecjqd3c5JK5HVJZViMsiRTCUAx/mhwXdCh0zHljA1KudAl98gZDlAyQIRgX4Sfjw
DbafPf3cYF37XZTtqk1884Bh1L/lCWDZbSgyTfmtBWX2GvDs7a0AnD9Cr8p+u8SQBGAoNu1HmS27
7fswjRijlUeHJfvH4JYPkO9W8QgpaqhKJBPEIKrd7tH6EEKY0IwgV31JqW/H7Yns0470CLA8GnFq
8IzHaXccgVqestVHJ0ffPuBIOWzLqpB3SZLW64fmfEawAflOC3bzurYVD7rAxi3v18ekA1jNv2yt
izwPwY1hc4ixveFi0sLlaBh95PGft9ecb7FvShbOtX1DsPupjL7IagCghqaEcGUPF/5+16XV22mq
5zjh4XFONQs7Dq/CedDBTcbHVRG4IYB8xr82+l2rJLox4miTtmlgD/2NCxWWlhGKa3un/E8WSWwY
mpuXhDmZMb8aXXJzIm+E1Ol7cPf/QXXieUHERkCiufCxNOQPjrd10abON7JlX0KcGC5TUrBUOYhK
JZX5qQwQKXn+sx55cSbyrN1ck3BiroxTih5b6uOnErmxPlMq2SJ6ra1835h7eHnuCDfZlbSUMZ6t
+oai7/97B2KmJNQ1JUMC2vPnIrKCxuGYFEH/6NIkhjKlx5pkNM3u0kieVZ0aUaKAlo8DlJxGnQe+
ZBTzxgidCASCwChaVrmIFFMagvqYnfpgHyZHCKfRpt8UF45v7FbhUI4b+aHIWcwgzG+lUZCiY3Kq
S0Gw4SRVnmWjwzOnNKuWAe1fAblRcpxIcqzhQjIRO9i3DLizdCZHRL/UFOIWDRUmk9y/z+nf3FSt
aiesGPRLPBozUZd7VHd9qdSPPwCf1wSggvESDvI/U/IM6t31ps+N9tUVJ0uVdLALil6l5swq930T
3LyJ5Zdkt39ZVS7d594RroRXGye91dfyKS48XurRFIsiLdG3YWj6XzeidNj1jvQq3N8TY6thLBUp
wyc5btJ7L1+aqTSV/kFFvs0Z4RaW3oQyqRJg84XY4qq1mQ4EO2/PhqcyLd76CH56MY64wvFb6iat
Ls8PUIuB34Nsm0T03cv6DUuZK3AzbvqdkwE020R51Nbov/1VSg+19FzrqZK6KDA/Hck9V6ATC72I
uiovHOISVTS0QcQRG9IV8kMEmju2lxo5LkbwwzpCvv/KKr1JaFdqc/1C+O5KpEPBKxl9JYB3gGds
FyAD2KN99LEV/YyIiwNxs/v7r35VYIRBqXhz4fHCO96bW1wX50cmzRwk9HQvnO8sF4wNXZVUdDHE
qbYfaxtcHaXL3XSPc9MjvqzPfh+EM3307ZxnkJajAfjy+pnqcjmCxafY3+UBbk5JEbhH2LaNqKoo
CE9E1X0q3VmGKPltoEyCyYErd6FGwAs8KuxjIQei3qD83nuiO81ZIwhMJc3ek1IF8kZ2qtRlB/EM
Minwp0cA+KKxU1k8bFYmdl9mT99tMm56c7VfEUCzAr2XAHn7nXB2XOAOHxFT28uYsw3Pj1tkJIzJ
59uD4Lq3fDbfB3c3Aj5eZjqM8Xiio/p+krnUGXiH3fZmwUEkLDRGO9iF6ghP6XcyNjIqigLJC1pp
jsoDMbci2zQV8NXX3tBOrNy+cHWuZR1e6pucMUAuISuCgxTBrKHp2zv4TmxieO24YP7xkSeNHdfw
m/CorVD1s0ih4aRwYC2YRZ1KtAHGvBCOaa7gqUWMNggQlRcdK418blsSjKKgCVNU0qJ0D3jIWGeL
IIpBzGWB0ZJNYiEp16Te6xdnwaI6kqMkmL5xODioS91/HiXPX3FuubzAUlZOvzQS1I28g7eM7i9j
+/LdzR0EQPKzv1j1/87cTinV3uv6sqG0EZWZmgPmxiOAzWXP0WoJGowPeER1vnQYMaxIEtzXJVPG
G3/DHse8EHuRj78Mt3z6gdkMsFACcf6wkmdtJT6uds3NsvesCf29ycyFhbxf7bGumGvBe6nZNrxc
ef7urwwkLdE2yBHIY3ILGdPvkdMRp8FAnEzh9qWbAwVmPZUGpllebQ4lDpyeRlB6kH+bgBirVhia
bbsbOyoT9zh9oKpQqkbLy36MF48sdu1ZGmoRk/gQz5Ig89DwxSI+xdyvlQl7OB7JwJx69vXe+upg
UIAx0EdSkWgx6BKIem4Z/sFVsNyHFtTFR3EfKRs4l+hCJ87CZvVNMk0ZgC/QLmL4Jv2hVBbBVl3p
22fKxL1icu/TvKn1tuNdSPGOsz5K8L/Z8tw5E/VUHf53JdQYh8mECDDtN5m02SAbMRZg1BjMU1Se
nHDBf0tIPWi0r6LrO6BMTrekG9CHllEDgGPzkE0OBSovcE7nmpoANHQm55HQ5gbdDM8P9Ej5634J
ihCEWbPENtHmrHAaueqh0uqoBksPE9Omwt1T2e7DpLnVCBSR12g/QTIXEuLIgzrvA954CG8pEHIJ
GLjFvQ7JZszgIYAFEURTl2a9bBVkjX3yPhIEL07o27gh3yNkmDZ4NBn1u2b7spco6aRyk4DIqivI
4lnJsYdU6TMSUxIDC+SP1hwDxbS+voam/5qng3Eo8BOeOm+ih3EwvHp1ChAvpqEjQv+tja5lTgsG
hzO6FTAaLUHGeJ2nDnHxEwEeXxuVcWteGUCTSlgalNoKsU010QlxsSZ5kG63vtCLTIwkqUP6F8QF
nmhdKcseFdL4bUWj4TJsxqHg3Ve5BpPDuuBoAgSq/CYvuRnvEGJhxWZK5oL2Ln2sq+qp571YI4Hz
zZzVbOAWqPk5tBmKr37Xt9SureG9bEB7mihggJgn19EKd6orhkmFYX7IqNFAu+lwCR6uxRifr0aW
vvCNRgYsCg7AtSQ8sgoTJIbmMB/tJW6toR/f3ERM7g1f+i+F31YiB0mOzQ/As/86nKy3YwpquRlh
VaTwlWFS4LiKOI1GkYfRQazelNFBOecXE1zSipyMJCQvjQcAGFVrkhuKAQ7BkknJ9TOYlrmjc6ok
SBb3Bd3i5rIpeH0ZuEe9CoeUSXhbxGGESe8mwBg5UYbK6ijOgRCk5GFF4nKbQRHaxzN2bXAagDQO
h3AVF+0UE4kAciXRXbLWIwIcfo0+MFWdA3u1/WEGOUS9KlfylltZt96SImyggw3U5A2/sGCAnLPY
3e7NrpCmQugWuTqdBlOn3AUQkD67Po2U8hmVrUVMGoPYFLUzl95QTvR9y1FfWyiGz/tGiIBdbwcF
iGLOCtrMwEgF4F1/l0BIq7+bFMtW6DSP2kueE8zZZJKVttitLO7bHdn1y6DwcCleOJ6Efbia16aM
cDovozE92biNtqN3NWTGrrxA/ifWUdzktr4M8W4USj1RH28JoUdqdMxesR+pEP79FEM0PgeGf1hR
Bs9HiGWqQX40/PbfUfCoMndNWdrbeoMmhU709MyHC9GwDwSsdDDny0a57UjEidCfpjh0htfAnId7
2mtAp17u0d9xMoMi8QaAAXoiD71Z1hdsojoTrs6x1IW7jjOQbQ2lnCvl6/oAAeK7czUKo7tZ9J+3
KUHyg7Ye6Vy/c9uWlpUwGnMlzAL0IIyrnzHwL40qPGY4NBzl4MsLN4swo1OgQr4sWrGeE6NUeCjq
X/DvJJdxvS0ESa3lxWQX73hXr5NydytOc+6aqsGk0Is1M4CgnHkRk82cd8icF96m7KuEHl46AYTr
h3vIAOMbPdgb/bY5gOz83gIzIgBMLEm3N2CmAtGpe9JRcczD67euMRsvVmDnm+WImwezgyBZshD1
NK5ulxhbnIbIl87+kgEBcvvivGv6bPLgkJt94SFssDAlBgd3w5f4AqIUV0zL2xzSElLGrRO+V4m/
pDGEk4ne+6zkjtpX7CUkPQ2EH8V5hWr4Z33QC60Xrsp7O1Skhm5q122/CA4eCMzAJma9osP3KnR+
oyAazBwAk7df5xSnWL4EDJTysrkhMj2U4KhZcPbgUt5apeexOLIoKPR5Tb7JX3cv1q6o3rWI+ZW/
5gGew8M45QERl0RN03NOcCO2BpRuz4EM1FnV8QLZPWau5rAsb9Nz/yN+DyrytW/+iawSt/WhsbW2
UwzKRph+H4kl9FpvcbzIujIoxAY/FavJ8XLBIl/jVVQyS2sfGTRe9fvjHnoz/i4MHemilsN2JYDr
cMV7gdACXS96sEjcO3+ebUYI1z4dobTVQOKG9so95x/ud+kj2TaUWLAfazrYJo5vTbuKWwO6qKL7
W4NHtdVkjE1CMY2zXiO5xFTLxaDYPjA+xV5sWb1gMrDHOTgK0n2VsAOtqlFpU91+xBJofh945fH9
psA1xrQuRZvIENwES1z7oCyL/0LOh436Y+TQ9xncQBwLumVcjlqI161UQBvrdX+4boEyfLZoQGXX
CJSH9SzF53SkQqOTp9RH2HbULiJHmLXgPAxnlLnvB43cJFFHseBD6uAEguqov4Q2LYoafTDld0q6
H5wZcCKovD01qyhj6QWan7gSUuSZLwwtjvyzPvsX6304Wx7UE5M7sDRgN+Fsx+wQSjSM4xno14eb
tadlbkYUhf09IDI9mDmTO6+5IxqYUDfd/z87yP/Tqy+PdvJfYb4doGJSBy6+fY+LZ+wzdmLwFmKX
fjmptMLCXqPX5/K4BPtXoiJFAy4Oun2njunZ1L+v5lb/BMQmo29mgfyCV49yznW1YzIUKYjCDpcA
42/L+82kQPrPJN3dAns1z76imZwXB8o18gdEVfjY+X+jYxY+TvRmTGygcFo9Fh42QNPvs2QXEFvn
uUyEbltI7Q46UwLp9g9AdF78my2nJTKhjmJtfbvbrjhUMdcr4L0nkYeTzvGNxVlHKkXRvm4J4a7Z
CQUTnCFFXNXCbnsxYvON8yOW/pJnW8513U6uNeWfYxdtE4D4b/A3ug7H/dFGbqRpHQJJevkiQnuN
xGmk5NKzDCmy84ijQdl4WFx2wHnRB6nqqgMYmGBZR6W7qS9ijrBfCbMbP14FOTs4aZXi8PFAgBH8
ms3lnNH0DI+90gFKDR2m70gWJb2RfkMwbmAJQD6P3JEmSCZ/h+q1L4YWeXDd3uL1zL5eOWZ/nQaS
KEPLpVyLqnrjDpG012mmXUSShU1NN7g78XFUQSqg4mEEOgsYlJQmiMk1rVuwq/vAF8UwN/e0hTT4
hHfUUbE2VxjkkJMBTlfsEklScscjK4flBlr7O2TQkFZRimUdBzJT1ARCtt4P03kei/arro+gcv5z
MOlLDiLbTiGfkyt4n0Lbo0jZweW2bCBJP2QBTSzrc74SYYPbCgWllnDr/Jr66kjg8jT/e0Spagoi
Z7C09lYHXDimmd+gJbw+3P97m+bUibRs6QS5u8tI9XnrFH8mno7Ks1LoSii/3I5SD5FiT4FHSqPt
0IOJIVo47UaAN/ONDMOtNUQWumX1s0SJQgs//glq8CHfukWifCVhvcB+1NFQ0aM2N0xwSU+ZnMba
jfAlTSYsfwqMne7C+Lt65g21q/BkVkbQeBRIiJD7+IQ3lz5VmUv5/1rf10sC0atXw1VtQpk8XMtM
xNDb0g0kXtV8uLuhdKK7T2iSCQu+hE3iCoqhvr6wy1GI1we6+COER3biNxeWw5Dhnorw/41J7Bn3
znZ8kxDbV/eYIZOAa8x6ex/ILKs2PTN/56ibcfXE2i49qs9+px2HdRhg3QLSLI7EgZQYfGqW/vxH
wFPerI8EFuFWyQY00qSq2dPrZNOuByRAJif7IDNI9yZraMQwH1i3R1QFVlFHHVvEIhVKrEdGU2iN
ToMAc91N1Z2JPUGNgI3EpIOuym276A6fmry3EPKYglhdVH2qn8CC6FbNOHjVytx/PT9034HABc7Q
Nj5xBEzbhp3uJjNlAI+lZTfyuCwdWi80YpWwm7kF4J/MXRCBRa96dQ8n3wI0OiHcCJlZ9e/ydVNp
sDEboQhZzAbGhXf73NoURDcuKStcYFlNG3dhVJu2H/dDd5m3omSfxzMVec9fJRiUykzUREG8aYcU
QT5AA8NM2THwxOf2VsVbQg4lIRD3zizXEdF3HGgfpgBQ7yNBfeIcIHhDd3jN04/6bdTtA9UFQ0OY
VAMaa3jHdrTeJNo9I89Bqgi0hpiDuNor32qtzHS9/LTzNwtRGyvP4Tv9sdw1926ImV8Mrm9mPBnl
SQua0QW5G+AnVRLpA2bMYTledEDzqXHDfTY4580PphKx2bfIu/3H568TFSniK5g0lQxVAYsMTyk4
uq0s5oiVmrAUqoREyUsxWs1BCAid3LtRwQYgc4z712TXk/df9OZScRTIj0EJC+NB9+t38SM9fwXf
p2kWOR72nmpHKiQNp3g0vFwXFasvMO3a/jxEFnXDqpBGqjuDixJWWEfmaQ3sWRxQJF21k2XfwDtE
ObGewqTpMY9vh9C12VEFEO+H8ihOyZeooSuXOaEkwhSiHJp94WtYAiH2CYAm0XWL5Dl98VH2f2W3
MoZ9O/uCFJQnZE+b5579ZzVQkjtwXZIbaIqImaV9uD52nj8itebKakML03muaCn6jbYO7vUsq574
0Jl1MqEkfVtmIghNvkwcGlxS0nEsAiD1UgL9FHgdc89kAgFX7AswLBSWYtVvZeWmeApj8vLzr2LH
NUo1PxKr36kvJaJcZ8xxEcj3Ss1c8UUArwXsmnqKjDRvnb19WnPG40S32NF9bphgU9K3f3uHDihp
z2RvpP5VtAyHfFAlVGEfPB/39ZJKDwf4ziqioqengaYdJsx4GXe1HstZriznezDfhdLHUD79pi6y
IjOzXKFmVnc2fA5tbAcn1qbwu73QSnVy+EsCiwWHsaTLeRs6/3Wfs7aP7GO+ReSN9BU+fjZJerlh
p7hi8YY8u4BgnHCDr1BHKFh9NSEKBJpV2mxyocqRLqYg+Nk3khCYlz9UmtjjmA/Y6ziEB6HmABrA
6Dmj+IMKh9HEnE50os6C+3KpmRS8pOVC5+l1RDXx9aDm9ed5PjvlVWaztrm7aq0c6cY+/j6uAVzK
kVkiYhcoZYGLQ4Ku+bQftODeqmA0MyNUHnGCjN/Z5CVmNMlOlwW8GV5X6da1YsGHviUdGdTt6aKF
STcS4WcpQKWF+7x5bwDvWv2psfSDKg4I7sZW7vBRt1GSQjZlMdPBMd5pprHMppO+q0+90wdSdorN
d+BDQurYqoHMK1o/mVqXfox4AjN+b4hA74ZM5j45NwItUXkpb6486yu08p8ycOqdcGs6WW0NUjWj
UK3RmENQqD9yrNNgwhJjUqHnnt/f6UmmYNnyFvQWFeaCpcsmZkXEiGh+LPHW/H2DOMFSVUNxkD/q
CdFDEc6NbtsAmtCAJB7lhJTnbyE/xzOyfPLBFskuUS+eaFSsXppgjeME3g+4/fRKv0NF8/J9uLev
xn99ypQM4SVXCQO8EQhJRbuR3eixUaOCkuPVKV5GGTsi2bQR6CiYiT06YYBWLiPLOS080W/qC/aD
0WI5cBm0mgAsuW7qB1wBq4BXvHLiPhBeaJ03V6nVUWxt/wlTbGZXCHdkEVvj+rve8QHwWyTS9Q+L
ZfJsOMtHBIJkUX1JQ4Ak84Pu5NZfRuQSxqtPMjNEoy00JtItcfDe/rifegx3G4LMluGVWRr6Wp5j
fk4hNM64YxElu4+O3G6Hps+kVB1aUflOPi8UC2+Rk1pVgCcZUW58kZJF0hxjh4imNP2+18GDThsZ
HavSwT4FrwV4/84GNMMPYzT3y5y/0Z5oYV5u6A3jVApUH/7B9k0J65ZbK/OoBunh771D/WUd/Ngi
oGUHihpSRhEymx4korZ2xdvwx3pxePW3VU8E9JF7ibaZMNm0zU0Pb14y4AOwhq6ifLP7k9IwWQ3M
RLzACsNow+cnOkPOa/kpsRxkx0cjferWLVDERFU9DGTq6TTrSWVkZ2hvA5wFAaigQZrA5MdJkpzz
y9KwBwTJgtwZ5bwdjp795pTanstIWKeeWwsLAWbTIeMsDYqCc4q2iK/exedjRqr4glLB4eZlqo8P
HEW+L3VOE7LycYxVsSMxG0odW8SkTw+kgWPPAscssCk766IzVRIuhyEeZWSL2E/iFxs6ErZ6KUAR
1pRvuu9veqaO8Fzgi/8Edg5TWIhVp2co9LYTkDVkB+fVeXmyiQa1+G3+BleAUtN4Ud9terbScOQ8
CDRtKyvGSzjVsObk61SAw7RRNeKRnVRSvAMk8L7VTzQ1GvOQxOqKS9LQIV1NtX3Axi2ABZBl3jVY
eRZFomiGFy7EEs+hTc5hAqIOtmqXUy8x9MuxxzJX1eSgaieK4L3ebQo8OezUxInBonEdU9krWXUK
tA85ZmcOgze6c060Oj7FUdSHJlJN/wp1GzYl1Cc253aI4XdUXdvN4PWeH2V2nmBD6PTGXTn3yQQn
Gd/KQgxI0i+XP6NSGAEraqFwJjkQGGi5AQej2Tjjx7HfD08N494ayzHvcVLwOjap7a0WI5iFhYuS
9sNaqHyd4gbQMsusCmUG5tpfHTbUbej6WXRqcvG0pPeDScRN62vOqYa6V+sdJYkcL7urt8d5QiQG
GS5kw6RJdGi6UNflhbv0aQtJLddcoyl5+Oyxubm87q15Yil2ZNit4qMjOXGTJLKQC2B/TXZw3wN1
z27o6Pg01fLwxnKuk5VRlojJC5cd9IkT2Zl1HHCu5228YvUP50i7pT4744svH1k1MvBhvrtpGYCo
2DGWaJ2KRrjti3sQHMt1sljPeZmq4sbmqiyI6mepGbl/Av1gn99kdmPR9EK4MFIwtyEkSl/2XeRo
yui1K5904epJM3N3d3PV/R0ao6R5amInTRxlDW55lpNu06uIn6ARIQxjz1mZf3nfufetfHODKDyO
CMUi/0BlGP45AcJJmujlhUqxpG887eOUMKYzK1sg5owE5mr3KkiSs+en3XS0x955AbY6N1AEytVm
Lm+P5c9798K4hAV695qdv5jlkKyojLpInLvfM2NT7zvOLuPLII1GnAkHx6sXn1fK7p5OQCAcm8WL
Pyma5Ko/wq1I5U5BrrcEXCNS5bvUMTPImrn2loGfx3zZT3vbmDT12c08UgYfrdt1m+DiPuZhoG9R
d47uMMOHKGCWLGSaMvFmFcuLPFU+CKmyJbNma/HFF1Yt6iz6QfcjCajnsGF2HdTSfgbyNm0SYWhi
d9eFPsatH8+HMiObc8WySQ0Ra/rdodeBksQ3qtQv2n5TjtkgLLtwBHchff/CAf6Ep8S/9D4gRxsi
h6yYD3FZDW51ieZ9xhQIVZCyIedqfZDcX72Nzek/EKk24hq9n44micwjIUBP0VGhPVDNTl10S4tH
zanyO1rjxuXdYqm/19tVxjvCP+wI6jM0YHdp1NOmfmXxf1cTcEO0CnQzQD6PPBwDBL7eP/beIOda
+LxlMtBdYAYQaNe+dNRA6qXLbNwsGEsI5AswWutMu5PaCYdwY/ekpZS1WxARgNaXy5nwLSqPk9CC
Q8tQWqK2vYPqEafEFdqgQDdsWJP/e1VANDujxeHmn9PrkL9ji59ufy9dIXV0eLDrK3K3BwnmMFU6
T4T8WsL1n6YUA7uYNlSth9gk2vMGxHY8y4UcT44u7nyvS5fGUsq29X2QucDh0drTd7v2iqt+EzUU
PoFWyCcXJWyT1FpzNYPllO/mVMeV5SmBPt8uShdxzY5M6pZmm6sbZkVK7f+zOW+q0+HviN7nJDnB
EF14lRju9xThnRR+5yFueMeHuRDUPbW0GJKYGukRA/nW0rwctaq+XmbMSFSdz0XrptBcr7qiZrh0
EXVgEkhvz8Qby2XzwBegZ6EakruAk6TkrNBJ79y7IT3rZf8BXEsQUVTfEB7omVCz62Uy78k8oQGm
6/smrhcuW0bUOUBD4SE7x4s05Pl/blqfvWDqVxFsFXU2kLlsWIpX2BDVwALFy0pCI/iJyEH4TQxG
cLJQ9nMMSGQ/5WOLTLW0tQVC+Y2AYXNhx6XiB8QDpay/ge3YeCGozHglGBOsMo5sAETOcpoO8OR6
1DT11XH31yXkQhaseP8xMhLOAPWoVHyvnKs+MeFAM01uFD2rSjjdfQxaIpJdb+gT/elssr1bRMxR
CiJgx///xawRPZYsZBZF9HA/gncj/+o1LM1NM453F6/wDp+Jt4NqIMqati+4GbbBr22YDaPra6EI
8s/SpnVul6kI4G26ZtWktSgWriLvmo30DBbNX1S3dT4kfzB3WvvR7z1kcDSyS/6fxbkcqj4teU0E
VRm+C9MnQRDG1xzlaxhgTTpBR2C1DvmK9b4XdFvPTgZXEaHL32hUgpnzd6zh82XHldcBCVtVSxtb
sUK1O9ieavVmgjUqxC8xwujheUq8JXEFhD5UW5KVamCQ8wdGLrd5gnuzSdAQbgIN0d1/mdBnGxoy
nSkw1AikA2HkU79jSyQKrdMW1o9Cyrhjw1o2XJBDNB4JnSACsoR2wdxwcv/kTdNhgCO6dLO/VZcA
ZCGaL9VoI662TgkIVePPee1lUtfPxM90+u/yimKCZhKtLezpBfDlcUu1D+PYeqDFDARThKy6eysP
ufEXXYexo8LBSVaUxnoFw27NiImYGtE04P6XVYy5EnS4wy+VkKf3AYPGhlnqny0D4Bkb0CIo5cI6
ZsUhoJqeWtK/xfvQWeoZHwlBPoXOQwBk+usAewXKe5I7nO2WfMevXOgixVjDkTWa3NpOuKS0dImP
KdxHL+NjBYzRdfBKGvZPVuYBXGzuPDmUrT8Sxfzygj3STZ+7LEMa6faknTlLG5bTzwswSGwigtIH
+ziUROlHxGADa7LMjXwFt/1mwFn5SXKGgzOBFRFOfe3/TSoXLyI2n81pnAe3myXwRqCN2+viN8Nr
/DmP7MW6xdYbEyHJIGeY3ZNxvtJYV5CkO2ECALHfyO/xMGmjuxloWDimHJEw8Itvwa+MAuopNfMn
V6gL2z/RCn7jMvqOx5aY7cb7mxWZfZn1gfs3dwg60OohEdfOZYBAmUvw4vQT/zL7+Z/WvwG7iSaW
OKmYpxThnRLoO1mTNzYy6TvHrN/iplew0gtSRTiweZukoPI/Qkv5cbVdPsann4Whto91fpcz4xPl
8mGOCoSp6FgHDKrHdr7NtycrYFxw1uUStYKFRJvWUwWYjvO4sExeQ02g3lQNqwIpKEGcyhKFF2PE
Z/frevVsBdb7yLfTX8gza1P2HY+PKHi06UATkLHAiIayDwI1p3VBzi8FYi5Pf9YFMDNVY3cJuyNW
pC2K3pIZW2+qI1kXjFhh3D7NxWKH6Sl/NDtebu7ILqpJ/++kOpX2/7tiPTtvod/VtK/M326/cMOR
1qpVH8jWO0v5TSn9ZmWlkobtjzpW6/xFM+6dZhxvCqTNgj8xnNjLm2h/+840e7smvnY56z7mcCGg
O8SQYjRtVibkLU9MXPdJ4J/3Y9iuXak1XsEdXsjw/owgGUzATqYKbhnSNvE5lZM1fznSce59D7WE
CXLcdBf+4dsRuarEz0LYTsMPR+XwEpkpJ2T3npqvSaixdJneVNLIfELOeGd7HLcglgk8XDknrBlZ
c2j36ze/5Xc6ZRPaoGglAASWl48/NspgAxWNnaNsI2cUQ81+kXflvINbUo7g14ljzrgmS3dC0Wak
1QbnwBWppop/Lq+KkczRHddB+hQ8h4JcXb1f4AXmv3EmdOPglD0kLXa6s8CTAeOW6maAHGRJIWdc
UlzXxnkAMrGuxAeg0Ts7nSBVUFs/lnALbKolyMhUJBGiWlocBznGalmY8YR6tiSXp3fv9+5KKmuY
ZLUVcgu2Odb2228pwZ1rYqDPJHKM02tSWC6MX1fKb4kaigCJbXat3yFUm3CLZs1lew3yW4cJKuQb
E1gpqQhDhU397KHypgizT1aFpZS6QmngptK0IyDf6Uq7B5/f2TbKzB0q76kUtruoORbe1b2N4o9W
m+3pvuBrbnYKaVr4ucbHrZY5KLMJswir/y/Y/9QblE2dt98XKHZEqKluw6UzGT7jIeMI8K8zKMKu
FofF4qnks3tIKEV4tqhATuupyr5tUp+eDhPB9EoJ0ApPm/WgvmaJEiumsIRCmm4vCBDuCgZc9S5f
ePjP1QUjfjgDEleyZieZF4cRoKEkUN+NgPggSqpl94CS7da7yNEqIxZc5OYssXCAUDEKQEZ2aqA0
nGKhfT3X0hHpPQ7LNCRGljrKwBGL74XBqyk4Hxw/H3CNfqJqnQmjKPgRT2+Ad6s3G+RkASk5mYOU
B1LUvV/1zf1vLfaEbazXRqo/2R79Qr7UKAx5dDegBKprJkPqQG2lMSpBPXFWDHxVJvxqoooLqe8L
4XpBpTCB3uaLshKjNVpTKf1WJHzdwj5GCS9Qt8Jw0vsqrM141z4kEudRPw7rOf79k+CD/lrnRogO
OCdETMQNC+9ROzhPLYkTFk8i1cGVvzp5zxgJ4yhHpiML+46Er2VI6/UEZjB07y9vuUSjpW1G/Q0s
TaDUbiMST9DYTdoBG6jH2mS3AdWOzL0lzoSzuXv04nx+NLsYZrZxGTZMbFqlkbJy5hl2Y5je8EYO
cC4xZ+2UTn0voY3sNESF+aP/4+a0cPE49CmBOX5MRdXlTy3NFBZHWjp45egpXbFgFrOEHHxjlxO2
gUfKh97YD1yscHErn8rQoSuQ30+m1WgiJ9L2xKc+x9R6klxyiny80cKBGBFAN0AVeJGdQexG8425
QoNdwx0l5lla1fLzPA8l8wWWZRWLP9pV8rUZigSqPdOa1uZKEzEFzpfs5nNRhAUy7QIdDXR87vuw
L8NK52NIOGvKTi8hlo+YdvId2fKVJx+dH6nsJZDbY/aT+W3HBZNPKoUY3nXZZCT/fJQ+9mMREozz
LFzNG2ilc/sktKZ+JYAAJqDsndVDnObx4ErqaFLaX0MVoDgYnXG5S3v+9UpZyjQxylY75aWBcH2t
6llB+W+STSMaqJZi3mHINdoUjnBALrvQFod8ncBdYQZSCy64n4aXaY0cEsGfzAyATlRaP6fdXE/G
SmPLerg4Fa1q5bSpRlsMcKmxCgWHOCdSwBIzjEfnk5GVsn+0l60I+k1vyuo3nme86mU/pQoH+WnD
peKLNCV4ky2HS0VlnfTvpjfszbuS+wlTF9w73n7Dub4p+r/G6tRnMY7o48agSz8LynfZ+Amhmymu
eCS14rvx7XzGIjXSgdP5ndEiQfuOdHU9A8ncVo0oxtwlwORmBuMGm30rOXrmzUMvnjHhH0KJIK1/
hy689aSzJ5SKlHS3zN1Lj4QyP/AfF9EUeoBv2eamNwWJvEutdsPhTAhAS1kOUWA5FGKuH7+rIUDf
JFZ73mLTmxCljliiGt61oYjsdXd2SdO0C/+WClR57q+qrReoLj+jeheTWPGRioAyzRGNN2EsUHwK
EFpoH+0I0KMvxLNwqzimtPaDagfsU0mxERpjwjJGMh4eJklL33nXj8S/65NHwwjv5l50nQlKrDV3
sfr7JP+1udqJhOcP9QHjJsxaYbB/CaANZdBqqnbPwhHODrO5tS3hLr+BrqgoR4R/BgAd1b08Y/oc
9phHrkYS1dd7pTAc8Js7L4RfUWxxn5ye34kh63YMuC438GJiYnEKaGY3RJna4h3aqpgzrPKk729G
tJizOnl1x79m8Xt8YXwr5gxO1z1C8n6IQ5nMzAd65Ai22gtiXBBSmJF6GKk4WctU8r1DNSuM6blB
KKGGzLr8K8TbxyoCl1WyD14feCrM7ilN6vUAiNmAvYrLYeEOj+JEUfpqdZGzqmtLTwrmwUApjCLt
7j/zVa0VYQqzcR9eZnWkrj2ZCWJirtIaz0P6Uxx6TPnDwJ+zBBKM7UbC5QgK1ap2Unq+NZxBLbdl
JJY12XenMEAws4pfpRP/T9liUQ8dlKXnq9OYgnExdZjbCgn+hYx8AmbPg4xIlpT4Jgw01jYVLxpg
kIXXLsi+8N/+8TmxGmE5YOO1efxG+HQz9Lkyx3Lb0KaUlE4zqZ4PsecIfMOhqhIstRfj3JvaW4Uf
14jpAicoCixCdY8rIgeTWN6TjB04tKJMQmMiLhifySmQ//Ee5v9QNGnj8mdJW1ExNn23hgEpFWTy
uam/WwoCbBmgKJbNkpCYg2co8YA3jk8p/nZHBJPaEEhS24Th0VbEo4IFDrqXX4vsTNm74Tt4wp3L
G+ZuUDN3SRAKNWuO//O6xoMTr7LKi0QdlpLCQWZ97JyHc6g3BJN/QCBt9c5GMMwNPg+N05n3BAzx
KiSMikz/88mPKde10HL72xfK2i6wmZ85OihXof9RaAE+Q8nm6RRdXGuNZ980QxB73rHV0Ijs/vIS
owNwga0U+GbS5jgD0oG5NmMYR0p2x2/HJQNxRdv9UKJKYkRN/R4YmX35FVz7w78uJB4PuJL6H2Dn
xFB/BOm3HS8uai5E/ud8TO0LAXLJFatNH2e4BXtzwkFADtmGDKub9uJ9Ipa+yDqy4+0mZywQsfg5
+jt63eHsMG95IqQATg5o+x51Fx4IAZbO4kbE87fsnjBT/u0mvjzNUDe6rfKUtbTJ4dtIlQI9+Jwa
ok8u/2Yf0jaSozBstZ7dbpmf/fp3t270jljM3okfL/egFv/+nM1D+dcX5pJOaB8W8aY4eii3482Q
MXTQe6W5QZ1om+KJ/Ixubj5ny0wfq5Y9INSBw5VG8D9xHM8Gho5aYoB8TMgRacA+XPwGo6E2pgFa
xUSpCOy8W3qdrVDfKjrgnJqQXLm8LEagCok+zqXbGHitxa98vWnT7d2uEBtXsll9GDR2k0pzk5Gb
mrux7W7ik2DNhPJptwIfYhrKccFMjsTDvond1khTQzQNLl9lum7gtUvPwjXczhkKv3nHcjOTCRmH
BxZLtRley5twYFULrm1SluT/cA5htjUvAVqi6XGNhIwmvLgdSdF6J1HNq80KqLaJ7nFKIhG6Mv2c
mt7shYuCL4fjXkGC+RBMZGiaiz8PL/r1xgqHinjqAI7T2yNUu66OQ3XtqHOPZGQVZeJh61auqhNM
WDO6PGpXKeG7xSNtXL2CVIQ4rOXtbRiETQ0GhV3FYIN5jvydxVxxbdVLcgoP1SYnj71HSBVBPfWR
+wDxqxB3l6zsCMBC9GuaayGEIuKsFIzUaR34r+o75CC6CmueVR5i5g0KmRJyOg8RGjAle7+TZnoH
4Czng+gfex9JanDor6bQnyIxuHLqxZScoIePyDWaQzGyK4ubSdFU50DaMlBEROe89eDIJN06yYhh
9vwuGMiIl/7xYp8HF3Wes4VT0Lpg4vjOW0w7YZlzF1UY13bvXhfzzz7iCrmFZwZiUSkQ/j2lY4u/
ic1wLksyovbGn7+B/iS2QL8TyniVx8h+Z3gLWJzLmbFjjYbnGAFJG69MaUE8jz4gqGsKZ5isBkhp
ziZgLqZAYvmnLymaEJ0/vZTDV/PFPSL8ES7+CiQ9At62sxiXTDjceIstNwk0NDlPgNCU0y0RjBMk
hanvGtdNLf17cHlY6U217U6Lbe8H3/0ROKB4Sm1JCxc8dG9g4d6WBr/cHMDbz1tRoH1AfXsF5JCx
uVXnoDuR+9ZDniZzLR6B8PMoMr9qRAL28WVyyYU2C8083wE0D9KCuvNeFn9WEnJ8gDym+usAgELE
l4GjQ/JKk3kzvVWiItRa0Zbk/+s/3RdlFy6MjRSGBrKcZ3NuBUr6has+IFqQ4RKUcV7K8xJpEuvS
eL8MdPd77BL3XCuud7UdIrSPvUSaCdhnWyePqWgmwrH9NDB3+QhkI2MNdogVcSC2qGYh648pu0lr
O7J97r71RSsdbovM6ryWAOhHwVl5feLohJY/GR4aa6MH/4DzaWjDLSow8wx1NizyN0Vqn8n/pGF+
E3tKQf7DjRpShY8cy766ffWCjbwvJIiIDSNBpGUxAr9l5sE7ah8NlBQ3Jl4Wb7CDW47+CnxRBUVq
YNucWzt5DcMjMQSaoN6C1bljkmBhPqaDe+n4pZe+hkTI2NOjWzWtkT9Bj2ehzklHBkxgaZoACHrj
WJxsJeTZ5eJF9pqAbSrifS6rA97OrUMrK+pig4xRcCxgwJsR8UA2bKELLYBYucGUOlcbc/x7xH4g
Qug+yHmn+EIjWqbq6Kmmgpl75efFsKceKQJpcVUHpVxJHFlLdgJfBaXoVWyhI8fh06QOdRS/+SvV
ZtTo8n8NmYnIlMSOWZK0amVNQFeZB3vYOUjc8Sqf3uAH9okGNQZuw1LuWQxzud7Sdb6jtob7qLt9
JQb2x/fumsiQZ5VhF/atvDu+H5/0/YhUZJIDUdCgxUfbKu9clB27jR0jBlmjZcI4mCBgWG8+5S/5
ucQOvU7IuA2Ew5XKCdSBzIlfRzSJPD/iQvU1gSB26BhinAF6jUAirvF4ubAAV5xNNLw/GXwsIzpi
idFxNyyOUjewpIwG50MWwZtrc/h0SIlpcWzyetg3TPomkQZVOTue130QUIT9nC7J3Kbk8lQTCu6l
4w3gPJKL+n9iBx18cEMEe14NdJrJSZKMGRV8d+UQvECgKlk2C3Y0nSGzw0hGvZIFATbJ/2L08tBV
zwZuKLaYR5vxElUA9LaTuqkeRRCIg2ezyQ/RZSbTCFLrMOBtNLH2p4fIkkt462lL1goQnt8qT9iS
iitd8yRr5SFjedGMO1H/qQjeOrwJwDxEPntD9OUU5pCwxt3mlr4JJKDc7X+JzCDEAF5oT4q5g5b2
mQrZ/f6RrM4CCcLFv4qHNX8Cfc1gOhcPBQcdw0Hq6G8DIx53eQyy4oW+DcZll8D4YJ3AV/Rfq4dE
z6jjU7p/s7GYCp/vimsctTQA+eyvtoUzHThmXLUlY4jPcsLkqzMC+TPvaGKv24gti6eD417W37hV
ho5MnBWvEkEa2CIp+ZYVmEso/NstwFVWNBHqLPL+Nm5tQ3is7V6tI5eU6dT1eSJWORsanpOZrucO
WEqhDNjXRU99uLfdzgpHMzza+pdvm1nguyQxuHdgjKOEw9o54N37xoADa+ydw2FM2EdQ6YFNofIC
VUAfKTdTPMSC4DPg+IreUaRBPb+ZlgudqW0hVjq+Od7vCeIiUMbaSWVcFNAEAXLdQh2Lc/98Nb+P
Z+sMhYWnrR23bZd/xHD2LVhDVnlijVzU66/19LbuiUH1TXQpmq6/v8JRp3vfj2QIhA+zvoSW5MuJ
jc5YEzfyAOybMcJx8uOm6Igdf/yB+NLxWTOGYy/EqEZ7gX8CvGblSEu5RihNfUx9TKZWsgtKxM0M
xPq3/jM3lOGXGRJO54Ws+DbmdWdamyDTeJB68KEkPCbBjre4YNQyMIQcNxu4zj6WHOw/pQMKIqh6
8pG16P9F0FcFeDujSEHB7evlREX6Xb8ao3M38r13ZiBRMgweibx5CPP9gq9DklaMIDhw++84JYh9
GdTlIKKKMBR1We+CtbNkdL0EWUy1cHbsl0XHwW/E12HEDRWb80ljx/PJdmryUJp9oXGdY/Mo9dOT
uQIHFcWIsxIjKSV1zwA1kC/M3dbb6esIlqnQS4wZKuv1LbsYG96JGMD2UURZJWFrWDRqfONr2sFT
LyAWehi27FekEhyDk4T11RqsNYFZ3tkYmhzEcNODbFrMBjjnBdJ6PCd/mOAgrTyokrucrcvpTlHL
SCSus/Yk+NLewYrW4Ew9y8o3a4NW9q2iJdj4NB1li3DvLPRKtRfQ00DVYousUd2Inmh75eQMU9kM
pEjk/aH5CouXOPpvdWcie8zWfSt6K3zlM+D5aKaNqQVEFedI1FWHHiJLlU7lALqISjk5d9BnpGDo
5hmu6mVl5FmCv/pSszHnvs2rNh9jEnnx1H+o1bKZ3GTolXB5CZd+pb/DwOUbhQ5iMyYIgVvaoTOR
mleMDyu2HhsJq6olu3j+dqu/1zvzb/01LZjxOmbnXE+rkUaCUeEhG0e+DqKBBzYD7rLMg7DftVV7
zMB6sOxiTrtVJXcLxnorFOB3ByeFDlZIVSbXCsdsw0fT3Mkb20hOku4Dyl8MUX6yXhYmc7CR1F/4
Tx1XAKE0FVRlCsBoC7e3AMKzBYTOTEnJRqjC5mGk1qu6eyOA/c2wWjhkoqQQN6GMuGv6ESTJ7dj6
DZ29jKuKZSCDNwVpbjIQFiWRcCTCZH7QEFMQkG8ezi5AP8Wm1pvY0yLsG5bolXSWx0IaNJ/Z7uLf
SL7OR4ZmkkZ2W4LAybVUM6aMHmjsHwZ6Tr+SRk5JWMMkjuMC/VSN0UgXEgf5hPRWITKwQYGaQwOj
RzBC1XYO6G9AWf3IwV0t5p479gkIrPvgPoQCYQbYWU8EWJ2eWJritqJI61WzMNqfGRCMipEqWpu2
UgU09xXdJuODVKFTAYR360tSwG0wU8ae/3fYswJPccR6/wdSKvhkjL3VhGvuj/ZlLP+erB2t4voI
XGitptifkLlAVK2mUPEBh+5bC5M8jpVuF2ttehGwSIhUZviaP9GOl6YRKE16wSLdqcgMAtLEtUer
gLoC6gfxoh93yQ+hFkYYzbYns5QurD+/VibeP207/3dOeiyPrna1ViFm3DjhFdiGP7uPgVxasp33
4Y/PhT2/clQECMjiFOSi8332VSiuUJiEUEr/k+4SYK72pZn8gSAv3XlPVFG6hYT9scld/BFa7anx
BQ511+ckwka7E9ZZeu5h52MeNqwDSZ3G4OGvn4vqk0MQDdBXDb3S/B+o9YJ8ABxk8q2adtEAX/1N
Wx3CrcukThluSNoMrskMk3uYYgxGZ29435u2Pw7rvw5xqydClfPWI/o6sWb/5Cz4nECJCXa3lCKs
3KmMfvHfe5B3fHrqTOioDiWS6k2L9hD+Xu/PumiJNIxTHYimIvu3g7HDL0DdFTo7Is2KKEIdTuKV
iz2Jqx/lBTeSSZvNr6uTbjlOIhq1XwvrudxYzLS+GUR5fQokfSnD9yCSh33IcPybyBJaORAZG7l2
nApGpb5k0Fy6p4mmxYxR/ELwwgtCQWEPoswn0gSnVw1zvR5AR5cV3Wv6Eq1jH+v8SWbzUIncZucV
Bp5BQcR8pQ9DUd/8TYCv9fWowcKFFPmCXVRIgA4wkdUD7+Ty/DMhRq9xiwJJtS0PDFtFryJuDAm2
ns0yKQzsMyQb/CvkWghzlORL3r367aNoCNNZwTvWBhYVIWFjQfA+cpIJitr2faoXb2L1IC2fogmB
DO6fb1vpi75PWu/YQa269/oNLn+IRCeaP7+0z+/ttSS0u8U+iaG3Ub7PiwMWv99UW95e+jUUGUeM
0j86jOKcurIKWo45Tuk9MsgdX41QrhzYlpTUGr6f0H2yJNDHBYmHn8HvI1HsJ6FDLnd/+kX3WQcR
PHVTV6IT56t7NS2uFdGu0ZJufrDwntCn4mJslqNoe8iqqAC7wwf7Bk4W/77bgEk78BPeZogwfmJu
0NteiqCktgq8NtjpJ8oI2wxwF6z4AhFfDwWRkdbw9ps8XRON1Q9/B9C1srB0ySUI+t9R5yANEOyw
p0AoS/CXXEcwVBpDo329QtARItFvwIc/WZVxG70OXINFqBXmDWqo9TNeVG5BWargSmkcpVohtQlA
iaEzqcD6itkthc/wKypiEeT97kby/sNQjtgdcjB/u5bvwJQL2IY/1s7uFbCoPOlIGW9tlfXG4QZJ
1YRrHYWvi+o/eE02WEvMdSVkzAy+c9PjUF3+gGUax0LXQVB5OB+CEUorlvrcIPvxWSORCf0D3NwT
SOEGYLNKwA798xANuFjHiYi7zkH/sXu8xrh/QwORXLxG+/GqJetikscZjhwnTpDOHpzu/tsF1KfE
6I3SNrYCcBTjluDcc0coAVimdarkMhpBo5qKvX6u+V3G1oYuR//qs5VPeUeorf73QkoKjDANAhAs
PlkSuZMSf3d5pj0lJGjn0wIi7cZNJj5ic42n2tfJvEhFjI/Kr+yLugTtfvUaFiVYPsXg6mulC2Hb
S3pZHqsbUOjoMwxM/bmpmkoAC2M451sa2UuLcU4ESRMXO+1t/Zdlv78mrkrVN7Ow/zT7lQsH2ZfH
ZJHJ6Eh5/CY6P4cRcE2nPsfKRtE1AoninBtXsuRvVD3/G4IkrKEM2vi4AJbccT8F0Cm82Ht6oFIR
xKCcZAOyq/CjNLi+oNmITZJE9nVdV1QagVIBU77E6l3M/Nt9F54KEfgTf/IEOlfwS1Pwv9S45CPd
F0Fm9/5Pmx47jXYEV2nI51kCcrSnYq4w0oEb8E7OKKIwxUxzI18ZZhcHJqqmoaCEEZmHF624N/kA
Vfb8ezUWUBr+AH5aia0wmT9aeYTYQvUXB0X9F7ZzlaAd3dPM/TX8kn7G+mzUyaKX4BCfbzq9guh6
Qr9hBfhy/3eWEQZ/QBlkN/qTYQw8sYzVhmdxwWzjppDXIPiXVRgCuCoNvts7rjsJC6dWkfddC5PY
BY0wKePeEYq/Vp7bRu9yjUbgt4US+YEHM9cddjxfjxyLjrHozXg8QaEsg3mPozZfUU6DtDHRYZfl
dfhFZnkhfbGxLPdfenLzKm7aFluDCEb3tdv9UpeGCXV38xeIe9uyY9gu1NkS1cCVrZ64l6vPkvW6
v0lMWjjzR0+pU30jExBbodMFWN5TuEHv7wOHasScG6pusljslspcZfivFwNyzmi2uDk+YgGXgykM
wcmQvbB91bs/5UdNp2hx2TtGA4yEel7zSBqXIm3ksaF8c13tARSmXFAOlPy3PYRrSa4//KoT473i
yiCfaRdWcoHZFmb3Z2Il46HfYwGZQyXYMDCaGr1sw4dPbMU0SJH08eHIqGp+/8hlsHh2OIawNwAf
41+KqgJRiCM/Ert4FFx+lfmXq0+OXjCBQZngCq0HDErbsbOQTbE2f1H7IgI1JCNHhslUL4W8RaCs
xzmYrkH7zcIoKFrEVD5ApZq4KTfl7goMpSzgygMDKEqWLHa8khiIRTwec7M0LSy7Gru929lpmQwA
FrfTZBFZmNieWOSkZUZvw8IUNFhjDHTpJgPta1tCOULp2PP7jRAZM3/kKn3nRc5hIymn4LJz2P9m
TUquAyXXzAtN200nGmqygJ14GiAm4XvVXnOxM2/Qj13KZNnZmZEw0zPhKd2gtmZ2uhqcnt7EWIbs
JlXMF4aMTC+kbKwZ/MPF5ug7l1unwgTCDLP1OlIPf3jjPrWG/m7/IgL+1Yyb0diNXYx4MywYwaOg
9qk7mGq/I71M9PaheaG6LGmsHmgLYObgX28Dv6vZdz8L2EUiTr5GTzJlhkoDpIn+1QIYzjS2a65o
0vyjFzmNU1xmJCzsKoHFR2l0+2ogM/3eWk2EsZqWVFAsFkulN6dynAW9TkYaiEjhAOMkoptqvUxW
thgRuhf4Nnw0IMoYolKb63+FvlCE4gzc6Fnj5q1aOde5sLEkHl09AZKt0PFcaayQSQoI7elfbiGl
8TDekn65rz/Z+xp2wGOXuSrSnGlv7U6UEXxp8WTAnTo7eVcKmVLk0KVBZdgCfLVEv0HZlARi/TXK
onzVn9RdcPcEShr7NgSoX/eyFZAjjwFgKiH6JfSHldlr4LNp+K69sKE8xV08p89ShJeg5nzgo45I
FjhNRg5p3S9cNJCqezE61qNGuOQStnMBbQxvIPppR9GfP722qDkGqD04L3zgZLe0NgPTEQh7m89q
xseFmZDlSYkbKKp198wnVJEC6zEaic0hpoh5/4hZ2uq5dksq5GNezslc9cHlx80SGhpChYrDZo4b
T66C+gsFalrMFM407H0viuo9SVSIzsudoov7RJxC90CEuntkOM/qvWODBUxwt1g7zWMqF3CMmqIx
rMYaq7SHOAvVKFb/ucPUInzzelKuR+MaC5MzzGinYZbp//NgiqI8xeLxbMOQA20Nzt9RbnwgZ5Gq
fwD2t2y5V5Mhb2a062tKc/lsuG/Y6JYu63OhGFOTyDMoljLaKAuXe9DdV4vTODz8APTDB0oH0vTy
zgNpRsihaIUCFvTwlL7LsnJOlqDv0PhDavrXiUbKPkPU3ato5SYd8pwI7nRsehgamNNLc5JbUP6x
O1VbckYjHGlTsCpzBE4QCxVd7ZHziJHIePY7SeGoI2BbzHt96sUQ33AJOrS/vn3O6BuljWAB366w
lE5ez4ZFmoXLpTNSHJm7pfygtTyoQU/k5pOEN4CxW9oAFQM2QbgfFLCgr3ooY1vT8Eq4sx7tkFoe
uy78h3gFAQmeg93J7LkECxti2auNsLavPrtI/VpmN7QgJZt71d2CWlMK5h3Tjj7MO6Zevr6dUbsb
QhqeTVdKI0HWLgtKB4Ehmby4TqXfBpsBFzMKSHQ452c96TuP8IFczrjGhrcV8WUhZ/d8f/JbP4if
uzmVQEBB81ausYLBVHkCiui5rnHxHZEZprF+yh/5qhQ6DRCLOfdsQmUgoy5G1mPve2TNts5h5B4d
1ETuwo5K0HGnxKRnMHSvITw6V4oTP0+/XdYl0E5Z+IuRFI7qhIlb8NonOeJDUKQoURwaqY6E7GAo
Q5LBC3nfw32eg00psFEbR8GZwfTfksD+ymNhMdo1n7gzQlmPF1i+Q5tWfEefJMIie5WnYlzXpJaO
4YfXkMLS4KHy8zkg9r3AXb3orsKKJc8mDguACZYe3zzn6wVgs0xQf//i15xNFIrdDm6y0KQstYe5
0kIqyaZ3qMLk0Wecbm0PT0n5EByBix7NCc/jwh0Q3N6reeJHm30xq7MShVxbz2KX2LRMAJ+/Skc0
OF/FTVFECKa4kSN9gdSEuRqPBlGWIEVZ/DVmXuzNw6sZONWrrlDJJ2Yy1eQqJLDQnERhusrm7IDP
YTlaeE+/67LwmGlkl0ljNGiMMWhMSdQN95hhdv4e83QGHy3DWTwJ9OFqWr26SisdC56wDC/9Hufm
Q3gUNCDDK1psn6qSwRL0cTjwNARKJr0UbJAuhX4gKYqt8oVQPAFE1BTcw3uzl49tWU12uh4Zjra/
7U6k3xohcPP2/niXKoXjvIoHGvmwNXLErjVBiyy9RkZv7WeQHxR4/s/LTy+z5l+qIBxDyzQ5L7Ff
6mL/TvknbCs+fI2OXkS3+G7qbE67GLkFc5QYKQlLvEjUfyv+cpPpb0XvRU/G09+HkiL6qN/Fwf09
C10/1yWUVN+bWpN5S1ZKyWnXEHMXDVliU2GZqWkzv1bi4oHUo3XXFRFRYSaTofbCWBuMlZ2Yc6i+
bpyTenoMo+n428cKFwqS7Q+dnxrRoyxn0fwx/6C6j7/Lb+JiPFo/zq+IFSl3XM4GQav+CpAcbhFs
Hs5drGokE3sbmjI4SqotPjxWSSyk36v3h3F5gbd4JEdp3x2knx/fA53OImHlxWXQAe0JT9nWA2Q3
1eX9K6x/81M161aXt9h3LMD4jiBL+lu590ZDK2cUF++wgSDesBdx0xC2oqrSNs/8hxrdEuFMX3jD
GlOoZzUjwma38i6jgO1EOA6e2Cony+TUC6MbA0qbo1PB4Rzz0tJmVLDdOFqcBqHxm70tJH9Cz8uG
4v57LAS2OPxqPChnHHKresNTdirjK8JlKkpE3mqR+QNgfct4yaboPZqClJKQoUlp/V5TOo1IquDj
eEwtWEMYlBGZHvfWVFyEUZLY53yxSVx7NIXMHK7OQ+y+IC0MuS4h0CFHofbyHzXZ4osdrw67tfCq
IIdXRyj4L+X8CYjWF2C/WHLk3yATgoa+EyxnAXOpCa11zRIHo5+Lfh0vsle0CfCtxHhc9VU3FsjM
ALHopvqPqevuaSw959cf9c5jNqc5EALdEodNZTYIPqQ6wNz/FD2A+Jgf2kfFr4pQOAWc5vRMRUuG
TpmGxakMa1flBPBUH9sj4E+g4h46apWndyt2Anpd0Ee7C/f2B1ROo9Jfco55HLXbIVam8hMVbmzH
DBkvneMII6GiVw8VStX8LYy2873cOWRJitOoNKr5sgGdeeQV0UHeJuFuWZuTkZ6sIgO56wfwd9ah
Ps3Z83qCsXaa0NQToDziCkSHA4iTOsHbLjNN8Stw5rkPYOleJsdfqqHciRcRLbOBF1/kKPTsERSD
/dASrxFF/lmAmOrdCBMKrKMzkX1PeYbaLiJOsqvtJzPnhal/70yR+6jUEkorkGVmtiOEZ6/kRQkh
PhWlSCFil3QJHi/mNS0k8eO+Rp1+4d8DjphpNYINfewDxrbRHjcu/7RM/nzSM2LClWEXVJ/E6c5g
e2bnuWKOFbhc4xv8DuIqlnAIskWrr5HEKfwbpthot6EFlnQxNSdpqxW3kByqDqczQRDXVpmG4Tzt
DseAOyCyc47axm1XFGGPrb6xcDEiNZtagokAgP/HJvl62Ctv2S3ZcOy46PbvKUZii6tEOSywO0DK
Ns+bkwuMSG82I5ssbmAQgKws4RtidEQKNW+rC6nUaXaI9KdnuZpK6r5KzLz70cnYZiDUL/60I3oc
WLY5CmhlFTii6fnXYOH+dsLVhq6xQZ24pfpXFxbBwiX8602lPywIFJh8GmH1ZGPDaynwhO+rILZ0
VhSvPS8pS9B95J9pyIOD5Bcbwguak1Y2/JDEUHcYk7pf8JFuQwika4IfmWI88dyAUkzT1qZtK7WC
FhWoyCQFrItfPNfH63x872k/bd5HN+1rn1fJcNng5hXZJZIqSJj2uiG8cTWsy3TkzuJIzEkTAKFR
aYYu6cnpANzH/95t/+sdz7o2wK2c4fbQludp3TnWlRoirb1N9ILqJC1wEfGLJEP8dZyWDLmNeRVB
ckvDZWvOFqgWzECmcrHbLZKmg3wuY4mUycUtPNiXiWYjaaptztxqPYaIPM4W+nXTmG7Kg0TZ85ST
OXE868mXosYuW6MjXSfObfxn1RJ5QXCAb+SYplmLvAdbLAufXiOnkTHG2ajGTQujYoCzjEZ04TWy
jYN/Q56bW8Pkz62WFzNExGeW5VZMBcWmUx95sMf5ptCmd5YOYreL6ZHa4N++iMZOYzZamI9U3Gc6
X88j/JsBTuqLNDMrxbemkGUQjvwEzrEBKpL3/RbJhnl5yNZOsRCUqD4t9OJ05Nrov5lJGWZBXfow
D968mzDhGg48Lkqf2uyKMxH0GwiTy51y2hL3AjfpbkWn0rajIFBTrPwauSdIYT+t4TQQe8PrH6/X
tWq9/Xr2hqxf5ToBkSkekJtVFqA8i5Wm311zqY4Zdt78vlKDe4SkkIBUhmJ2qJbRvGHlHakX15Wy
uaenwA3do845mHo/ZVo88139w40o0zp/QNfIBEJoNk1tQVM2T3W4YwlwtgXHP8k4V9ne6s+4nNGM
XmZ5iLTme3nrCJhPjN8L3scI5yovFwfDbwugi6Xz0rsF1AcbwbpLnqjNYfSk0/WP8ZfEh82lE13I
1evt5hhiRo4zUP98d5Ry4SIQYdVJFOpRl/V2tBimM70rb7Iws0u5VVSAyFp+hBIk8sIJ9xDzoOv+
K/3Z/MxSDlpyz9Q48rDd1xfu2G1azng6Vb3mirXi4UBRCQPAIYHVBZGbWj8IDuV3DXYKPT/PSn+3
+dmk8kJREFBRbTQpdze/FGEGUAfaHlle9mnoOvbHi16xTcuzm3kusb9tPE24j5tqNmnAMH4tMO6R
Cc4AXq8s+07bG68gPta2yxveypid1aYuzNzneheqCdVV3zQrsrlj7ejHo58upAV38WkPbZeOca6k
qvu/dorEZ/XDsdRMU3dT7X5ZsiHCmhLqPMjRVUMj+w1ZVC2zvkKmiAZWQe1P++WJHEYnd0zZLxZ8
XbY1nXEeAP49PcB2ECI5H4nZDbGRu+4zUVxoW6tHVKdqs19eMYzaFu7nJQ6l6ugZCadtaOZx2/hU
ix/oYR+tP88cq5Mh1f3UI0wXq766O878uP4+9MMjEcwrzFFgz+70/A2sjIBJXpANstI+cWz2JlZL
yNxGSCY98yGQxrEcCWrapNu2HQLDuhkEGbA+Q9iB1Gtbwu7N2ly83plfDhMR5Rv79b0TpmzJzVRS
QfXDUVlX+G5Kdu/ITPsnk6O3+H0si1rWiNe6HAiEHy0aZQTfzmRsWOoVAdbhZ3VTW94vaN3a+ddq
2dIxZjntL/KoNSiUQLmpFDtJndCuNtYW0LFqHDrol6yC5HLJh4A0dxBcP9wP+ojcXLxmyTHyp0WB
EcndhfpUxLX/fV1dxHEfbv+XRbgMJz9hOkj0FoRR54w0/XMXgF4ClhRO9H6POpvOh9NLf+b+6mrY
w6mPKyIFGXI9DHV2DoLbZjf8etaM/dh6syxmGBwxQHqvDG8ELk8EPq/1OG1yu4S7wNZnupiFGevS
H0WSVE3TXAnxtBjdIo7HjY8weiDa5tmMzzbEpbrAWYozj2ajNdI2kOzBWqUeQZqFwgG77BBKw/GC
lE2c980CLxYZA1aUGk9TzaMCRKNWwIukeymS+KHkrAKtsqjYRT5Lt8mAahcZT4JfPVkAN8qgYci3
kvD8uuWB+qc4+ol6t4RQ4mEEsGk7Ym9coV5Iz/5Rn/LqT0lPkDDt1rAWexBB0jmwzg4eNLlRzT+Q
VivG3Ssbqo85UZU13dlxEXwY40T8ghUG9IfcgvS2yRKXP3ItuG3t7RSWkNUKk671a3iFB94Qy0Vt
Yu2rg2ok7Ng2Gp8iT47q2J6lWDFPVB5PYG82Us0cH+bqHhWOEZYorzMts7eqYF//HdsdTtT5paow
c4G4S77Qh2oS3zefYTgTO2Pv9baamG9GiyMRRpnIx+ZMkwvvn/cyRVuvEGyMQ5rdZRz/J4naYlr5
jdAnSNYCvXyBoWpiPYwOWXVHMfX2qywbjuHZzWuLGGguwr4vK6tRJP2YFLfsvynTpKw00M54JcLp
DkXcctZhXnC7Obq7Y6pu4Luw57B8gyspZmzucGvc0LNlszIT/xI6vSDY3Gi2SiN8LIf6GQjI3OSz
1SWaYg/Z+8p6uTFOfL6H31X/sKgc24ctztHYP3qKQAWJRkpolZk8NC0j1cwg8xJdKN6fMV0xRw/b
Oh6MvHkdvAPaOQThYx0t0MS3US4w85NRGuHFd2UAgK3VBfZZcAgCf1cwxipWn/nkuDwflGVEE7FW
ct6/MIbIIsROAZUC5Ipj3AuQpUhlH7H01t12IP62IKsxav9QlKvMd5x/eFTZqE+ontxbrZjPwR/E
OKZlVl884sTn3CVIMbpYQADO1PqQeZqTL6TaEFnCLBIdezcvIgJeUZ0BeLN7mO2eZkfVcWq5XmD7
kMIEz37o2yCngr5OPsg0TAFXaiC4QuXWlZerYSqJN4Nn0lIzzGQXuhXkvslPlahUjhV+VhABLnbr
qb0g1FGbBNl+Ufv8yFLmXw3BlHcBq+GYr60Ic053sPTKj0wyphjVgf8Fu8yeZCzdptm2JzSrulUE
iRafKFQJ0QsbRrb3Hi9gl/p9p0fnjraRjihb/5NbbdHrRg8+8TQ8JSGshFfz1I+e06dLyufc+618
y/o6USZ20LvTmF6CfdPNIIZQ27dudViGY4HDOy1CZXtMdow7S+lnPNq/QmBiw8LQolDbFFdqFPS/
kC1MFgF1/iQDV2t5288n7Vv0jPbRE8dG2xWU5mniMqW18bCDgxh2DtWIJydpYjWAbhPYNmpJRQ6W
hA6Us54TuVD1fDRKK6SXS853n4nIf/s0M4K/m+SVH3bqPKJoqXlPcXJcdhGxZoPSELiunkEmd+v8
oG0akQ7ybyqm6S1q+6AxVuNpsjGVfSS9xrpMi2X6kWkwoUFu87rSeHhrUfkutV+ne6yA/VFJvG+q
Nobx8pXOgmOjqCTQrtoziSL5Fpw5OZ0QiIj2tv/g2koDdvFDWrw/PJxl0hJDnEeLDUaGxQO9B9F3
/iDHtpBapTm870zZshhxAiWbGqYL/Ml8qPDwao6KKGs6OQtkamTQh3hsXBac9C2EPOnoMVURlXoj
8fjyRD5BRge/r6IEwHnpFi1k0celk0ET4jgSxBrVf0sRBEq/OHyEsiScDXJMBMCsHsAYTLmIZOhp
4piQwhixRsKDFHrktLFKtxHiCwIhh6jODS0Dn4CyUwC8wsdbNaeXTlWOlnXy0HVowXYfaGxc67Yf
4kRFU5WOwUjC43VrO2e6rkmAiaa5kW4za70J4qjZQ9lx/ORhOluc49c33N7XiTZGyUnDlY2yNi+1
RYptvFIbGeWzSK2MISljiVTbB4h7B6V2G+KJOsYuEU80Y5BSGDg5wSA4524K9b0SRL2c9rUrw98w
G710pUs29sAKiViuodEbr/F4R+/jvz+KkYy3FoM185vUMjQGtak7riy5A8AO6amdxI7lTDo5p+JD
dSRImDIoKYGIbgJGwBY2cnE8uWVZEErG3yO4mH07qVBGfoloHTumjrdELG1QpBg/PMXObTk9ZJfY
5BoKC0SldVb4bwIcuJ1IldNLThS6EBDCR/GBjNe8C5ndkb2xXeAbgbqqIpZ2dp/xoZ9tiojas79m
3qBBfO4cDj41WtYOKnKYWbaHGzeDdOY+ARHBfSHTTPvHt9Pn0ggzEP2nlGmtnH/fEO1LIsY3bmnu
RsVPkw4vvdOyXp7OwGEDG+Ieq7lmVXcH+myRwDKfSb76WXscEXFhrWk9r4mqjIwgFyBXVhb3fmma
EOg22jEcQbNIG6WMZQ9TlFBjeeRm7ceV+jWFLKxgw3RHOb/jpqi0vYH6mBMv5onHroiPQJ0PqUfV
Ctk6h5CQ4Xi76pn/ssGFS2Legp9ecPOKentpgB9FVVxcP8UTl937MFdYREBsFSuF/hDX30Nk3s4b
CsThE8JYmPB2eAcjxKPVjm5sxEmQxiz4cNINBzDeIcIthU/mQHrvUq6HKTQJNc3ezybiCBYDJdm6
V2cT/lSfPC9dsqGoXMWbH69mPRaVL9YcAU4WvTRofS73zVgwtvWMKCHuf720TAx9Y/BbVOGE96om
VBZxsFBJG4P1YSrlLxdGRAA+B4cZag9HINaoULDgcwn94mIS0617OrmyPJJV4AF9/FEkgfrD03uQ
QosmunKl4+MA1SUekd/VYzanUmX7mTjOCbYjT4twyQ1GuuTkxZHTXEuJ0hOJlMS7HK797X1Bjb0+
ryhy2fAgvtF/3zCe6+LdiFepnZQTz/wKpZ1xzq+9XF5XyJ2TD53frDBIdyxepD4Jn1sUXfdJ2RRq
TWFJFyWBZpKCHdyp47dZcGcp8q5jL6LGIsoAmoA0zn5Cp80BrHU5bBQ4cELvZaHjVc98c8s26h6P
ns+bXWc26Sxn0yJeWKBfx/AiU0KngU/Gu+apl/+XhVHxlpogrmYq3AZipldsbMAeI6eDnHqsBDSw
obI92XMXs3epgMc2JgcJ01DqIFkV9KLD+CK6TTnZy1XN8xWTkBl1iKrUmMw8fR26hGe4ysORd2Im
AlY2DKm+N6s8PFpbY19cbae1IRZ+3w40WDjezGGOHv+t6kNABRm8NDbltoX+D8cSSyKIowSSND0e
T/echsowzMPHBR5ezoO2w2DELF7iVQ7PlTOMHn6YKaZdb2j9tHdSphapUjKnttMEKq/GbrfIkaKz
hOE6raWcBH/xLGNZ26obMKPDwYYkvC7XG0QRvMoDEm8Ao7h1dQ7XCrh+13aS59k/fHs0knl2D83T
BQe8FlcMYlsj2QbYX9o1Zrftg81JbQm8i1OA+As/08Bc3SkwmDQW2L1Y7mtJBISgKKWyoJIcqFZx
u+GcFe2e+4TTq4bSq6bJQ/VJxuOU4CZF2/VVm7u9TmkxOz6B1qlKlP2s0h4f+cx6p+sABXQFoboO
QujPiMjPcnE12Gci6ekIn1t2y6mkj/5smd1aYJd9dQEhQfM4oBg5+AU+26a4qfcs+HDfOjz0M7j7
ZZOzO7O9OMIT2YM+0FmZh7qHaQ24R8me6oMg+JYa7hJ29EHh1/M4J76PBrubh5U91+U6KN7ksjs8
alU+ZF8lPj3rQDSCxlk32e57UDJVAs2Pd5kD1Jltsi67MqdEBU40+lj2s2jbH133Dmfqp1sgbzx/
VFQt2t/5zTCzALdKwGFG4hlqY/CfBekaAwmq0IuC+VdeM6VVHIejuA0G45JMm+rJPxjbN9Ip4bVy
PbES4NHGychir6S2+iId33nZ4vxYuhk83/lb5QFRbySdcUESBU8cWOBq8NHOlH/4YldHu1TVp8GF
IG7lyrQ8T2G4Xo1wEyV1ANzydnNeJnFhG97RX8snZASwklvihOjXRuYnbT4A5Cs2Yo4O0e0NTh/l
Hs60gi6npJck5aQUY4x5zMXKWwilRt3P2fpgMa7iebESCF4J5xpuncT8o3tY+MY8wGnAQnQH4ej9
X4cFRYrG+lfhB88yc22e+dRZ5Bi5bezTiu+iixViIgYJbBwo16luqk6yS553KbJ13Ueyukw0QXXm
/Yxx2nwC5E3USzkaJAakohh7ynN6241+kA5BWlJVGAuYDhDsTU/tCaitWgzIIQNR6VvNDv+zGhIB
A3SJy9ZYlRBMbXDyxDj/ojQ99dXN0dqCWYlXoF5m/GYogiYD8NXbRLLLQ2gyuzyxjBNicrsTk7SH
Ho8bh3upA5oTs9DYUF0vLuz7Q52MBl8w5BvvdxGsGeCTegzRm8vKIEX+5BJToVfqDJb1gU7s9huw
Pc5MVFrzLwRJWr9NWbGqywGtRlJ6TiRvm6bzuy9dptD/FZBjOhdDczeWlgVV66GTWj7mydYjNHL3
sCNPCltmBwUNPAPXDzRz7oPzo5ZxRva1TMrEhNNdHK4VYMGBws1EWnsLO+dPy+Ax/Hy6bkaTKXdr
fm0Sb+c1fbjiFHjgwLkApZELBqfPc2GYHPFjyqTROjfeO23kRh3U30DlWsZGzlbjefEpLvCe8SXH
Bty6uf24VOifsMFCndAFf4JFEfxToLT5KQV6DR5rroA/tzuLWBaEQWHD7rfSqA2bx2WtY9RnubR3
0FMxyMybKb/NNwwNswMr0/JNT8iNzTG0Q7MwtFQ1vO7XulHKSVlk5boFBNyMZu5AFsFEHBK2cLO4
vY4+wBRJOpFw2oDXEYUcLGrfiv+tpIMtGosukXVZ2gTDJPwnri0HLXhDvXHMHCFLZIwXBK1P+hJs
dWkrVy5n2MePFMojk9hkqXh3Q12vSkQz1KiPKaiDI96bYr/wcZ+4o3uHeDKR/aMwp2pF0dcEQDyR
gGWYuZ51imR4haYsuCUWI+caFPOVY2EBZrCjP9glYsZkPUKSb47kUlBp/l/XZHOj90sjCOCWIrGO
mSyc9j+DSWEPmsnHgDE+funVsdeHGfyZpUzqozODeA+qsVn+Ot2KvV9QxBL/WRtIq798AJJrdCyp
dQ7FpKhYWvc+A2Y0iB/BF+KZsv2W+Uwj2G7Gzq0ZGliJX06cY9k/9/teaRiSFRlu9PoTPnh1JoiG
AKsDtYZJsReRCj0OcX88TBfRgdCzggqA1zGtjcC9UUWL6RBiP8YBqxdXRNJKW7UQby8we+xoS2+X
dmaHD7Ea44Na7QkLuSQkBobHYE2AsPFHZ7Vk62kPw4vqt/p5zYzbrawdlr5wB6oDCpljsl7OeLoZ
dEbFdXc95h4GKbE+iP+AkNwao7GL2gm2eYfiGFTJiBMcMVa/HRksDeqB8ClsvTYl+gq1OazRE4Dv
PKdMGPjnVXJriNxGRsmjtPS9HVDYNhHTKd9D8kdmwfT+8/RWERsgo9BtiSqyQBoXDYblAQSpop0Z
zgfCxDLqURCBLa094Q1gGbckT20gm7W5oFdfk0v5nhABCLxdfjeRxgCrwKLRLgMxtw2kbS604NbO
4BMasbJX3v7ZKRdivQyrpfSMXTFj2JJ2wqVh0paFifF+5QvpktydaburlrP1eFU+XBOcHQvfj1DL
xefab0/EO7+KxgfL2cRprks1ocjIaUuswrWUrmK3aksFQoBbUfuisOyuamy/8Wx60r1n8x/idznK
MMFNIs4+MyLjKFyk2YHoDsgRNzLmyvZpqtzG6VWcnP61XvA09szkmRGpEV8j7xw79u/AnHjLlbxq
l5sVdOV11D+2zde0VEozMuA3JZ0uxz6QYjJskF5R6AW9u7Vnek8iiX5Uesm4GR7LEc+ifBjqEmKW
sDSz/x3SQMzNPg4QjTVHMklPTUURVvCEE1uGRdU/w7rL5M/vCnoxpNfIxGgr7+SwGADbCsqPEU6o
DyhHQmiX6j0EuL8cVX2Z0HvHUCT1z3siWKUReqH8GwYH6vExSEbKtsTkN3bBJChBnGf33OKxuvZn
qDvUKvD2m7Rj+45aaTil1gKeo4O2NzNQlIQs88CcFxqz2PKFSBAuXanHGlL6LGh7rUDWqZ9tF2g0
o3YpKIbupXv52A1aadU9GNlxSzjCaYkOM/4Hrf9yQGgwtVzyb1PwE9QiDtpu1rgdy95nnryp1O4K
zNDMV1/LC8Glq5TorG1yo9g+PdW0X7SK6DMhr4WKpeaCmrPej7+LBdIqHjKYYfFbVP2R+yd8dZ9O
48Omv1/RFJejWGiI9F8eDxAqrpPQPplLbCRWzg+cQJ+4gT5SWdV1vakA8xtlIH/Sv4WOnVsg0YEt
4XEf4YkACaRwFg2z7iq+oSR7Qz1EKtM5Q5vVcXRSARvam9QWc35Xw5hXMsyeH03upX4cMBjZ8JRV
mnyjz821EqRvcsuKU6w1ueTJuxggOzOQCztYuZbeJ6buK2dKHGE5ehx5nWhe4S+I8CKtJjbuEtZi
SjpC5jEePG/YdRyhsBrVXXB3N5t0DFAfuZ7zIXCWlw/GKY4eF4NwIz4lk5ObroSSC8hLlbRsPWec
hH5A8bElIDZWd0SpkD4Nst1F214Ngl08bf2hqjcct32iK7c5CS5+GEJ03u/0gBrpvv4aPoLnRmu8
oVW1ZFapIyxpWnOJ9Lp7St+qVK6GqCqfptCSxHeAhi/f/i67cK6JCs5/VpUYvXMBmK+byoDZ0Jsn
rXLKxnAKr9l1RNVi8yQobvJlf7IaNxs6EPa02VQSPKs5/IITwvYpJjmuSHgY2u2WlrsOCTYO7ptG
Gumn4LJn5IXw77azMNZxadAr+9fw9ZF6WVJq+HQjDaH/fZENXHIyfKwABc4h7hoxO3pBzHj952DO
eK507YLEJhaKHlnFYMvefbyJvHVfUd3JFOOcIJucpIjRS3QcpkKTsvg19viYVvT1xeoqg3+eZfgy
G+5G5Nw2KhUBbY0iFYDqT4at4SbGacflGq/GeOaBZplPiKR9MW8/kAnuYIbFMSW6gmotCy/6oC+X
7ejbcocF8sOW6MQBv257VJjjUxd82HXmkMgtkh/FKFGGbuvtayWM8CBYv+tWzXFLfW/SouopSjM0
dXngsi6wuDe1cAaNFbrHrhQGsCSI+ZqKF+Ms8R7nHx4clrBMWj7WZPhCrvLkn3vQV1oRlZWAtToq
CXu4mBCLYbs3tQhHw9vDiyoYrxpHoSUhOr1akm0argQrNWk/zH7Ic3LpBamWI2oKCbvMM2pB18P1
pxvgs6UkwW4pMddi4aURo/ogFORon3AUzdZybpm90iFTr19stTXBNdtmAg5mHZ22gm2NflGTjbPC
R9QP8W+7sQgL+4HHmCNrZZ4FNeBwngavCgcY1vE6bDTpSJPeSJywnCMAM6mMABYsrVTw/LaKSTpw
thp48FU6OZfX7oNFSYLQgmIb8C8DwCn5A1zSWyit93Zx6h2MkFQBO28j90ZZG/gkmxLEtlvVmUFu
XwH+RKwAWL2HO1qZfAUKw0XRK5sVGDiFmvIiYab1ljEjcj0qSDJLZomz66njgdBJAggluf5CWEN1
so4ZIcES2T9sOzRrnPtnnZR2leoIXTMslKnDGFlt7a9dHzyqtgbPjmdwQnwldoY4sJT6kGwIj4Hm
lwPPhkHAHFcr7Nm+PcLPjXnhrx4bkYeJFhD4zmyEh6Ifo72WU4KA742s4xzY3B9ho0RwAc81hIkk
fBVgEiJXggp3a321NJZ24q/Nk8ewqrBrQv86etXtXaKwD7peKeJKABtszkK1yj/2VqKxggmdnXQL
H53OW7zouctt4mAHSZFFDo6hQkDQQbFYqeGJdnmHTqXhe31kL9gZmcDzz3jbOEr/FFIZuoHWA5xk
0E7V9ONPzxJikcwS4K+rm2j0c5KOI+noEbKNiURicC1U1eS4YjF3M0do6SA5r1CQjPbAnf6C1Lbk
UqxYMz2ysyumwn7sfOnDBQOhNa8qQF6lsF4lv5KjybzEkS35J0n1i9+vj4ceKnknKORZEgckAMh0
Qcfb0ErbWk/lveeNi6wQkJSfZPS94X10dKYymLlQZ+AcxQw8tq30WW2qrPuNKIan58rfF2WsNt2V
UhmBJhO115Lt1vLQ761tGt1v4O1WPn3Rjrg3y0g7SkgPnP/wQN0nuHmIwgvAcpJXhiBGxWeVv7Qi
goAk03uiLvEkzAomqs53Xevy7I9Z72k/DLt/RhvTQg9WuyuFJNO7fTj1dUCjc0qlCk+Ti6wtkbTQ
uEREYxANi2AsKnp9kM/vSWZFV696+lpIqydYQFmxOX8hqxFQomhFrmhwRpZ2CTNYRYcOUJbbgpOz
Y3HbjpUuuovav3Yp9mDHmtjF6tkJGkl8zNENcU9KgeGYEnPbb6JQg39tsTM4U0RBfrSA4mjDBzNe
n3NVNzfdn2VXsqDSxhni2zGhjBvp+X+ca6qY+UENmgZuOYYkQaatwDjJhWzCDaeGHWjmkhYDTAmM
AYTfD/Do92jNA6c0IpZZp7Qg1FOA7sOwL22sHHEQapfij4YMU6rtEYGjykisGlrOCSh/6PBAjFBr
U+A4ouDwS5eiRscgvHmuCQg+/lLadLExBvX0Nn+h96MDETYLt5J66ANPCSOn3jObQ3jGlWhvrigm
B/tMkp8wZXdVnvF3NgriM6JI7h2PpqPimugfhhUDEmUwKkktLZ9zfCESGPuMOTUXoPvbZ4K0o5sS
A4u3mQI0WnAs21Sbih8qRTNhnXxOx2ywdgzn7LPk/CbQarAxzOuFdUJv9TbWcRUAoqy4S/W6EW7Y
lYypQPopSqNMlqnbdrcdWlVbPdDMuXFNDN4dijn53Ey1xsF4RYCBLgYVjfHDMMu8eEsA2lFXTmS8
038kkiRoGftYA+cPq5yJPOoR1L6ISh5BuB6zkzpaAlij2DvUDDMjuEbRf++BAgy+sGE/821A/Gf3
B4TJD3OhVjMDfel4C0HT/Bs3CpvP5yG//ihBCMAhczVfBwO5Z8yz5F2CctKuDrq0bLHqD1U7q2lt
N1HSFn+T+3gLtUU5KJWYQiD1/18QPxjOuKGgXIioOlkUriY5huJ4lluekLklHrg/i4Xbx8E1ZdI7
xv3PzjVYXv+5uHzE/oOE/DccWzn7aNvOiB+tbu7K/Y5tjf6lRuWhIoGbLMxnIEwS382ERXyFHUEz
TFCQmV8aBubtXnqpImY0cf2buRFpLIg/mdRoTyln/O1KxoyfJMKr/AGCvwt2Yj4VVKA3Y+mn0991
cT/ZnmD6UtekNS9lHpKxNYQGexdr7gR80qbPApNduuqwlLMTm13GlKREMxbhDyEiUVYyIGsvjEkG
1Dx7KRb7xaLjL3EHbpI91gz9KGviylgXhip9iv6RrGw9lLDMOXLQExBBIR9ch4HlKM3N3U0UgTwu
oCFLvOkiKFImzIT5NQ5XZpN6+NyP/qwtEZ6mS62FrLDqetM9sVokBtHzZHM14Ct2bGvhobNooqNv
LTBOsy85TOGIJ1Oc2X1B0WQRRpGVHw++eowHWr6e7WlDKXAKdbQLS2yYWGgJP6qO41jCjom5lKGl
UPM9SZIi86BERl+p6KkRJZeWjajz/ZjNWwJhEeyXId8FQSwXlG6qhBrc5rUM0oRYLKbFIELegtSX
gzT0tMI96H2DEEMpP3KLa3NIbVvRSOP/ThR17Bvys2yzAiVAbOZoNysf6mi9aVjJyBgAVuIabZxe
xtEci7zSWmP9kcuPGWcG5YVRqp56CAqd7qge7wgJBpMc/pczdsn/JsXBgmnoXWVxOVMxJfdjrKPy
bFgwfNwuX1GTJNcKoHniGaJAHGCVQjm0CPfimGh22+yRgRnKb1+fCLu0s2aj5WKK3bfk/iWisj3N
9g5ET3OlHKQUxx9pTU+qWxonJIrapF8VUPcl60Mc0wXcZUgSFUNZHMMzc0nFKPlmpXBZj2qn94ua
JV2Id+zr3DGVluRVhomapOkCZ7s1ZUMewG3D7/qhxXaqbjAd9cfj/n1XqWyAwj0o6mNbFz6g/7pP
4KcJppOS1/+mZ3RIsHuBI6gcDwNd5+1yDWjujQrnQGhn2jPCOdNcVecNbwOjxIAoFeZhHk5jL9RJ
hpDTTGPoPu1p/dO3UWEhboFxlhNLB8gJLW+NWrE1Jp2qbW7hWlUBpLkVoMWCJyeL+3NtIQ0DSx+d
WEeyd5hfy3JqRxusmMFHAQR2MbocLoZmWHg0C2EfgKUfI9Xhk5s0GwSTWqeRvBdqh4AQinKmYVUT
9MltxZR0AEPKM71aE4CGRpkCEdGw2vD3Ya6PYwqoaGQ5prW0EnunzK4rqFymciQOBvbwNV/1H23d
jc63jaMoc4t4MPOBhhVPpI1gfleASiKwMtWhJDgiuhoBdU0+RMQRT1sQxK3hVn3avu5nPU09fPzd
hrbRZYqYtel4met/lKUmGCfDAQwYhJarJPELheMVLJ4unxh7n9Up4XAaVjJWb0rHPQYab/vkqI5l
WtoKmtHPMYYMKRe0hqDqYtWUNvvODw7CJMEMR6Gtq7Bqf2Xgk4JETE84Ih7FL8sAcBo9D6arBCHz
bMBCwX/iKj870ZJ8YjaMybeylxuP8yuvKGGJDwJbgpiNMIWp0E01LwLFnLEjb1iCJzzfajrh/z0C
GlimUl+5gMVYtfFno88pSB/UrhRFNxP60qZmkxiKAcd0xcOzKI9KmF6d81BE4lxouFaPPEUftWVK
FIXipy7ihnkc/LckaNrIjHxgg470wnTHL/hJsI1fShIk8W5zALU0T9IG4y2U4wE9aRyU5IlYurRp
NobbE/EF/UFNnaMm2trGek/jUCTNxz9IZ75f6Qw8naKFL0jap8HPSWve9kj7lsE2fEzrxsDn4SIv
kEGbBPhKF+PtEduBizWZlDCmWLMIxAP9Is18FxssfusH6veFKuKKBb/ZBv/5WSidfCnGt9mJ5H7h
zxQxCvoi3g9CdOQ/4ZAkX5A1zjME240iZfnruymYxYcAAMz6oqrlZtXUm5+EeQEjFoSxpoBScLHR
Q7nEG+SP8cZQ7BOFIt72RDtvuW9H7Y9FUa1WFdJD+iuLNmvTvQ0ngAcg0n7wNgopL+Bu+FO0rnDj
WICc9rf2SpcA0DwDHVxaEM/NBv4VuN5DNRAt9QwzbpDtOQBslOKDgqUJ4ZqcK02Jrr+ezL7q17db
lUfcjKgkRhpJPC+Lcev9UOpvoLDSQ/LgcWLLp1s93XEFv+Ey3JHodWRFREnen5w9FjU0MhVeUB7X
z+iIR1VLhNqWbigq7NQqN72qtPv7YhMknRpD6NiVT7YPG7NkNiivfJ2DwGN68AQXlOssXoiM3H0v
S36eiYgqhVT5+zZyeYNYbo8TDGtNxSUoXyMyRIBsf6pki/nsX6xijS7M8765ZhvwtvJ+U5xwT84k
p6/UbVDaeGvDNvAS5P2KjgxtYfDrYVcZoPGqyUy6w/43Rx1pAl4GwQLV0um+pwhn2iYAgJfINdsM
4TnFkahPVy2P3O4XZr0ezxc2le5bkOgb9Gy3Yu6iDHV9cpo0nlTBAx4KTB1d7wWtWNBaz3Fj9e+s
U0WB3BkDOSefEbSzWOd+lmOO191TF7cskJ8ddLW1K3zmqfLe+ld2j7cupTgzLGY8E6/x8QReNzWY
ed9+RyhqJxb4oUWt2VTQKsJq8bodF0rsrdy+NfjsAZ0ffH7uRuwUlYey2wByYINPY3o61DjqgbjO
MkNPcGA6V8s/vw+E4t3SBhgBQh/rQ0XHe7EFHM+k0wwfDZkXPBfDTQQebzs1rHx5zXxp6ZTw0DOl
w94PgVsBEpqAV4tZdr3i7bz/YCv5ONNFjwM/onUm0rUAXI25BR/qYcERcWXRIOE4DNVBlI4zwN6j
KdOzcrnQr9L/n2wpU+vxYeCgPSO0Pg1JwpOAvKLfKKtvqk+B0TeQOlkElTUPrc6G2LnkCXCApqY8
oIsLJjNKkFkBgKC/R6/2tkHMjLrDd1/bVUkr91qVlshBhQsmB8szcUGM7vnOrXzawns5uQRAUdrw
2eA8t9CyN79CSJs0X2jvkxwsuSfueLuvNlstmvvAOJwxEcZCxuSvh6nfgwlB0FKZ2ZWwuNb1iucp
m/XFw96OacmF95mYxA0ffc64zhxC0R+G3OoardBX1MbCvgck7S73s+Dzeq4tGqkd2tSgvLpl2/cf
PtDpJAYIYb5YQz4WMrVgARPiItKgxfocKcIHU/4oG7uO5anr3AEp7kbx8pyz6KQTrkC2vGWtn+kg
Thc05EzbFjgxL9nzAFsolHf24YEZd+AaGlxkA5kpqxCn9HJxEK/9oLZZx5BgJvhsp+k4IKubEf9u
5CNRSabkkICK776U2OFnA+0g3awY5G10yrNwqwJLJudWtJqkNKWjmEZCIQYtQYKzLVwwK5fJk8fj
u1SleWLvF9/bAOuxwJHlLFQCdSMIUgQQ+0voQHVUcueFa43gRDDmdZxjX02jBNGZhpKeqCuUZTlZ
1jNn2NA3yeoPgaB+p0RAhmDlBEy26c0YderSEOztK125lQs2rcwRdZCWsBR20ID1h5WEPJvosCN1
rfTPO+Co4XBv6ZcRreedq00DLQXRemsX1ucF2Ujf9hgJ/gBQh1m9MS96Evgsj2HOkXVw/MwP+RjA
dCIdziDOWXPmf+cNo45xPm/S14oXoihiLqywv9y9aM/JnaNndCsVGVGM+Vx+bb1IzonLZKGxjkIX
3uO9iVlDqtX+Jj/u1PNFrH5xZ/OrRXEiPNbFxfQFya08LUL+W6iYu6EX1wNF+zdW3oTlzW1KsQ/6
r5noJ5hzbc2vpgpjMJ5poYr+hGNLPyTbdYc38h3sZrblpNU8dVOdi/cLDwl1uZIuCzfRIADh8kR5
+NbWuEZfDfhk3sD8xjo/6JZGoAnWvuqDOiZHbyyyfGL0n6xo3jlI4zZCQ7TBD4H2gsr3iYPmtNKz
iz59G4YKHutaQVleUSUOIiXt58ofJgLcLFKvVJVxmFwYDUIiA+AHVlstiN13wEgVEPpwoBexJK43
cfvRLhz0OtHOGINR7LqjDWnHmu5PWFru1ndZdrBeqHHEndtFr0/xD27cHEYT2locyd1reUiHjBqZ
uM80ZKAaxA9zpzwJDtEpL2sgx4LIFbizh5lWWww05mPIO3lgCXz7mCAYABpLgxqThRPSaNKv9lXN
h/mq/+5AC1udnaIJuhURZ8e85qi/NtNMJuNfH72ZWOQSvTPJ6PFfdJ58pIQVRtsFAuFzEoJGdltZ
U0da7G2HHcndRDV5TVuS2iVWSvlqJ7dNSzRf7N1l7RYSwLT9J6l/aAePrC4iyocOl9ab6tmoSaIt
IU0pE29AzPcHjhCBkBxiGThPkIjBRfIXoywM68Git+1/X9mr6cZbio8cFdYOZOSKod3eT++KpqDO
01yC+cUG9DUYvQXJxeWJeYV8Fpj5RFbkRR8u6DEVFr//g95begPeDXUmvDdXkeim1ImILIBtlfT5
mX/el7knDsLfp3HM4gp0wVaPnHCiQlLS44ZuPhbtpX88znVLKx13AfOaoQmn7AKJZg3qO/Gm+ka4
UW9erU+UhNIQZWMVhAL3e3kJz09E7YMCFRE8ftO0J2Ijk+SIGJSLpjZQwpyBZ3B6Trt7Dnvt/Yts
MKa2LDv2VqP8HMtwUneEVtThOM5Pnf5LctsNV96ACL+V2UzP/WuR3llL0l4Wc+DnQo12Ecqq54+C
fj9Y6mE80FTeZlZbyc9Cwi4iVVNDM6nDGXnxrzD6lYa2yub5z2n7M6xJmRx24FrBeS9CVRrYNDdB
1mal61gsN0/2UPxPegU1cxvlGfAt7S7Ax31hVlSC4Xk5CF+/UcwrLu/407mYQxS+FsgsM+tq6wsk
kHlG9ZPtXSlvmAyS04ot6iQE2p1LY2XrH11UY5gPreHLQBqjsx8dVc0FZVXKG3ypw3XUHOER22y7
yuC5LxTGi7Wl9ldgJwdwpp5El9gXUVnahYzxjVX0x50dP2g4RIFI82I0/F82RJsg+5V+9EYIZQ1j
VRCxoccZsgpUbvVk8TOzq/w4LEm+yfvyK2qkQPWO6IKOqR2cLdc/gGGezyBzAapFm8sgamT4olov
oFVyRQliukaoRx3eRfV9GzZqufJZQC02O6x0pF99WaogbpdzGPImK0TUiVBjkZFIPcUDAI+vczpU
vH2BCckcpwjlNnkuzETOQ5z9L2ZJaiFBYJ5zBfnlxn06EEEk1qZRQ5AsMbeokJxA1cek3wXIl3g/
wTlHcMjI1gKEntcluVti58viaJyqEV9HgGskTWJIyuHmLwZOZJ5jE7wzOAptxDJyngQV34Z1yUXm
iHsQIWK7g5RfhfGYvHlCYoegZUMvPNY+tgl3DQDopSxmZiCI6T7U8MAyNjPvZ8lSpsiwmt0RZJ7d
ctB87krMFx6wYgRoa2JgodTZMO4MtROpq5ciCIruXW4QC5HBe43I77NH9mdQygLYFSDesQTC/7iA
rzPgrBNh5G4nbpPYwXf8u2LH/7Xhe4jtB+q3sejwwFcsLccI2H25nR9/XhkH5hI10M3lnQSGiYNa
YYTNDHideqi3Ay/K84/fa3DJ4RrHjsEOYqFDqKCPH2anVDyBfXEHJVPAbhXI3vTFmL7XDonJGTgp
shS4yTS14YwatFfMhvCxdl4OWwib7N64KpERTlnW4a6xvizqU4u8NihIB/rfCX1cAcI6hNtbrF9l
j1zmL1EaNqLJ7uQoEB6cJw/7/0ebNPZLQUE+kmLBQQkDce70SJFvvfcNq16AAA980w8lO9YwkJiv
ntznh0vDLhMRdytrJc7dtaiNL1UTcrijq0vk4bOnDyYSIdxzO2eAiID3cUsTyHRBC+ZF1hAMYBc/
kVOy+A3TmJ5mkGrganKVRTI6BSKklI4tipZLmEIV4AhVjQd6okD83Hc58pWCXwFXZMRlHEP8CZI2
1gUURTwo1wEzICZCma/PdrgVYLxKRf00bDDOrVe7BZodPjopbpsR6WhEvcfiqhtzaC1oG+4A8vlu
pgjHmFa7/w7XsYCTOy9fiOKyUbuT4hS/kr+yhriiir1Q0x9sVV7nB0yUcbTGZvvhvGuZ811/ctHL
lQYOjnT6vGWCqtxzvOXefcv7l0gj6BU0A72p0H4lNWnfabT3JgK4LV1MMtIy3k6+fvYsyRIj0ee6
jpyAArWdGjpvh7AZRemuV0PqNWVeJJ4zx2f8Bi/HXXdUr0RsGr8oG3TLOdD5qlL+713me7lZtfIU
Wl6eHXqEsNa3Jza8Ew3+6NNpuyPtEqwMiHiJuRXW8Ktek94oKasUgYz/b+qsSkPLkvNcPleSFbVi
A2Seh1YtUiSya4bR5LrNTf0/kGmIEjH8+3YLpn5cIEMYTDu36EpIswS+6kSynz/JTpmgGLOWMUAN
yIBPAQ1TL418G0w/VHBXk48AX3wBK0NsJXcIwROSpF79bz7sRCu53AQFutdVNm8mjolw27xfjOuO
S22pNdmWHhuyXecegjZJCWRY7Me3FKn72DYLqaXB1xDmaLbKFlnds49n1kFDCg2xwEjqSGmP+14c
yPabVHPJqJnRsRCb3GbxwhMFKyZv9RZhFEDZNzt4++a5uiEggtmihaVC77ovSMJnt5zYW+CXrWgz
7iqd3oYu79uo+bEUITw63SnPmI4I8ClzE1Je2TOjunPJaokr3r13Jx5yOS7p7WxBR68Itj9QFrSQ
jZIgP2UOr+BQ3tWNxVXTIankLTwkXKUqW2bMD7qotSoDUb2x+LABaw+3/g0cT/y+Wt9tyw0vqpBk
OKJ7ps1TLVHL9FowWe5d58MTaLXjojkkE/BoGBWS5Qly/0ZMh5HnX2xjemlzTkeerMWSo1JZVzKD
oBLCrHR7OokqqGtb3om4BdjIiHO8BkJCjXOKfQGGf13ipgG41Qi3su+HUFvZkX4ZERZrWfa60mJo
84ugTmYjXf4px66Vf552MS7xVWv9gHCMyCilISWRzEfmT8DygpEd4TmuoqkqcBQTWNrhRbiZv79+
Bb2sFhZ+rsBc+FFy7rGqehHStqbE26Y5yqBVGoc8OO+mjkD70iGo0YuRaBXrTWm08vHC4FoX1hbG
RWORrY/F2vzRwbF/ujtHu9bPZIv08hDycc7u9aBhOk1GDUsLqd9IerQea+mM7+Kb5FmdDbTUtHEU
QPebBZdzishuevjCZKRd6sxmIEl/lfDfwa8Lum+5S4JLExr1lHQP49+UAz286PXII+W2aK0hnmuV
6GkiGlAfGJ7x7z8CMkaW21ZSkpZlsgZAUvpUjDQbFMwchy1L6oLi8d5YRPkVDaiI03EXD9Hn5whx
fra4Wap/HfcsTG8/offS6J5ECLGqpg4S99IgAhdV7/titcDCNgRZGit8f8LAdB9haL/jumO28PLi
Op0dJYmn/+yC3lX+h9gUNs3rbmgBdZ9ydtn7GoEtrbn2sCoAUKyyoZxXMxC/mKDQCF8xP8+/ZRH0
6WDvLr9hilTz+EuX6plAlVAuULPsYjXpmc0IN6H5NampUa94VFSK29c7XK3NFguNj127rrsf2s/C
8dbgwDKV1aHxKKuS1Rf4B53xEc3RHVvNR13BEkf6mwk4Z0lG646UMEVjps8eDyFuau3sf9ojftSK
4XhxmE9WZT6IeEjI5PnriUOoPU1VKMUfJOs4OfUNdIZ4phP6Fn2CsYwwoghalSFmzchcT8C89M6n
lGgYMxLZChvRDUrDhrq/dfOsrWaz4xQt4R/JwNUQDJRxjSTRmIOlbsMwvZm/Em8zuXF9hdHZrJtc
Rn4AcrfEbVmERvqwdakIYahuyy2YL9Av4d9EHJeEGRYy7EXt7ZAdAL8svfmepP0vayBvO6pBl2lF
bQBSvKu8YgiTf4WItKat3qBP5GklQzXI5vLS48X7kLCM9UfghZtZKGK43OBSCAT/3/87s2+gz469
DM306H1FDLEGxiZXB0V2AXOLSVOpGrT4E7w+1HTJHuMEEyTiYkHEN1P27rq91G2GO7aAV9CDUTzr
WOcSco549K9pVyy1Vq6PCHMhl3Q2HGkQrcodmlkKDd0xvrpUTyQ8a6znoDQ7c695weAcgL10CNt9
35ZgkyJsYGkeedaeMNu5mSu8iZrhb2auQZBlZl7vbZ46IiGl1CZUp0Dv2E1rHTLHi18Np/LXRzDh
YW6wBs4y0NG+Q3EZ2zk923w+K1sOeEK6+R+8B3wqDXiJ3aoPKYyC1DMKiFEVwKkdHwIe1cEzjWdC
tCqpkcDd9W7G0VhwyUeqcA3LhNG0fpfNCgATYHrs/MfewnPYfudc/2Tke2Q3q2e8Qsv+tQm6r0pX
HGnzTrlDt779rcyq8Aea1yXEiDcBVZfd3rU0BsChEz/wWNmfyScowVlgO0Ura2Oxfcapbrq21Rh6
DSE2rFsAZS/vwjBj0UI1/tXHDYLV/sLrDkoFBnCtoCjbes/9C2M5L9+SLXZi/GEot4TIc5c9ylCP
5Q2kv8xWATiNIpoGd07RcM/tDtGgC7R0hb47zGQsa1+WvtiQ7v1kYfwm8rzuJ5XmUK0VgphtX1/z
BDSU6Hh/89ipPbFapZ/Td7GfBL+NoAFj5rVUII/nNd2oSYhm0ymtvlUASeAgBytLAx6tQ7Py1b3J
8zWFjflMglYvOJ69cDI45anvjy1hp1svc9BNj9XXFGrpP9Pt4sKiGz4lX8nm8llcCpEXFfAm0bUj
h6fdSD5JhlCJiQScr15hBgzCVcSt0ZbeRAgfjaXLbijAeyZdZBxbaDaXEw1pQ803NrnOC8XhNphX
Y1dYIQDt67x4TMkXBOVDo4Jmn8i38ZSBJa8WKa+y0Y3AhPEcjs0n5wSCTZYbAKMjdGbrlXnGCYsY
1LY8HTSNRTCS3KkfgXKCbgxkqeBIfeUunRypZQ9JdegkpCVn1jNWM4g7vcku0T6sJrlzNq347DCs
VDeEW4bL515N8wnF+5K4ptyCwdfQrj2Op7wz6SmXZpg7s+7JU7T83iCfvGxqn/H0BjHNlWfqb2l/
Jov2gQ+18RkfiZGbEafXVsBX+SE5pEWQ7EH5Wo686jRO7yJ/e+yAPv9EYTgJdiv15t2KzMpksp3O
GB9zmT8gKZyK8AO8BcE7tceJJX1BTF6zJNYpS5zYZw55/zR73hipS96BRzP9g5XcDhIzDDVFxGl+
FKHtcDMDb6MrLdGWIX2jhOZvJbJbwINNGqVumMG41Ug3tGFcnJszC6IzdmGLDzgkGXmWpyhixBs0
Rz/z2O/2GBypuRuoEXOLg7QWV/lR5r9JC3IJU46L0qAA7l2O1J45itIGf3VI2mTyXapmofYBX8sS
IftsMxj4ew0ypHXVshKDeL3fwiNjvdoRWW5OmP4XvHkTTLheUgQEB0N0EY1kGFvD7lcTfnUMxe8B
FWBZtp75BV9TiTHryb6xrDyp/2uKZw8slDnyvTgeM1UxLKdi5xxcRXVWarzOndgtr5cOZ8TlTVV0
VcmYtpzUHBxpnmTn+X7lqvw6XMdUGAo0ysWI18ejmL4P+haWdkdC+Lnw38fJIxKt0LL+o1ZFSd3j
nyuEKnAEJT0C9AWr9ZwzVWhhl65hGbY3P+2EA5mjaiOQgMsxkA8tukxOSBEtHzGLnPQjZUot5jpS
C4yeD93JBy9STJguEZH9y7ZtWITGvLWkS9rigQ94lJQDgvAIX6XWceQARwk3QE80Hwc9WhWhZ24I
1mNz6VGWuQZHIHGdTclh0pYRBoq6cVOEB6hdpT8VbTVAJSoMCGecqgKlkX64aAqy+DuCzAd7dwMq
NUPfFI88DgOgxxbw+doT9eShzkPEyfYcW+R7QFPy5hT8rqpDJooDb7Q6X9HC7lGwa0Ur4zEdI2sQ
Gh2WMWOnADfXV0T7VWHfTOAMTQ5nVjGiDGGpZvLqY3wvrsa0GXOQWw6VHYVHes2kb8q/vJj3XyOQ
isjCHx/cWpKzpEdXfsP9s/NDuhicyW4HgTtzasSPDzAW5Sl53HkzgC0htxUrjM8ezj06DYc0N/ZQ
MCKMRK3sV1TO7KqdjzJ7hy9nMfCyOvllONR9KqtiOJEHzqAut8nEucXpFSBHofiHHpLQSxebN34P
MCAbtMwMuw2T0DkcRBwFGjpEJi0hhrrzaP9ZJp1asaFaJlqBEU63lLYHmp9dn+k/HK0XRbDtRX+n
PUKpR/yxXxBp4bdWbXnrVZvi4eTGDcocbfiwUkl46oFcemMTByYwNfc2TN2xZt5vUvolhpi8RVxg
JqvAPOZItC7RYuozHFQjUIU9AQeLY2WrlwZZgE2txdYnNeZg/DaO3f0M42v6+dcFuElN9cKY7V9T
aNOLU4Jlh8qXXRncJoNEW+E3ODNxiIplWKe+mpZZ+t4JNuFWeaofrkd+sN9jG1Ha6b5vC51ZTpOp
qcvXe2DUu+I2ZJ8LA6V5c7XY/9SoEnLmx+9F1aUuJCuWhGROYUkg3y6gv20JmtGsvECpZ01A/rGM
5BAvTPVSbLf9Jg+rLv5bss9TpLZkHoZ/1tIvjaBLdvng+htwXM3l+a2Ws6xjEGt0gtmenE1XWPJa
qyXAn4u1kQ26UsoehgAKp1F+Ia5F1vtl7GDJmEtn+qB2PbG6kW4QoBL3IFkv1EBBhG4d8n/DuIrH
BUZ+gfPyRMxc/3JCkECMDL418uJBFKbNmpBii+/990Qha4bwaKtiuDucQaj+Nf58/PyBDds9dwdj
YRePyXei/izXmZjcueQpg23u6QGVm7DpLJ4wZ0Eeqs+LNJX0lJIYy6biBNkIebMt+kfaeM1Y16et
obrZrLN59qoaBL2oKw+KicYV/AqFNnXsALDjM/DulEfCQkFJTGnU6W8cuLhvCDMZ/u7aoMyeVeW+
EzC6bhFO6WBifa1x1hwAvxQXbFtSCEzjFzHemSg3Su42gCyNRXfNEtkgwe3fb2uo+q3y/Ub3ljS2
Upf/DkpS/NwMC9LM4XmSaFyR5e5VfzgUYIG70xlHeyrnuP8l7wLcaRVExuvlevJI+XsGIk0U7PTM
En46wTvDL8NK6v2gzH2NkEy5P1tuEyxkRNrueEuRIhqVoralB3B+gnqus5/lt5dAdhYQrHz2K3qh
Huqvn6VpzZdN+7Tsq+VxRcPLEOrsFCD9GDx2mP+U/JhMiTU09MrelQIATt5RGmcjGWS8+98TJKPk
9Jn8YMiHGysbnTYxneHR2vZXOILKJZ/5qqIsX9Ans8qg1VD89Fq5+sTt6N4GQNrCIcJ8RlrPyUb8
4uQh7lMtY8Wp474VabB5waamLgCqtoSrjswIv1zzcK4bOOONCgzZ9n6GY6OmqpgEzpq162Im93Qv
xquwlr1HRXBR7E2FJZtC5aOhqB40CsVauqLk5rZwOMy3DpSoPT9LFNOvY8FQ9ZtAFGHdJaXGhGFX
6m7Sb9avx1L69pMIxGKtGcHRdzvG4PqOoliyZjqnZQoXGxvzTfw3gV9UIMy40fjlehZ4M3ud0vp+
XVCHIfjH2ctfrxVR+OkZRKYj3RiMThpwM7tJCSaSUcvNssftq0OpTYItV6wjHpGRwyKikahYmTSu
UwIXPi1grdGZrWTgvXASI0dSLD3Ek8gSwdTa317Exbwa035tglyI+Asl/v6B2T9PU5vEGwC9WXW9
CmpCLunScWq6wR5zaw/tiPRGrNLXBAMmvrc47jRMfx+TOqSa9iywv8xcA6DnlBkBoAQIESgUiJsQ
K3gfwB+qMM8JOzsXX2oJx3soR17nV3SLPvP0jCK25+l+nZdnIWYWxHsuCxbQ0tT2ny7JmYtGknqW
ntYhpwuj0/EUfPzxQkpW+HmAzv7/q30bFglLmWjq687XcAEgcSfLJmLQ1xHj+btIKSws+4u74E05
h0hujBDVz1O3Ol0xudGYzvN76T2Ko6d40h+m16BHo19SkfmEV+rGjwpYuzuCxt3b1Eq/vqo2uujy
D9X96IJtrTFThIPFVkzg88w7A4MBrwWhEyc69jhg2V8yh7q79ttvZQWfCHvqDPL3k5Qo8FLQAu7q
/ogsZRJWs1QTrlMaAKSNf7GESYnohzqwR3UboN4f76o47foyTo8ln7X5Sbkdm3DJpqLdy90OcAvA
ZLYn+DlKK2imFNscwG22ijo9e2P1PAnmKlrYh7zlfBwaLJK0bfqIcYroErGvqb0aAKM1THDCsaJi
quFj0mnaRoatxWE7X/jHnqtjapZVFIO0IFVMjY/vdRkBP8gaMyuUQhpY2BMemNExsllJCtMz7pki
/UTjV4jWGs8bFgxrzdk6P52INHqBv324fX5t2GQWwacUWAuC8kCqI9A1me80TBuG9qVkIQUHFkqp
0GdERGKRic+OTbjO/Dx9Qx8f8HpS9yKiQRSgbv8+QzsWqtK1fwWSsAGG1735uAy9PjE0XmRYubRn
1/CMyDE+Go9nwR69EHOWF6wSiGU++o9NgE9k4KjHOLzeOpxmVBQCMT7dK7fGBBfulk84TJIe6Xow
czdSj1U2krfse3T7eYFSk549wnmwcmF/rXT1Wnri5hM4q7h9Z6ydaqbehE7VaxdTHLmvkqD4prqo
ZiV7wkVSmlk9zp5BfrckjtElrwFpWb8vbSoc079kcVutJ4hREi65CEzK3CxHDBxrAitO5qZNAaSU
LH89KQbTEQ0rVBQZiTMXxTtY1/wC140xerxJEQknqtcaswYWgXXV83g6WBdn+zoyyf4Xnh4rwTnY
KOfntVCPKevaOogrTT12uRVWdiRoygx8/k3DOCs+MZxHjT4bvMPcfovkr1tLJty0KQjg/CAsxpxQ
RGoQSej6JZBy2jKXZ0WHv9VbDp7Av3B8+enD1o6QoFdT6RPfW/W0alCCXy9tMH0wZe5xVKxmRYSs
i+B+lMVmm3ciA77jSsFww8OU9VZC5Vd8PCq4BMLHsW/aYn/npwpVyVrIn+LVI6tzDty9F8+WQ6Uc
xD4PZWIiFWBhuNQ7Z/njPJ9Vi8sbYXt+zggEV5eBN8pHn4/nmfwDlnlRwG2iBwxWTrKlbp88Vy4S
UpS26ZigOvVRNh27jeEv0tFBd36Jn0uFc4MnvJzPLgN/4ik2B/AiIRWKsLduOEp/D0Cup+AEjYpK
7V1vyLgv9gLeA9BSlZYuAxYdL5zG3JdbJZmqcG6fdCQJBk0+04UZfdlrh1r3aTlL/9yAFlOeVTSh
CakrosVdLJxRvDGrHY8yxbBToHM3A9KJAGpxKW3606KInxmw7qOhI1fquEcyOzVQP3mAiRdyox/8
JmlhTv5JaBEznsrN4vag4+ucv99K916clVmD5mfI0+/qPlZrB7XiyRQEnO0s9Ar2yJui/cnW6xWr
jfGRK4qWN0gRIpZb/edqodI8112JFDheTX6zEIecpvtLt0Y2kW/o269WkXheUGDS94ectten3BxW
gJ6Ui+QX9wHpthXcC11nKWIo6ulPtfpWSOvHNMDpNll0rrTCRu3xXsgdKchtju88GeQWzGw0VZfe
75jrHtKCUcJuLCo01s48G65urfaHw0w3AVa/j4CFUQlya2cgTPtaRC49lmTPi8Rxf2wpnbnzWwvL
KFXaqY1FjlXlEt8vwBaRvvGmX6HLY3oInSG7kcyk1G2ZcXGJuOou9C6dcPqebCUi+zpli9+aPzcR
k6J//v4PUGI5C2iCl+/xdwq/1si/ZGgXGM3azIlpEr8uhLXFYmEWeK92h2GSvIJN09MS4viQQA57
j0FwjWxRVWNUKW8PYQDBAZuLsqWKik5GXtyIcEwegSXRlMyNCOcaNRxjvjPf1qV5oJh/c+/xjNZP
+bH23iU+Xr0rQQIGkTrkRu7EGQA3IcIf4Fj1qtTPPFekeD+4K511K6paThhoMJm+g2a7qBW2PUhS
ggh3xUsVXPjoxfoRldM7ZiNrY0hQPvL3jB2yx+N0fHITdJNqJqwWaNTIWaJXX4VYX7oPtApmiz9d
mb8VwZuQ6EeCpA6E7zsTpj6O7sPtuuSL7wGApNvbJvinZv71cjgBKI8mU24Q+oeBCIkDYFXiDL5F
Jbm8xLRPnOp/Ujst4HfqdrVBF6KOs6H9uIUKSdI7miLFxMqvgDTjiYOuxW4seh74PVIDEzQh4HPP
uOrtohifgZVzyfunjz6m0LYpTh6AI8iQfYfA3XShvTgOpkYaYKQPtYk35Y8nmcYpSbpAHJ6PuiaT
pDR/xtwB/xzSRfH3T7WmU9NFyn+omCoXqvcSyH1IjFMyuRzvX56OlUbIsThwZXlA4P8WJ4h8wkma
+dkPbvPoTPIi5GtiRRo/aoHwp7+graW3TG15BcExw+u381+5JyYvJtmRtYHHM3xLfziLvC5katkG
8JcL/ipkj+kvwMq2nNGT6655BmE6fOr6SEW/KxvNZ3Qyq7zoz3Zt47BE0QqkHxpCZ180rt0d6m0k
rualwp6OLrRlFYPuA1Yyfkrr8TOMdwUz0u2vQkYiJX0SDnAk78opkblWu6Ta8pR0dot977CCxz+0
trH74FV4HvrKqcFIvUm1Al4bSdZOUCM/wZomUkbT6TYVV1BSIHsQXnebCAjGxSGd+mZKi6AODD1p
S4VM+/e7UwVki2lPaFj6/QEkoeqegrkiAUGidBELgyZfuUjC9dGXWZmLN7MkjnqfM0NUTh760Eb5
Vz9urBJ4Nr9Ih4rs+8SqFZ5LH+IculEO1bG/JPHSF0n1padL8NmYR9VMgcOolvPzl3hUnerGt7ra
vanKPtZLoF0myn/XyYAa8KwWx8JCQm7kPHrlHrJHRdUEsAPqwmsWkhoE1QenX280dJnMpgjkWKOD
nZh6di5HiM+9xg3BthLXguLphd1PXq0LaV44rQg8ACNR5VHTWnXfflygQkgOIzGcV9xJpV6E1t15
6qv/S08/EWWk729UVXza1BVVibRHcsgi6KpkMvp0XIgb9MoYtDGcpjBLpDpBCaQ77BwUYJ/p1+Sq
w/WZKSmLkt7cqn+mG3DHOXe2bmNQHXY7xegNuuxMEU6isHDBQPExfgF+cTaQVZoWoqKnuxbl3tqb
T31WKE5lb2el3SFygvJ5aI8Dgs1P6HlvpyuH/3FPK5RFQQ46WjB7JYcx2FvYIThgq10wIAofWQv1
LW0eB3NfsneSSVEL2v8imMOLDPK3M5i7k5yT96A5u8t6Dat8W6m8Ju7124EuzGLwl+fXPcZAY6tv
7eku4acd38leieq91zWweDwFfJlcWufg7DoyZPA6vaU42+hB7OBJ9MJ6+s/Cmi4mGg8qQDEc6gX2
nI6Z/8oftZxFCPfo2i+uySS5TQ/EwHSMAYV5jolgWHYIr4vnCwT6G7wQGZtRY3yz0KoVMoo0fHnZ
K+2YeJPlHzIdL/c5kD5/reoei7ZwYjC6y5Mqtk6ERMl/SqvnFEYG0ZA2AR0cwEmysvX5U8OnS4kb
JaQWlH17ySIjyEgKIKTW1elOn1/5lZApmNPYqGkY9D4Mr4rcn5v3DuZ6CcdbviT9F70nvmy0ZII9
HoSPiFfH5c2L4wW7+VZ0rQAp4vDFBdc+rTTxYp5bxdeTy3bU8P9dHx5H6lx7bv5F69DO3wvMDfLt
ANdt1jG8qtb7ZQfqjdM0Y3ZZjycYnKxj3B4+S9T68kMOnS/9IxpIgTZdaBURbKZY3GE5Su6xxUG/
bbunjvS47O7EhLd5U4+0fUoDqh4zLbeK3YD6gRldpgnmhk6M3TMDqM97hSn8Il6ENmSBhPjAYhBF
vNLRLWmzrdgvWiN9PFFKbASK3WYPyWHLejofJaslAEzZ+/FRTUpXKtQtHMxsYYMDFvra1VyTiNR4
PkwKPVfxglDsiSfKgybMCuOObfmozB5hNCqaFEe14koI6khStONRIkxZxZQyp2YPCqWrjn28XNBs
fprXgHhinC7fsKqDO+QAyowcfWH75Rb5cHDdYjWdmr3YXDzA2iIPIfjg8Ct53aDg9vZq3869um3/
Ldb3BvvO4cLMDbFgzafhykDRA2lE/BYSzn3ttkwBB0cEW8UuvaxaUs6EypaioGUBJHrNjxNiMp2G
vguyQ5l4F59TS2guuDMpdp/EfgbQ1DNDpweGTucrFlFVZ6IXqmcF6HoYQKNU4QMXhgNOmL8oMay6
Cv5Km6KiWWsdheMDke5QAH6JYBAPZrMuTXh6ISnMvjyOzz4WvBViDdbdvXT1GUMLcCdef0sx9yE/
lu496vMIHvT7Bu4RM+Fhi0+9Rgtu2HguBZKJp4oBcD+QoRP/kHJr5B1Uzah4oRMceVDZ1SoyEtTV
3SF5BYMjonSyqIW8mALtBO4c3BdcraTZL6cCBg9MbVUiSOQP+BOaM/5CnE9QHfmQxXmWSJVGTVY6
YUElSp7kEOUqIcmYzzZarpszhebf6JovKhu8vqz0dzsUDrkPa7LiUZHJF6HtxS6+ikDqTNd0IRxf
k4zGUUIUJ4ua91GAHC/Aa5P4uF20i/4N8XTKbK6yRwZB135c5rDh6varE0Vn+3MzQsr91Qm+do8y
4b+5Wwd7QTcDiNggIqeUyYaOxG8TMju1a37rKg0axPgP92vZMJ9j7RlJ3yqv0MxLXOnKb2m5/L2q
hOEFlijqF56rfD8hSQoDFGVcKe8noZBATRES7pW70awz3O8YnpfhMN/urna4mjRIDno1MCruMEg7
l6AbkWgrmdTVtADU2DU4HZsYs9SgfYYMwnedT6H7+gqN6RrAm4ZRtSbXmPg0fb2nRIkVl3Rgzv1Y
+X/qTFXRwVeUlMH/SyYFLiQwagmFFM8n0Mphbc6fykdblHRTiG9s/e6+mQWmcs6tHDFtK9+jRKsy
Hl+laiA26bJ3oONSaFTyXD05a88tdF6rPm/dDTeIptMyO0vgIjjTxj18HCfG4CyE18UUFfL39GV4
gxVwb99atLWHsKocv99FEvNHo9r44a/rMMD6C6lCoKWjgBUq9Xoq2BRmm0CnIjBixCNgFA0shGnN
k/rRXaoCG0JAjhdcd3sILBZVu2Ulkxn1cRN/OUR9NlNecZPWNP61G24m86w4xXo9FHcH+r45Nqlw
KQ1/+SRrkf5l/RIYYrBki+CDGJpgXuj2W+vXXgbngmUJ4mdE4vCCinJnjtNkwILmk6YdaGb6wmW+
sUofTHdyTo4qJx8z74DFOiOUh4wF1E6FbJHumOIKQ7ULtveP7g7rRs4FkQMTvb9D9V7f6IC6pSTb
ka9B7j/oKvte5TEPk3EZ9Hp1Jq7yBkyWcF13nLqJr37X2FnuBYYpq6aiDThNPpDDCGN+Y83XvPR9
08Rci+LxE8/ZQTKK4Da9Vlq3vpxFxeAqTKrhm0Ri25cH5pkjEp7o4dVSR8cNttM26YLiZpVKpAOw
nvi+esxf1dhuCBqNYn9rvquDcORBrFFpgoxqLdjdDH5A0YXI2jxBR8tTE7DHQ2dWu14UFnxcnmgA
PN22tTXW1qqXCgDNsPRPLk1Y8ZoZZTJGMYHzOrjPJtTUxpPaMRvcPqBLBOH9GcF0dS5FJN1jzBtb
vBmH895GHdcQUElgzqdnt/JfEO6SqjccsYK0whlUUZirPBp3JVex1ooA1GKCG2uuU2xLCIPdZzJn
B/FnsIllwGXTa71XQPhx6SoQ7yHsptpkWsH+9XIC6oqo4d8fVe1fGHRhi9UaaJ0u7XhvxI6n3Y8n
U2LjwP8qpItMWFJjOvu2DvnosvlHV549zg5ZPw1ITWXma47XmvFM1Acb3UG1hXjTD8fO0LrdWF/a
fARTeRDcXb6Z66I72PU1+5Os/f0fApl59S/YiFLgsmtCgiNEeEZVislMGKm//+XfV9Sox5++HbRS
rh1lqRBe7jIVFgjy4gSeD0L/wmdlBiDORf0gWzmZKzzozBemCjJcjyyIDMreidP3WC+VC5RFDvAq
WkMfkk3Gxs/OFeZLfne+cVeg3qkXtfT6wKbMjEK2x+nrwzAmK4FWMiuBOM8DNsoKiLICtfWzLb0Y
n65ODuhCU9R+1IyJJgZ+Gily2c9Hd9SsMljK3yqUITPzAgs/GGDO4V3VICG6GVFu/wRhLOZJKHhJ
mg5LzRaAJ0N1mRVSdBrZ+u67P5eOVpd8yJ7Q058oeioEUzUR2cG82g8qGUt8Q8RlI5b98bYIsXzB
weSkhe0wQQKbNiHn3ke/Ou9yCk2nGFOaXSouLrvva8qzfHTxdkTNouEbNDdbKWOutA0PijPj7ccx
Gybi3s5NwUZYHB888CljdWSlga2/ti9btMWe/e74R2Un/Q8c6vSSufJjYfVnVpoHgVYNOCzKoBRZ
Nf30zyG7UHtpPXTE8qOo9H2/y1n9ZxQJuENWejgJdkiAtaC1qS4dYfeHKOKaHarJWxKuRhQYn+HC
cF+OTqNzf/ZWAehf8gdcAVXD35m7RAVDjWdfPvZJO8Y6sE+PhcpiP95nCpIoQdbPeCShwMjhMLRx
gcZHDMdc9654e1K07Mb+HEYk67Hcsqk8gV/zxbKhPBvCdOduZVDlndQ+pn1nVWq6R3cZ8NMTjprh
Qcx8ZlVPQP3Q3q8hG2xQ125WwBzgC0WVz/IEIb+TGlHYo+K3vjHmLmRGVXWe7rxUqo9AU3iu+CLM
e/+40JYFM9ZoxzCL690iQXGCVhuI1sDwLiAd1w1e0GGLrqOx6TjiPERm4ZM2HLJQ50fxl1wBHJjz
ermmr7kJFZICjGSqKA5mOThg0seHXR6n1jGOuUcanVW93KGxAtL9eur0OD0nSwvSl+CSfUIbXHvH
NEFxNwWkCrvuezF/7cVdys5doGt0H2MJw7giPTm8wyvsZg9j1DgMdqe7adBuvgP5g8ailTIgoMVB
DBbFBf5HubGhpskFM4nRSdhmJ/JYzPbS6b3YfzQLprVqad9pS6LEHqnnJdS1eOc7C5E/cF0oEQDf
Vo6R8r7bKtn8QBbVuUZPWnZZO7UZxIYP0wnrqt7IcaKhxe8Uy0usxozlULCPYy1SLW8YVFI2tIxG
9e7D0DS+3/fvHCvQXcYIcg9PijVHfiNTW+/gf60bLSCyLfFmVWECopDMPVu0C5LFPMCS3kDJfQaj
sredwHap+5Ht0ZdMQpc4RO53IxIj7FARjAFTZOMgcg0p7rGnhcJ9MUfto1lANo2qjZcYCsZ12pFd
PJBCy3TK5oPSqSXOc8vi0Ec6orx8CNSVNv2jJ1G6cEkNx5eJCvx09pzGm8z14+C1CONjuh5WhBff
Rjd5bLnWPKX8rj8kryJeOGRJgzja/84YCyugE/JKKWYn/UTWjgDMIhBMrIlPwofVVsBhKa/EetYq
VFZledjPyoEZuyl3kjBhsV+5a2CphHb3QzWGRpur1AGfJEeYAzdYGL6b7aiH+0blNj2TFKSqg9h2
dQjPmgV7vPZXj/ntJ2GAzIPheu5YBYTzdGOurtKXNL6GKCZZn2LRC3Bikbp7ft5wBCZ76Lj0WvGp
C9hJKdUonX0je0psaIxAlg/df4xi8gEDw9U6JJiciCKVnm9wl+9LSpmyrZPK+EA06XY1seI3WPGg
TFYwD2Eqehd0YHxIbpjyBbQEMz9nHuRCs4RnLOEnLOkJGfYYv3CoYdn5ezcwZhzWs7TWMOrjuRI2
HI33n9y+ZWWTUrKzEV7RsFbN5N0+oCNivMCgphbbGY5oE8S89HQMfgUPEMqduhXFlC5jHiFF4vRs
MVOi3p90c4pTqd+eMLGOILT2C2F+5a7aV2zuc0UVt/DRz5ZhH1iF4ykjzPdWAHxkoZ+xasBFoIBm
X+k7/91yn7deRjgGjmw00azzLc2Wr4bjnkkPXCd+g+ySSk9CuC2YSjl/QLfYO6WSCiAYjlKMdBKz
OJ9Gd5F0yHxFFIKu3d8CRpFd4Un7knY3bJXnms45fHWvxzM8wkmKet6SBvi/M+UJH75vzvv2o2pk
Y9kstW9VfTvEpMiMXpYK2yOQFph0FQPsycIJIGraRa8njYTQCdmjbE618ykTCm4016d1ylrKA8gE
lpXEkoYG8FWKjl7BGVn6GfZ/5dmisSfyaiRuP++ZutQ5j8pTSBv+czl2081l07quonaJZeQfqS8s
onetmmgaaNe9MwchrMXd0wOAmMbY6AdRkFuWzc8Ti+/XzmBGCvOokEjWHje4f/M2oyRWqF0cgqvQ
KfjWNjEuz/dZVIi3VIMA8O2oFAIxrhR/D7NeLAPWmgAIbTwnQ8xa9WyzpDQOGVpSAaasJ6bgg4ch
EIyYk1CfEnReiB66Axtl1jWytTT+2ePL0YdiKmOqrqxxkAKzrRCzw82W+24wkJmxRTkNE79Heo9n
lJZ+azYy8tlAXqZq7pFpSokWuy+saIPW5OSX6BneQt9AUlZjPis6A4kGYxnaGvudpb4mrTgWdMEJ
BkLn9ZOfrysWQWJsuafeYSf9tcNOVApgJ5RCki54QJX2TEkX5RKtmHBf5ffAvxImplxemirJWkiv
g+Tep9RNbPucu9EY6J3PcfMWMkirdtiESpwj66WR8JRGi12Xk63LlfREwSNW5nQ0MvZGFzeQUqEb
lCO9OUGBjDKc06fFWGjPGedC3WUkIYl7MQfgPi7rjbmQtfzqsTZ+XuZVcBuhOGF0exxY4tknOXw3
I2qzVxIPNnq3+o1uFZehXowmLGZUKr83gWGX3meYJ+pD/A4EWTGjh27ohymln6oezfyPzAAweELj
19eCjOeqL6kaLD8sm+GwvwhBp9w8dnQ3iC1FGQ/DeRgZ96OajCEoz8iSuY86t16/obHrYxuXwuw0
Z0y0zB7gJ4Oek8mlzoh23atkJbZJUmBPl6ktzYtAIlQPFalvQMkXPjZ9gs90hAf8hD2Kzc4gjQLv
lZ2A7dIz/5pM9pivokUGU3wf4EVo2tZGUH6Qf+YZ6bSuAzIvDddYOXB7lYRpAvt0A3ZeyM1Fl0To
qxoRKMp+SdZPHgSGy2qjOTRzPODJ3BQyvEiy44ZdbSyMg8sBArRcrcEMRmgoAgtuyyVgbIwlkGfj
oeMoZ+rqj5Lj3HU4U7m/7InKZ4gzk5cbwPLzQlwDe1obMyp//BmIx8SpQkP5YpCxP6vA96NDj0Bh
/+jspQP6KXN8Ft8EagYeGZIyiiiKh2n8ZDiMIY7uAqyNfiuUV40g89adKdj3+PmTJaKGWKcSmoFI
cIItoLbNVGfgZrTEFKYmkjlC2veyNctcoSAddsShIc4Jjs/BQFhLO0T9ptqqyDJw9gmkHKM9Sirp
pxFEEO/1G+fO/75EbkjFjpsrCV6Wf5IQSrs+BzKxPnjphCpZvvnXKLuJE0Ng5RAncglxWNNphStq
BMQNbgqJSoSYsgJzhZtjOl4x/SrjMZNtnYU6eJeQKzykD6QC25yOdvP7iVcKBGJyXyZtrxgRS6Pk
EIDIGoD03biZ0oS2kuK7Oqr6rHujoiuLv/ulBChJot8ZkG0uWDEp50aK2OJpQCxaIn4Pud+XnIk/
zSWFv97PKq/nMUgNkZ2oe1QvxacmqB3NNWwvfRI8B+sQEic+o+PL2cfSDv7pCiAhnfeSym263IYp
HM9IBlzISCC+5MaiUPm7zngm+R5UNmxgREoueDkJ6fxgo+C1NnLNPH3vbBUhyDr4lt5wxWk710FC
LJnHV94nSR+UUA8M33Q0U3v+kPZCtfexQzV9gufx2iWbP8NeXMgJ8OAkS9E8fGzHtLWFG2Vp6DJv
2NTr/1LYWzCy5LFfdF0lOLCGA/nXXqV6QMgCJJZZmLd0/5ZbDnYIsjkR8s+qVrAunKojGxGJb+6P
3nSjxyM7HIxuXI2Gt21JEi/GhxxA87gdA7OqCtECXNUWrJxuKTSdCaAhr2ZBE9BdVQfZpNrQCBqn
2k3ZiI//Zq8M128OwE6I3Lfjfw8SJTGMoK8i5Rx40pD9JPYnxottW1xkSy9vRazrtCZfxwFdHLpX
y64dTgTWnUiKWh/uHjwJ/y71auwr6XEtqwiVRd8f5mAZnjGkt5pzIOVqjfs0c7o2oBe1JgbnGuws
E2m8GMzeSOBOCUD+4z+zkbNrlNmQZyvYAXXi37YipXZ5Lh5xgxnRRv/5Lb/hBEgREHmgzGojWQvH
L3IAEUScFIOjhOoy9dlA9m8H4gxx8Sk3xi+ANYWgAfxScBHIspxY42vvUsbCdDTVc+82lnrvtwob
5AB8tkozFrQ4vwv2EDGakSEPfxL6PpoCPfKxwn+h3JfhWcgzBacb4UENkMhHzH3SqcYf71HjDrre
/jc/Gcep3+TJUqtKtV76yuvyqwYZUGr2X0uYrMTbsODk0n2+wfJ6xugIHjsTXqvlkJK52DTIjSfJ
OwSlPIWMyLQcu+ouxd9eNjD0iEkCuIxL1MeURzWFNorzqY2bQspz0c8gVkaDNyY+KV66ihgGobTr
fe5c9JvaXxKaIjw60qzeUPh38ZgFe/+0JxY+OB6fsYAIKf5f5axUKV1CP/o35E2xYhX4nPUQlHN9
QrLwaSl2DbnRTQs7FHy5LD9lxq3B5xofFBx3mGciTCObJ7JAB5UXWZn/40fZD7MkwQWRiPnv4SEd
9uDXmJyK7u/A/QGq5/Qj1GszdzJ8CMkFL0xOJt6FwPyd39hgUsJRSG4nOdIHFlvr2Ev1uhY78bVq
7wAJxyGBdOrsizxlzyXkk5CUq5pQS8FoeBVX17EuMERHot2X5Sr9y+HptmUAKoM0OGvuHLqG5Jqp
/WTsCNbzMLTHyF8RxNI0oNIMkQ8KkND+444aSnDRzkukwNWWbjsp+p3vwCn/vLXS6SbjUQx3WeNy
WcBmkAsKX6fS+OHLkuMyUkL5swCrkQMarv1s2ANhVFHnEKSRIQiEaj8ZDNVszE2cO5clpGyeM0qn
eaOZXE02NZvNPIYLOIX6YUhKORzpHNvrJAjli0b4lTs2brNzbJAe6ViXvfE7i4lRA9Fi84HV2HBx
+DWEyvpRaUPAb4Hlzj82bgLwiEhqC/9SoqCoU4q6zeQQzxRVdX7lqRucLrRkWa8Zh/AuHOTy7vjN
sKA9E3AmX+1grlXZfV/+HX+LAcu5/QEHjOcrAEdq4n6Ap8UhvhbC6Zo7vg902YlvOIQm9tvLTy5P
AsndITy+Muzr1sqmk7Qww8GXN8/LKgzFZbja19V/nIU+g/qaI/X+ojF7B5SGB/DU3Xh43XCcO7LP
sKB+61OSw97fCR0yNoa4Pi4INGHlXjwoIvjbidhFuLhY/p8Pj6iZEKStl0/AtiHX3VoahwQNkEx+
8TtX3lpMr7nwOQ2E+DBQepDouYkJU/04+FAiRfKAi9YEANvoxQwNTg0jEELxWW8/Qvsnz299F3Mh
9PlRBjBX8cItsvAVoC73EyvBnNT5tRy53ydQE6ZE4DCKe3Q2WtRzdc49lbQTUy0pjhHAt81a18bv
rYk33y0RUrG2HWMAB6MPFXM5kQuy3Q+xEeVscTei4i2zgkqAqO4iRJlsXwvMPNGsS87scd8yWx24
2B/ZHd5YTcPgjkwnl6t8BZ25IVPTXubpaIDiHHZvYG6flZaRIN3D5Xgpna/5k1L25yMr1Z2JnKzz
jvyE9Rjp20Vk/10F+g5oY96pMPM0/xZ6TrRd87G2DGcdwVhvYg4RKMEm4ysv2ch3NX7XRt6f6aWt
4XZIiYDrCSlbsJHQH6yoYgrU4XngWS2AwJv1Bsz0VdiNx1sa1ngqh3CU5lZyObOwriCeAEHM7dXS
TAlPxJJTpYN/TMdBlSL6aikSyzhV3KlwhmnpUfO7bilud5rohk/uLvJCMkGHjC8+hAC+QWhOgPq9
m7gmtwPn06OZu1rw4SmVEPtDuMPWBPJehiS3Fq47hMkEcFssKTq8Fbnt5u7DSm5eFTQ1MYxeScA4
LyqBtygJncqInqPMwU6i0e62ygOutKxbaIsfvFgXnY99e1WCBYgHuxS7LqRbYVa7wZVtgzA6iwWd
OmEbbTQd4uhBCMU0qJ2h/ll92aVD8dZgPxT0ZPD+zSzThWLU6UJCH+OQrnaMchWcTI+FXYvL+2oE
s+ri+vqVLX4+r5kdtClOZRcI/LU7NWz0+rFCz5kXD87rax9Io0CIBZ1a7jyiZc3gvYWzWUxtk73a
vKQ7WAN+B0DWWbOEmHNbCGlHzea9Akd0B/eCbcq6UMWX07fCFdC8PH24QmxsY+y38nCCiKphyJ0u
eZelxBnzngqHyOs5vmY2+k4YpMYwv3+LWyjjnUWmGdPRD+BWzaHV2pnLuYYyrSF3gRxs15DtUcrf
xaRJHxZhM5csslKV+v3UB9Kp+4741ECnA6206eAjnxBdHcfNgPbZsWkHRwiLzu4tzQkiQd4b4aEn
lyqBDR1DyDdlnEYo1sOW2mdmoGQ06CGGSPtpLxmPYDJNkbVUaTPsT98yMsSaq1dCISA0IYNe3Caj
T3tzvHXWbgkCBM4w1JrII/nTTb2679mn0sV81wyAhNPS8lSurZAkHTvz879P481/9K6v0yyFi/Wn
MRFCidjf2m7sD4J+plx3XQje6DqgNGp1o3RMvKHfGufENVjoxhpOxi0+5w5dFLRjCl9RD0YhHCHd
tE5zb9N+9VvcFhpPEw6UyVw5VdgHeLsS3rMWIVGtGueqPQV38y3q1zaqE8OLV8uoqd5t/ienVJyS
b6smcjD5JynQhLLNo2aqDqqPFkiGrokMhTNiv+NJuaJXBdYQr49D/k6a8p3oh9BHoseJnboL6+Gn
PL9bmeJSz9GlyLC2ADn6baN92HAZpDxQbVDULBrO/n2X/dgss5iYKLVybeSPcFrd/39BdE5GToX/
Nda2cBYMhtGTdbXDbb2F87kQgmQQKw1oYTQv4ly0t6cjL0ek/AuXeAxs4vlKmVPt9zf6jVagtELa
MglBoHwEtU51XqUtXSlDagLgVdvH1GbHBel66MPufPIm3MD7uq6rIewTXwo7aKC1sNOZpNxMyXa+
cVRw7Kot8tBGtVb7M5lCXIORz9jAgyfyHcEAVoZsp0BoWXg9p944O2M+eo2YukpJXFDMJvbJv8fX
axWRXmCHL2L/JLUVo3f6fA9fh/o+ZcYGsKVjD+IDQKGH/m9lnoWCyuhMpEyqp9itCU0hhlFsBGZO
q3Pyg+93xzBNen5gE+jMhIhIjsKZLq3zLPVply1qhZNmbRIhU5pFLrvPvmGbDUs44r6q5AAQC4iV
ikHG40IZH4gC0/Oo6nFlT0/6Hpfgge9X7OcNCyo4rNLJtoJyqC2rZEaJGIcwZptNAKpSjOsT2mN6
g1h79fCXt9ErGny3e+AaioFURimo0HaWpI6bDdez0db2iBlN+Q/L0ef3KAKOWxo7undM8ZAu42sR
eX/RH9vWB5oKx8sgOa4vmcfKHVD/ABSZjwRSQTpq9/1pFx4vpiahFepmn20fc0BhlD9jTSsTcZ4p
X3tC160fDzGMYske+NA7WwtSFw2wBYJyiZLbN7bRL8x3Ib4fUGdjP7lqnhUjuuHLnybxt8Xg3+LV
SdKv5Jw385V/lYegS19xYOl9Trlbci+Y0dUDWj4s6axbMwz8Pf+zpHvoLjg5Ue+vg/K9eCh3m1XU
C03/m42SAlryFW2n07Fdm/Zy6UrUn7lbInTfMPhcOaMJ3DEdy0eW4mQ4VLcL49Gxzn3fqFVtaMkz
5uXF0vMFOSp4W/REOvA69Wx/ZT2CvVvSWKgx1hCt0X4TL/cLMKjiVf5PW2RoC59dh9cjyAZQMpCh
ND+WcpE69JO1rd4AQwLM6eC0nyvIvEZqek1bp3nGMOH7sAgxcKQTnxxvOWPy9+VPxnkoeGbkHie2
mnArDg0Y6TGg9sYlEtGC4gSgJWqg8z2Xjdh4LOXrC4MKrMCOmGQbOQplYCNoDfaz4TtZVEKzwqju
kzyk9eDtr1An/Vr61ZK8XjdZqYMGOg0V4dQ+3s1GNhk+UZeERwJEQlwM/zzPuKRZlMlIGhjMzXZb
82+zfklKg7MEACLh6oy3wOhTfA7EcofQDWO7PL/MtrVRzwqlPJKviqg6eFEIQkyhOPkl7X1kumLJ
fCelGtkQpxUZ191apf8u4bLzP3zXQMsTallNoB1Q3H7G+IcWKkIzVjFxBKxOCtKFtxXK/hq7iGA8
Bmauu88hSC1gk3zXyj/s8DrDHJ6VmlYs6w7WtAyhPaM2vOymA428qnmPSbs60VxPFSXkx40My3Kw
aXqkFLRp1DNLjaU8FP+woweOz3NvSc8QKth6VXI8C72/sba68vd3ze/INvvysFLV/bgqPurLoea5
tu8tnXtyG7ifJd2YODYb/JP3Q3mF6zHPP+gU4rxUSwis0U6GS621K4JCGKLC1RiKXqM+XiOj1W/t
61h9wMUq5rLFbmYlhIqfOBYICCgeF8I2i79JM/OgV37F4SgvK3mckIDXEauTKCNJmFJyKYRXkwXq
BIBRPz5A9B9AXyK1FRYJCq1Jt6xZKWzjIfRZhBV/kX6bs9WfnFSHMJxGoy1EZj+GUdaoig0/z8Nv
wvecyjift60lD2JmchIJdLgw+siZrwlWpvAXjvvh9+z6DT/6brOcthX2SVQxyExvpiBsbwiSWOZl
+/NZyiR0vTsfMCRlLakXuSdY5rtpxHKfQ+QHA8Yg1hmxJ55kRTnixfE6l7jZnW+v0InwROLmIugW
voK6c2elPjsbomp64wT+5VscVJoltdj0gpgjS1dM+c/S9+rrof6eG9Ngq8vbuU90CdXzMmxWs17C
+UccIb+55bbU43CBchoc/+6ZNVibrem/Kjv+Gkn9jLF7hMiWEgjacCWiGHUJ3SblIuSHX9/JMO2X
hWnSPPm9LyskERNwhH7O2W0R5/Abni/dF1qT3s2x+RkL8xO5+oBgXwQWY4fvrpxTZ3v0D1gh+9tw
HyY5P5G7pjzROOLqbICQZ/TWFcSAy0FUpFz9odxvCvQ427i+4WAgqckjaVms6HyItiVJWYqjQI4D
CdgEOxQLis16FV0redyltRpKsppJvvN9ufzKEQtovF2cyMqYPi8ZlFYVHzwzKSvVEiS3+DT6kHiL
cJvyf9fZvNR3dNuxb6DHaLqpIU0fZf+pGRy4jZvhStVCi5gTsj84zUj6Q3Vmm97fQlGhFT0xgZU5
EEcM+O49ELh/lBsv4tmk3LmlVQliwQGyP+S6Hy5CdNg3g9/Vwna6tLDZkH2oo4Co13Q9vULP4LuQ
cNqn+jlIOg4mhTXcy57049h2fX6htjX41kbrFzPL3r0CaENoHS2OkZMC8a8gyj7CCuZfSgAca51v
6LJu10jdWcYCVEI0RKshIF+boKtP6FpOtI0smG5D3fuHXqqbJ3j8pzk8vL7Jm1yHMwqv8haWO0bw
mg/etJjO68D/PXiJR9GBL9EortGwyzB2VsODxK6nsENdlwRtt4heZrL432pNrp6jT988S5Bg9Ebs
HpFDtVO7rYQDFGF4VzYqdLD+HWXwbW++rhV/j1+W5Qe/DeIknC4BvZYFYHmf3pS9r0w+UqAk5aF0
nuurO9CNMNvZQcq3Jtn3a2qTUmPmyhKHYVX/GeRdwE41+VmsAmmDZPVTsPIhTYm8fU9gypYB2ImO
twfrPWlURUJKakOylSx8wc10CqkZHFGNrn4g50yvTTYXM75EteiAQcHUzBL4CO3SbW2L07d39vc0
ATT9LWOkodFMVNJT62Yp9h+Mmc6QTWdQOwWI5x35jwpmTlGxW8bkABDoxZPbBraAvHrmUBQ+g7HH
eh+hAfFsTekSEilV3zKoW2TLcJranNsOykHB21OatCoh7FbtN1K3Sp+uhJG2J+Ev1llThfqFikti
b0881GdE/DVpFevPnwlmlGyBmvhdwKC7ixT3/CODBwCAe3f5sGm5WYw4wSyEAvF+FREtOD8V0ip4
i1vh7dpB5/lAlBMB8V29YMgxdBz3pTarICcmubWN+EVB0VDVn7Ed2QdIWmuDXYfenqI2U8LvExp3
wW539ariObI8dIcgmVYaG0Rne3rEqvYkutaIdsc+vqJnfPPCZ5MgdP3S3m9hJddNHOsUubYiRu7s
+O/t/KPhSxcJHZkffp/6DqWxBFkVYAHpwJYIuz0nKaPvYZAUOzkUUS2hMscPsXTeUraf/Q0+7Isi
0VIfbxr08URmz8o1PE2bcbx5XD/J1mNSbPZ/SpYPz1aLSPHHq6Cuc4TDmevw0PklVuvVHX2MOQtX
amTpmQTaST7SwCXs4v1872Y62B+9kRHMmhtwKxEePwW+4BHdRcQMsqm5azII48Zycn0e1C7KUmNb
uEUnmGT9FZASAzl0E/mgUjZmo9EYUbTWaduJ2ROlik8a7jIBeysWbaCzsX4dWg8A/1rNdmpNEqoO
XV1ladIaIkYbVPFaNriccqcgjca+80OqABxHWKky5lcYmt7jffzc3W3VQCRL14+s6L5F/E5VOxIv
nlaE4iRDKqwVdc3Za3nDaAZDUFQ9e0Ys8V5iseMz+eDGboVNXdpWZ9NYR+/bgxIpE2bxI/kkgafL
Ahl4w4QtyiepdAozi5LGUd3JaB8OE52Vo8Jh5DOXoA+5Jaa2TbLn3n7pFMHg972DVSTKpGLTblb5
yNrz5afLvL22Xc9hit8P/BTfm8uOPFiJ0W0vK4X73FM/RbHPZxDjbM+S8/QJk8u6THDmSohjFdqM
ajCBauhXuyInIJZkz36SD0cwh4Rn6tXVs+b3wRalFg/mt8xQtTuJHADQZ/fjBoC3Tm5+XjeEjZYL
Tj4nUBZ6C4c1i1DqCmvScAleUCte+c8dl4xZl0QncJA2/kSYYWU/98jJCLlrJtr8UfQ50e88velC
RPXrKdrz/x4FtPWTF1TVSFfCpZ+WxEmp1korj2lmVhXelarYIEkAn2EZuOZr2LhiF7Bycfkn9njM
JtJS1yItExCObFxupPR2ARKQJTkyV2cJU7vjEYm1AFDCRIrToHQVLz1lihIQQdgvJwE7Yj2Jv9Tc
CGex757W25/hvd7LOsD5gS8cbuOZj9jng6goCZLtALkjznfZmzhYjR+NtwahKWFfi4G5U7XXsls4
clUJHiOcOdGnnpBfMdZec41AKBqp9fkpq74rYLKK8fz3aULBIAna9RurEnkrGYz40GRSULqzRPXe
mxIfj2LF9F4dqCF/EiGkgTBBkcpaskK6aUW+v7Tpp2tzxW0LHQNuGcKfeKzO/M4B3ttyZY3CwpMl
w3Xw/k4DbyBEKVehxvtFvtcp1gUqqCytQJ1qnoth5naYGBKA3gUFaUzERt6WRSmPgY61xBougac6
uPv/lMlHZsLEYn0f3wOJyKZIhREPOAat0B2hkmty/Lack0xgwTcMHq0Dd01w6N3RkzY7Vf50vFqj
NbW2GFAFIdad3USKiT+yhU43Ci7lYg6Yguzm5QZL3wDU98QiMZ6f1t8W/hDl/POeG5sr6stAoedX
vLBlz5viWYmhv22NFI5IBi2SMJI7ISg/5ioMKmZR2Kgtgy4zKEmeM19RW9yDI7AAK6jlLtFrOgNB
e0h4OlOG9Y8fllMhRwHDwpuuYBz/dsgJjACwkoRWaNw103stOJnKHJSgBBvhcJgeIwr3MevTlZLG
LebGonaRpFsm+mIT0SPLCAOYuQtVtQ9vahOQo1kiAjdKiqcEulyN7TU0KwHQ/dKK1MyYZHxuh7p6
3hJQ0m5Ynfkn1gqbFjxeG/JbekZWBo5B0cVw5pfxV4rHuRfFPn8Sw4ZUAeGhHBqhbxpT2c9kDrJb
Q5jumY0QECzef76U+EGXVIRxKh4/PCbQPBw+DJzQPINAXRSCD06/II6AcQmznxxYofYDf5OFPaIh
0P1/drLkymE1uYM0zMEzrvj+TM1+3LcR6+0Uukl0ptRW798TaBzFQKJiOKJUb6Lb2U/5j2KHI5pF
WcJ20S43oNzJGsiDXZKyfMBugtDNJKfGiRU5jL1BbFAnldhcoMJxu9MBMdASqR2rsaDGQn5G7OH1
cVMPKKTjcycdGLXFakRv512trdNwf5HGo8t42rP0SUSp8CvlGoIGXsZZcNFq6jaf3i1aH0kNgbvb
Zuo6blbWjAIl6h2/9zZiVC1+Astxiq3wBUVRh30M59UZGBL3/drXAY1mn8JYXMr3E+YtBnatmUIp
45Tr/+1lnchsfpQrhvPi7mf/dwyf4G3YNOfVB56Tg2kR2BWfgJ9WYz+DHFBNKV1EOiWXvisgwotB
G7QExa5+xWh2WhcOkeUPvfBnd6B9/tSLp8ef3VWTLLW4qtndOiq0Nildu2dWFUip2e9TzK6FfaMW
QhWOjyk+Vucydr/PHrnpx3i8oYDYsVMD88uIbgh7+etlpSsxbOvZ2UKsN8XnGsV6WGrGDYtjGKpX
v6gd+IDT7HuKfOTRvgon/lIjLk8xGf88fitjQHAS/HdwnQaNh9WsqWrMHh1L2b2MPz9mfm2sblVB
mEcS5ye9iP5x0rJ0dGb7vvIUjclgmIphJEwTUGeTQVvugOJyWbxpLYSWtPBkBmjm2vcRlXVWNX4P
tncUISKIzdcwpxrrZEJQasGgSgJ1J/H7xV4bMjulpZTMb1LFw9zD5Ot/2bk2vqhzW8Vx5pGNYwmP
/ewUhSh7gUwe3SRsiPgK9Rp8Xqt05DEff0TVNfe89ldEvQd1QMkZYy3NOvNWCe55EPeYHGAw8Czd
IQdWvvv5HXvfcQ192ztZiIrJ0iBtTTGdL273pi90vuFPSuaz+MSUnTXownb30xkWiAxF5yKxNKN/
8BL87a5ym/HmfXe1fncyjfYSzKQVsOXSlgwVJeuyXfxxzZK2L+zd9vXbPFZGeXbiQATKMxh+hS/a
A4nwWe9xOn1SYlzAFIA54y5/fzzUHp0XRgZf8Nd111F9csF5dtFNWaM/MOxOF6eL7IrXDRnh5ZKF
z5ERTN6/t/D0Poo/qU2aMXFoUhtd2sKV5RUym1dngi6eHH2dZVmPMebAsQVhLrSKGhD3dexFrYHK
QwtU8hdMxdkMGM1HW1QWrRYXa3Jh2ccs7L7H8twlawQSzHWeYl4mXaljQwJw/4Y7HviMUVqbE3GJ
cE5G3btu9HPxkCJqiymvCa/+Y2Hh5T8GatgU8ium1xeh98gYrELKUXMx3Dml8EZ0Wa5aVBsX5ViR
Di307gB4oashLL9Dii1+Yqmgrf5vmNYwuuR4FWdRf2WdeR/tfhHETna1IL9N9PCMsQHnizBkjNge
h5b2gFXWO3stXxyvcF5CDPQBPOw660rIe/Evf5tSA/LWEnKG81rwpCJTP2YG/pNGEc46ez0+DgHt
/KjR4p8KZyNamoKt98Wldzumeii1BJxCT2eYAgQRhvhpdANn9E6JnpCJ+WR15vJrq568toPk1FAb
9dch5EwPj/0ncrhLI+CnHdWMe6fKE+0LN7BzHR+RpTWlmE6xnUTirb38De2YhmmUp7A/I3/G1ML8
v4JJbpm9vEwGzc0/u2bgPBb10dfNa1ZkR/U5+deAYzAwqYjvIlQ2Y/RdGHnRIzTZU/o6mgESVLfH
9+wJctovaBo69CTHIoT42wB/7jk0PI7biAuAgOtYGAxIySNxEfOQHpp81OEvqmfJ1TbXgGb3kulr
0OQO3Db+cIzwex+qeCAvL/kayHuo7mYUXQ9qlGaTEzkFcLgfCGZe8Fl1DG5NVUqYpX3JVd3KQlBY
gOormtz4fHu1aybKOPxbrl88lzaQxO3ft5wU29YIGfLlJy7TwwyeHhNV8PjVKuLTOpGhPutWpE1C
wZ3zvtX2PuYoRNmGlxmL4KXsViax1Rt3nF1nlc1M57Cy3V9+DSrA4uq+y7Ykqr1I1s6mZHrjCuuk
XmIa2Vy59ptfo59t7ONo0k7sn2h+gZXZh4Wnc7xKyouNyM5bZ25kM6hzohIoOi1epgDXSxLmTsl2
RRDfCMliWTLEn4FaiKu/s+95P7t4n+BGIebAxZ7qKFgyjlodceulDAPJgBBXSdGLqfVvcx8h/vhR
EA++8zAM+W4x+ZavEAPNMaxtYsyKqhQ+S++k8L2WcSbHZgWQKu7GTEMEwZNcFiJNrSoaVsMGDjnN
rPycR7kK3lGOHtEDRWoDAc1J1r2KHngP7kWnYyFNRx5A6XgAKP5pU8wpSpiIJ0znSLecxVHLkk92
SyDjsv0qhShC32SVefkE4XS0G9IVsJ5U1BKIw0IfY3f4KZ5ojfpBGIGOhjZjK9QjuB2PvO2i82tA
4l//HytWWN9jLLebMsT7QVT5DwQmUVeCvBI84O9axZrJIB+owFtS3ts/NmS5Q98E/PJOYUC2MMEy
Y/LaIRZBuld8IbAFc8A4f1Gl/SGQrA18VW44YOCI2mTZeFytZZ0Wkghe08RO2ivRmVzobATu/3fp
ZW3V1asJCeXctbFDGFmr6UPVT3PzehZXl4XBIgz1skmsS+3+0t0OXp6cMXZYfH0kE4WPZXicurgB
EG0lSEUZYdLWYRiMM4jdK+aaU6zux1qQHYLE3JgE/SLOFs1Jy/thZhWkrmAv98h5gndxPpYtBuei
Hyp29oaT2NAv5VLfwNhLY1MlQ/vZty4PLVkwe3KrJtJzKpvbSH+q0MJ9HkACzn9D7myHyMz2VGEU
xtociX01fInW2vYMbVE6f1WbUefdjsQGRn/A2YMtNQGj8A6TRuXuyVqLr+mHDwlt4E7JU+H8yFJb
gA+L0l0/5ge864csboZGHQm+r9oDoJx/gc745vaBsBWMrd2ns1KrN6lLS/b8ZPWC0Eo0u4QqEC9a
LGFEgN4ylfty80Flm6TX9MvHFICUras0dhbukGAhbne5/fphL8lLgDS3juXjPAxarM9kv24QB+cc
xqVeB1ZrFxPfAAMfPH8+ZIf8E4maoliDTlSc+YHTBAY/VQe6cVuatuSzANzEU+jJYPm5E+rZexn8
dvqTsiCUXEQO12+CyN8rBH5xLZSPXOzC8QAbKJH/sXQ9g2JCS3pY+FggWKg4JdI6t4CyWV6MXK8X
iuZDNQPnMNa1CmtmMOUe9NXOewXMgBBICJmZFWLCkYaLJSWZwUk4igejpaXM2xptgQ1ZIx08mltH
MbTwhHej6+/Dx8hRZsN27dacL8zxh30bxr/aTjJfLoVDiFTO6qKJB008xIdTsSG8WNcMSBvSBVsX
Q3Q2SpsMLRMicU2HMLYnHaqixwokYxMFsRDx3zdvdY51dYbEKlWHoKR8UWCi44oyDJIs7xsZymr9
qLuvS7E1lrCHcHieJlLwYtWRCMar6mpflDoypcjjQlJExw0hsq4Y+eDW1enTpGUFBhUxpLv00Tql
zn7/4x2fMH2auJZmh4u0vPip7F3wN2lMEXMq2JWSQ2e0yPo3f4Ta649ta+FGL82Bzg539o7Pi8Ts
0BXreI9UwJZmAZ6qC32L893cqobXOoWDs+duUYN4ct3RcjhQHWixqEIJI1q/KiObzrwjKXaswbkp
SVGO/JMerOh9VK22u/HQ+BjXr0bbWE2E7HC/Aj2nl7BuJYwQ411HwysYmKFat2gk3Zj59OjYjaq9
ZgZBZLpZgn+5FFoMG5pArfW6pdJPodcEj5D/CF1GGqQIMSkl6ZymCMITTTwMm94oiiGUcTooYdSG
VbYpY+OVuG8zgjJlveR8w129qJFcT5Cab9mEYwoXtB98NBuXpT7GgxfxX4KDkrQttr9+S8pj400I
jX8SF/FAzIr9EehH31yT8RmtyIb3j7UoYqOxDV0KinkrdZI3QncGyMXtPVyr05/sY0p9PBWpydSY
mIAogdcamVY+Ck1QSFDESLCrDzX4HvloA4wWXiolckosoaM/S5nX6k1PH0bRnJtusy+lRF48t+0S
Ifr2Y/pKkFKXAKFmcfdngqjsbaCQNTa41vp2gokvUYi8YLhhPwCWxMDm7IYfh12QfR6kBUd8bFQk
PqVwQsyn3mAfEVAg+nxMvr25K555MRwtbu6rJn3T/dh4E7Xz7wFFhwl7A3fs3L3PSd6tDvc9Z4CB
9jLB1YD8pq0e7mAo4ym6tY20o01mH1YOYejTCjVbxDFrO1YhPkxP3Z9WxP2DTFbqdsYswA7LxxCG
oA0xc9+VhPJ1CQOOcLqCNjPeyTBxAfWuoO7owkF5Bnz4fNA6mmofjVEm/srnqwG1MueaTP1vhTlW
u3UISLiQfc4RrVFKqRxH7WWmIOdM9c8RYhbnE8p6L/jendDeEKt5SaKW9ggiAfdS7lkzpKIpZcov
oQKB4B+Xm7IFO2X4IlxRzpd/Msw1UZOK7UtQVVomnqEOXf39/XsN65uu4gF9xB6U5Ogt5D0uld+z
TaidwsBpEJUibmeije0lES0uPl+0+eu+lgSZ+CLAuPOG1gjEhIho+N8iF6HmLicRmAOFjUBV74lr
J+wGTvvmT3j2NkNhcSjOH86tQY5lr2nuRDGCQzA/FEFy0WinW1w9YetWx9a2xylGVXOOBfpUiYLe
SaZdQj+VcRr0ANJwWBaO928kZBOLHc5tCeqO92dpijc4nhgt3micXNRUH4IrKTxCUI351PGG8d7J
WgjODxs1UH57Lgpwvx0zA9bKAtSwjH6rx295OlW9J5C1t2ND4f4QhpL40uumTC/eXf3NLc8rmi9t
8f8DkOxQySRWbRqmjEj1cw/imlQgDAeGxVRo+raYmSbBEKDtd+roUwh8e6I1o7scucrbMWPYcLFy
7kWh9+tnqopky9cm621wClq06IRm/vknHpTwk+Y6i6z0WaTANtNcu0Ou6uzfXazM/X5NBij79UEJ
p5RppSLjTsCwQxfhQLGlWW5KlsuYAiYknTvRtxRoiwFz4lIGylwXJF6C1kxim64VHLIiH2hooH/v
Sut9tfvl8U0HCH23T/XQGevOGjYNAD5MwF/wB0WnJIBdg6SsswJPHRVo9XAnHx8LQ6ianDyypKV5
Qh/sC+Cfj3PbV6BdPr795lktc2u/3LwO2DO5/wdAxIFn6JD45ZuiOSysb6Wb9GveAnurz1cf/9cx
rRaL78sP0V2fLG1A+NFeYDS+tfoHwP//98iSQs2EkSHhfRY8/RqszX9v8oIGMmGMEr1ecWE0nz+G
KGXgNhGj9wqywcZ8Fj3Q408HkAszbo0RoW0sMjVbSdTbjZx86Ww6bQD6sA5u0yCf2AqVwWppOuAg
pWFV8Ac0gfVzDDFEovII0HCKUllrLU3dc1IwRHzoYXz90xPFzH+Skd3wyTaSpo0dM9CorOAFI/am
geS8T2TtEtkj58h3kJ96JPlXcwYY315buApJaoWRwWGeSJCzydFn338BKj35+4/tKWLPc2XGd3Pe
Wwn0uTtfZxYL5eqRKbnklI2Qo6wu7xI57WAlv5MygPDXAPCMul22fBnzy8fjHh3wktxcJa72UeJo
KFRzp/CS8uR7CD8dGfgMScfJj66Co/DVnP8AwEF9+0wSHF9YN3sAeCDM1+Sm3DLDpmQBhMnt5ul7
FE4rwZfrw3QIPRkDpJ+4w59XdJXZz0PC3aHF4tpCPYhsej8w7viI+soxaCdS4Gtas9jT8P8RKKdi
kN1daams7U223lFTEOni7NL19jAhpVnosMjRjUpP1C+VwOvolb6OP8ilww4jEeeYCgIoYnDldYj4
0SKk5VZGCal6jr8OrIiZL96KrppmWxBnrMdPEYeKJQHKFCMzdv9DcNtESWGzQrk+L/r4Ml7ffrBZ
WcBqDNqp1jdjj3ese8oQCPvb9RWTVCtFPocitJqR3jdlUebYc/pSY3YUL1EDaK6wKIlMWTbgDk13
h+Dh4sGRk075gxpr50xqwHKV/uYS6gZdU7mznyY1NufXeLmqI0mOS1oZJ+hO65p26d2hpBKlrlfo
7VWZkhOwpdp1+Ryd30WPDqPZxdZfW7wh30OcRmazxKMx8yyjx9l58N2P1usZbvr/xxEWxrgBy6/C
gpywkig9eLkdlAqqBWQtFFe+a08z6vFFa35lOXafS1wnRIIkWItdlys6SclF9PYSeanYK0rdjgic
TiTs3kzfKJJBsorSYpZ+2PsiuCrG2Gt42F3+vxPVoIxX1Tm/XlFNQqu85Lf5QqniJ9gASsp0Hv1+
l8Ce5QkAHo4RkvBv4kYDSsURWBwvddXz1M3VTkdHGDnPW7IqJbVgdBM4xgvViITOkFQhxTUV+hSK
WPwfUrD0q3U0638fTwbr6ACXgJZMGNWpAyRqGqt4V1GkjSvcAY4upNkBAmqBx4kqzZDZVujpKJDa
MEIHpO/7wYNItjkP3F+NbqoG0TENlTigNsgCrIS4eLW9uAkZ47rF9N36xPrGy8QSyZpNCwGFcz7/
Z0hRWxjO/1AN/qODM4RdhMBgPGxkc/OvtwleFvOGQXLVs0wifWJrjc4LSOkUxZfjT6EvrWlj/NSI
rWZSymypIoYpbxMRajPhNVJZ/5piuTAnKxEP7T/mDw71LZp8qKhjmD59WvCCxHE0OwkwLmeZ+tHE
cZ/0QykpVyeyXZ2kMGkNs2XKEB1zvmHaRSGSNF3jncob/mzojOMbyY4k96GpNn627hYJWjcdfx8/
Uv0UQMxjyNUKZivwS2qVCpD1URJhJzoLsPhVe+tL9UgxUjSG+2WaeajjW7vDjVaBciVcjanMMMiS
albq7+h18BtxXEw9Ynyqnaaqm6pV5LDKsfoKnBiRDfuIpVHKqZ1jnSBweOMye1BQtiMJpAmRD7hq
rpqUf6qG02xa3sirEuHl/Df+tclJPN5LsLJwvfceudspEH64je9Qa2d/xRw300F41dA2is3GcIiQ
JVC1Pj3amE2DFEKAGsU0j1IgdDlwIwvsLCw/mkzKntbok31/A2h0w7RoaX6Lp5mvKTdF1kirJaJW
Q5+75xs4fYsqNPXhxOLRS40giGVYryExejABp7ETRPc/g1K4X8g16GPamRDOuUQk9EInMpE+B05S
rSWMnWU45qlDzikstrphBXd1QsqfLaAMctnNzrsNqS/JMTewTXKKFhWHpNcGSltRaHzZJUuR6Qt5
VixozNNlgLl9oTNiDsBI9AE09Y5uqtUMyj7ClpqhnUXTvPOdSpQCTWzjXY86rGdg9Y/o4HaKCjpI
zzdpFsZHE3+zcfEURAKM8TtNh+q23IA7HAFv2ZReUeiqiBTzlgdwJ1IrfOSTzvp+tx0lG9ckHpJ7
VX3hMtej/uggzKw30n9byd3ONzbIKzYMwIUOEKOaOAVJbVc2StDN2wHsZNMBSmJw7ll20r/IUsGJ
v7/fF6VTb8VTDpCW6BTJJ4l6ueozv9zQHFjrChuFhoUSWFFooCaksNXPD6DSPtI+kqLQ5k1rPwBi
WRjGGYK+EaxROlo5wNKqPK2OuvssI+E20tX03OYvhm7vT2ude60vq2uikUkaXW48RSPhTjPk8SG5
M8v1mpoix+eJipnXhbS5ufPjMIvC4ho7epRaCxQurmjKjIV+09Y1TRjYFTaC+SuHiYl2O1bVZs0j
CgoP3LZUbAcLvfWameYk92tBqoHnBvJZIv0am1DWe7QuC6jhCMbJBODXLou6zMUOidSC1VXa5+C3
LHIuFWoQ8QsS6Pn4ide77Lv0xbLJHYKylbJzC2x04AWLatO7oZlMPFQ6cg90lDaEqg7D3VVKlXh9
iEVgNa1rleeZLVsN+kwdsMhEouQlItb9ZNbGUeoy7ODpQ85ABbPXwIzmDinRHzGjIcscoVU7rYqh
Qg3u7xcZ6hEb9nYj/JkQSby5IvDhvFu1qV9OCrK9KKC2C/mVe8KoTggNwtnwoxXYR/20nWpFMDe5
1+HlNta1dSTOcAJJmuTixoLNemuRtib6SjxzUkDm8FOHtRP3/zpKuepgOVBF+6CG8I0GbiBAwN9h
GInPSDaSJtUd0dBraKWjku8wv6QdSZrMLouX1DCDD/K1yUGM21awOYVwm9jViC9KAwZ4lPGgRX8x
92I7p6005PVosZ9U4hdWxR17UnUwj4H1tldN47/JXaL4s+6uyMCRz/WvojvWdpNYXc17E1f3IaQ1
TK6QY/jvjk468mYBqkayuyvf4N+lNMGfF+gRcUh2XGs760Dg+Xehcyl2vcxDG7zEHzXeshMHu1yZ
5bWUO21VZ1NBUPpUco5/X/YnBsjH1TGtSYMR1A6mBen2vCgep48WE5uq9SpCC/ni9eCy7NOYLr80
BD89mirxd69S96ZQWyKjl8H0KkWEDjnbeEmohqpYAIPWeqtZcUsKkYsTnZAyaZWPKTYzJpdrFlOv
CrMOYn8TVBJLWSNRqIZHCa4lOvzw0HYWsbQkJmDL9R2uT6Q0jh0s0KyKpBS1upZuK3qtgUONxfT0
kLRkwZxxZAZos+X0Zq9b+wKZRj24HQKgI2KNUqsIa/+nMeScpMb0wyJDVzpmhSM3KJX6PU+nxl3g
QE4beGxypJDlHzvHsRG8vW9D/RVztUBjJ7xizjwEdzS3kc9U19JShN4vOnkVM4vRUVqs4EeyPdrx
gda0Nsm3a9DcGrmf+zsxK3B9N9uFYsa11XAkXdDk2E0wPL9pKlvpdgms7jQCo5FkTQuPabaxRgVK
ggz/ou+CFF6PMOt6wxWW3GjpGa1m3fa9KwCm7Bqc9FqyyXHBPAWwPLpqKk2e6S+QYBYq/T7sdl1Y
cFYt5ohfoz0bdxX+cZg/6Lsy1kQqHQAUwOmeWQh6KtwPiKGojOwN1w3sgbRnh3QHqW+1P8I6UAcn
i4O1xk4WGJyiwzA05U0J6HqwKPf+/4SMRJW4KbqAD+h9my/zB08Vk3USjwKMsS5umWEv8/J6xoet
YdN8EW9/HeJBFU+Ds33lZk08MBfNiRMIXINoGT1cnjdlVSs7c7oM9FnWKPH34Yxdji3v0szG/N0F
VLnYPOmrL2u256DvvqzTTYPvwqzPv17P4ikqtTdZufInJVMry+AfHf6xOeFgWlz37BtsKnxqgol5
OThnRy1VDErPLNC9aUPBq7+C8x2txfPu3txbPgvxETbh+UX5c86o7Oh51GqkCx5It81K7h3Kxul9
i5jXjjrR44Eeyq9aZIc+KtojUVQ42zmEd7UtePSEi5TbmnFdmrDHL8MDRGHzaR5A4NWuAE8srGh4
ZR66PjZy2Xw9cHSbmqo3e9ipbd9QDE+17GZtVMR3AkqeSf9KRFeQJtY/R6ZYgEK2ya5Nu8+qkSva
+RTOoaY/QPPQr8U3hqL4G86sJnSBgYTAPIMk0klgn0YZCcr8zoanOPqd35/Wl9rBF6Xts+h5ikAL
qxdcX1fvNaDn51Jgxnd+Zuhwfq6GDPTwqm1EG2ewjHP7MBlFPqIiKOMexi3Ygtxmw+IiDNqUmhal
aKjqIYNJbmXVH8ETLlhk3P/xbgTD9vJtTD60HltQKN1dB0enVWX6GzL+a6x1yrhpV8aXGPQUwK5c
IuGNSMD2m0UB0H+Pw7AgGcd8TeJgRwcoupFGqiFiEOmV4ud+c1MtZ7eojrJdJcK60nFfOsCdo7eA
8DNi0eJgB0+cjpZqu2OGW+qKX/vAnaVSMtWM6D1/xaK9EoLIiHNytybx3N1tgAk0Ng75nunMhCfF
ZM/a2FScrMuJwVmt6Av+bhxYI9lQAjWETvVLP7L8X/dNl30WqKRR1Dgt5Ru/HoMKXQ+gT9addRsX
goCPUfH0fhUGGngA8T1X/1n6k09mWZXxaW4DiXD32KV1FG31xLGquKiw2kwBWoKCUX3gq9PROBS0
VhdHaJ/uycWuYmm+G2PUKnEwl4zbUk3xdCJoStQCiifz47zbwH9Z7FCAw0Z2w68vFGMBSL3A62xE
1HeH1gFbYe1STbv4aH7L1mTs/YKiV4+GogzvccSRIy4PLwHWYJBE9J+kA9DhzxWH5jQdJJPT2ox2
EXZNdPf7nWhMxD3LTsg+NGuLzuZMf17zYVsB4oN6gKNA3vboUp0FnXDNtWa1vv+6eCNAMXICrbJg
s/QmdY/5X8Kipz6gf2Q7S6+lZBOzI5Irl+J7KtjZcu6rPmOCZ0antRENN0IbQOswppdbaG36Ii2J
MgUzd/3DeQcz1b5F9RVjGReVg3MxmKgl/AVZq9mn6+6DepaC/tbDT5vhh5ikH9N1Upc3vqhPVlV/
qETHqTtTj0Uy6RZZwMGKDPg6a3dHuOFEmY1GIzXVbXwI6iDaYI0TjGzBh3RmvYEeNi2p4PPJERem
+SbMPGjH1H7FzwTCuWSo65mxTFPouov2i9BdDmYkNE7hkekjLe9nZrUE+u8JsePLk1UWxHGsie2b
wmS5sRo9bw3so/1DAqnPVhyZQzaIBlw6odQcE9xHEYdeviySIgjlLydIFnVHpCB1nWtR8rJoIBwL
9CeiMwKfAGPBMEkdDEoVYgjBjAqS5Kr1dhXvgiNMHbohjoYwsHpg6/JZONOBx39gD64ofpf0gBF1
ptg/t5eDiXGx4Tg+CsWpW62SBMamWap58YcLkOyNw0wQl+SxSZ+bzXFFWeGPhJQEpW+qwpXMonoc
v8B3Yt/qZf+hisGezhQbN21AM91SypIpqQId0FCvsAocxUbh/HXBd/z/11EddrYbHnhMTcthbZNN
BQy+vEo4NqXU85SZRqmvHp/7a8sr8obKeTkYNtJwv6yrWUbeJWxHp98/Rl6zgVcfYA7lZD59uF8x
jzsLgZbWvHWbOVrfFaWKL/Vv6wsraqDrfLQWoIIdyF38IQ43giKh7PFyta14gfD1FEyLQlv1VXY9
60Kb1Wd391Q1aDN2uxqFeLb8StbLbHCqkCVHUAt5IS/lvfd4FEvHxSWTSbA5sLqczROu0jdT4gao
tcUYrU/6jHFXAYk3MxHOQdA1C7LTIZCoWW0b7503rtpjtyIAFn0eTbCBgZbO5Za8yd3BTuqhsWYK
GVO8PE26Sc0Cv0foNBz6Gu8hSYuz9MFZXM2kyITCZ7yo0h628Ei+soYha/Rrk8WE6AhcI+IblRAo
vYzWWqr85H8x5n5HhmT98hp9O4RVjD4H4GvAjMkExV+0ydd3aBrXYf+bj4Acg0ZRYslkg7UHmTMB
XwFnUmjq/zTTP+YlznCmy/v3DRAmDzj1bi+sthg4o7BpXgwvkpyMIzw3qIrBYsOdG9xKZoHEOlEi
dJw/9S3SeAnxl9g8QqMey3nomLi7Xf9cVpnw4Aq5/ZYzYJJGahMWoI12Ra470yMD/O8P0M/x68FD
wP/he4R6k0Q88ucQoBI/vmIGusqlVuXi+Mm8Rg8MPfoKhwYbt+RNM0kMKT1K/kjRVJa00iuquKnu
y7A9bjarFOs02v8hTjKIxkbzD6nVXUOCXPCe4I6mPg/xI7CZO9bGgkmAxXTG1T9vmqlalNt0i2mq
jD4umjOsyU08MIO3muGZ1hst4TdDGsChpoWCe8YdAwWTvBz058w1/JDVVQUkJaoanvutmDAH6ReS
GGnnm58AtMq/cPoXKeiRgQRNDNXgQ+7C6IN4Iut/NrtzEso33Zi3EwdYzcTmDHTGE4ZDYhjBRWv+
vzZW7KMIO+MaVc5KTXa+Nv5bIFXlCci6ORkOXtV6n/QfLh5lV5wvPKicv7HkO1olde46iCsFPNkF
BSg7WKtOlWT4IcLp7Rm28v+upPL875s1o5YAJafWZDYafsJhfTU2e9P+PLJJdCh4TnBHgi5TtVby
f0AAEpa4hiRdTB1coRaEqD5/pBJyWmwpc6XDl9Fhe9DgS9LgRMzqcFUwk2riMTPW7P/Y0mpaDxn5
JC4w+jXAG64zyzKfeQNIZ2aef8goWx72hqe8QRSwrY7pYI01IyI6Ie3QQ/noC8fxBKyNACcvgrfl
V58c+uPxHDiF3x4O1Lx5nA7aDr508x913u4Z3Obgdc/M60QLzSdnTHLjcdJ64qBwfJ7/eeJdrEQ+
aMQG8nmZargxQYxIa6h3qR65sLIzt/0BJBuPHYAcO2aWjO7u4sndDeeLwwWpokIwINwdgoKGaOma
8tQ8mupc4nVxlT3+riHUOqCZfWFVz1YFm23Af2LEiwMFspV8AkmvomSOsveocQoOCRotZyExi45H
8YshYLnC+kv+GFZyGSQQotSXITu/Wb1zfaEQRNuV0u2Vr2PxtrZqKjhydRXAAPsDV0HOW5PO9vHh
6pWCfoa50Zpq0yBLbFC9M978g0qSqHVjgoHyKZ7epTernSEgWjdYB8nXFczKIw7RovooEgyAV+15
Mnqy2UlYa0tjTEkDbPxhVN1Xo3joqX5MnyfgH8GAeHNpUPnVuMM5LMNNSk0o4JyJOf67h4pecu1B
0xAaqv/WnhuR9cV60JmozcAoJA1ZVa3o75PGaUSQkLSvklBksAed2KI36SmBKXyaceeKhtzSQK4J
qsbvvqmhBjE9Dn5ZLvI1RdM56LCYwVWcQJOh+GBShEf9y8p2gGNm92uon4u+0MwlXtcE4I3sTsso
ND9bpKkyyVegGUShmDVgA4Ms8TfLzBVUEZMhyU0pbE85YCdKatI4haTOZHuwZZU/nr28OAroepZX
cM81ACUHQ43B5Dx/dd9JkxU1xk4zlybtNJ3z2nfpi1dDPXdyiXMMH1SjOUaIAoqtApXt6HrrrY+e
PDLi8dNEkbOoVLfORgWJfdS8DFb9/HFYya9PZAfIK541jm0qAriW43TV5kWHHuJyX+Xs/kvSugNk
+CpBZwmsoEGdDA45U4N0md+lDqliiGEI0dXPMD425Fvr63/vNuVOFm2saWv2nkFIQ7F2N/XfmkA8
rxc8Y1yDBAmmLGIKBFojtNp8lYNjmGPZtStDWTQ7LvWP5KfcEM5IJQtbCg5e+bWlp1lcyZu2Lq9Z
f1XbRleV9MIcaOgQnSmEIy9Ut79NNVFjn82YXetbhb6UlopDZkv4n9OLJRXf5gK7JGTLHAfpGJAL
LJppGOjM6Xw2OA2VD7trLzoR45PTk91cuQIIN2HogKdOPzl86BnTM0ld9i4A5vRiwQK6mVPkeuaQ
BHyfAOverwrzBNxM7h0ATXB0CC5hknBPDXB2QINkEouiXsT02xqYhbyig7pdz1L9oE6DAxyDAs4V
QDvx8YT0cfzRkoZ90a31BA4kXJ089Lf9qeoRQToRR2FuRERnw6XXWbYaKhoJyYzyxeAh8NW3eoCL
GEQxW5WnmEviOHr+CsYJcPg5UV+OKMqp4Tn9EN9Ca1+RFz2epSUeEAoqMUZQgKD+Bz57Rc6Dqte9
BIoziRgRPRf2fmyW69hrZ/boo65J78BH3LMRtf71LsOfwto1vfFK1YNo8FySG0m/4Dg844/4JFHl
zvgsrUYhrquQMQT5VMBHoIETn1n0Rj86zXlAtpaW2ksZLvOypmhMDtCOu6/nfFAfIamuWvEeKsHU
p9gtmhTSjyU26TXvWJ/kL6hFy0iSimcfif8gaStgHJVeKt9PF+/XIZlRilNciQJ9m6m/ZTCt50am
/Y9ZNKDGbHobt8mMhe5vxZHmtwSevVg4bJ7g5bmdDBL/TMusAsPMCtmRsUkExErMY7lSvtYVUEmQ
ZzzYhgyh8oOADDW0GpOMToFBXh6/h3qa/tN+Ibr6PbfRLK+VdZjKtaSiuAKP1O6nJOnNw1NnlD8A
6d9cjRUQ5y3V3rzHJJJyl0YlZBaDASg+TQr+7Cd7IgM8vu7MQYFo+NJ2ejkxxlzaDJcRruJLg9od
4bKe8TOMdFOziC8mH3noBh+UBaGN3Km2iV83K7joavl/5CPdn9DK08bgA+jtIw5U93Lf9Qnh7gTn
MO+/bI5j/Y3WL0Z4otystd6b7JAKuWp91Ci93hbL3kqvsiiNMJCOrsuzMmaN7WApRcGelHOG3fpw
l8HpEUmKmSL3DNit1e6BLNpOy81ci8wttbDSOqjh+FpdBy0tW0DlfEGavr7CTHRZPHHIx2rGGwFp
7u9Q7RHF8sU8P8ZIMnuLjE0laxul144DRsFK7dCKPXHPFWy1aNb5cDCcKTFo1o3nKMNjyT5sOqVD
1IKA9Y0YdE1DYNgL1Y+C4ZdPCnHCoeoQV85RRomnePN0NLd/MU96OzUNNHI6iTNWSHbdiD28d/ou
UmuuWfwVhoW98tCAmuqdcqN2Dt2bvDkOMTgiiHyvUKRik6/SAq7v95Upx7FY9q3X/99QAA9qu/xO
8bB5qPyH1aKEw+0Daz81VoRI2LcrvVpzkWfOX+emn9ahfKHpCyzFPch0BBMOp6NqiSzpoke8CtGF
3esXp2ldq3KoAKAgr/0Cmobjj6vT0Bdy+Htw7TMTNiTL7PfK5QOj3QHR6NQ/nWcgRhOu4AZpWxK4
HeSZTCG7jQaT5BHtb8w1fYqy3jDQ+wjwyjTymp88jq2/zISHQzmZAScsmTtsHiTlIRDS8wznfAQT
L+NF8Wfqiwk1od8QclLEFpGezJCyCJtJHM9pt50HOkABi3FsmLvs64npMvylwawZUFmBvsq77prs
lXVgurIiTPb6xAT194SeuyQvoG0uXfYx0NeRIa27dAbJLuDLSEtu+2bT+H/x3eaGvSLI6k4JihvP
9TniFCAIgiUFW16gZKug9ZFbnWPWORWNo7DmN1x2fprSM9c4qMGhPDUuVoonZ4kaQKqqsq53zVUJ
B4nN3GpdF+kPQxUayBzvR3VdKTJa7wr+UhFrE8GPqAvQ7tdaqIkEOunXRmh66nbhMVApOy3froGD
7ace3hh0xWBOR026sgoGYfmzFDnkghblP8kiQ4Op6eiU7cyEZvtMIExUKlO/HvVvtdV05ZqV8QcP
C7djgqeuemLCUKtGInuo9DK1cfd0fawGF5qZTf4aJxKH2yBVyMjaAoWXq2GChUPtV1ctiQ70NAGF
Ee1hLGniH5+xN1N7Mk1I1Nl13FAhoLvFhTCBs3Tykx8gGV3KVE/ABvzvFzmoOycLvRKp27vkQ5C9
3D0e7NYoFBPy0MJ0GWhSH8dnOHFNMfRhu1R910aTUCM93tSk+ahoUbgJ+X/1STI5IcwEdORR8Na1
eTdVu7+p241Re0wB4etzJEafGFRs2Xw9Hcw3kcm3Ijhwec+Go6JPaKnihwZtAkG688RsR1nEMlGU
NKBSH91M9DGja2s39YPCpYQtpqp9vLbGewSYoookyV3d+d6PsjMBaqzlJp5+dT1ryv0HGEjxvrDw
4HOPSZEfa/YqAyImeFb86EZfA3cirC+nEyfYnPnO3/GfNRnuvecowFTp6MJYcZzBGL0reL3MKU6I
FfcVVsKlFBGSq7hsMr5apc5e/3WacSHIBvEEhbxGdIvFJnyrQXgl695fcXoo4UWNO5lfRmojH8vf
d383WCLHmqhnc19c3PGUjGmcJUYD8Tzn8QOFQ1JP89YvXfJ5uDza6S1xuWINMcUwBQ4Qb2qel4pc
qexSI7DE7vbewAGX8U0W6cuH/zEE1ox5FECBnAiqAqQXRW+qho0dgoCnqFgZU1RFdRms8mQ5iutD
DiPYB5O43pkPIQG8RP8JyoBUq05FHsAzR6+RuimT3crnr+UAeie0cxVFhojoYjV1mhvvyeHAbRQG
0uYCsTuHeW6hca/NW4QObXRhtNda9VYbkoSDvCt3/7t+hU5xbG+UBmRJiv7j5w8rgZWEm2pYdhBE
NAWXIQXNhS9MHamHaVC1EKJiC3cyts4fqsvfZR4/x+nQYZnAa7M9e2sUfGT2gy38yEHDlUo4fql4
esM3qdh3cdZM4ITz1uV8C5svteSJhvXGfM9JFs1MQFKg+wWfkGSyMFPfpYxRp9Sf3qZp8heSTUd9
OoMr8MINEnivNek5zI2Mh3tdevMv6ZRX6bxjFZFKENS98QIxVfq5/gc09XL23a1JMCKSrOmNFfM2
R/3bdQPAhv3WO+2DcTB0DOzUEYZssLjhbx4klIa9PI9qGTMDCNc0yrc/CkEmeAeRPzsEOvPGrzsu
o1UTf4up04NgYFe+XXbwGaznzGax8tnQVF0KNvChqMPYiwwFpN31mRlbtAVBes4kXbdmgnriQHom
nYWms6mmnFhX75dxBEH1GvHwodRnasrYuyoEsZTvEdVTxTP51BdqMBDAfVHrBEEZxaqKmhHjN04f
2dB9WzF0vNVxzYoqpiC0kvXwBttiESXc46yFodKBApmTvrylhIlsxTt6B49lnXRl1EKMCinwf6DD
olCy8OI4LOGbXt8iViXLH6pN+hkF31QgAxiRpazi/3XLUvuRugZIKNWzSRF5ZvhBYZ7FtpbNG46h
/Y4xWmfabAZwn4vm9XQbeyQl5pgsQnfcKHYaKbl+LwanlZIBJ92ndeoiNnIM6/9cr6YuUVV83yOl
+ckN0F9KvRndAGnjG/uDlUllxGnHO0EW/Nq1Ne1mBi9o/8yjgYvN8THlxDrEpKYRwFHMSYsB4bxF
dwDWsJpmVStmllQ0q6I16mmvDp6Dq/nYbo3uWa9jtzEUZsC9fNVR/rQ+mJpqjVE7LBzY5wic2nR/
V6RLQaZGXPSp11a5wuRL3eiYNEnIBpXicxQ8pyZwnItdI900s9X0Zt9wGfDuZn4bULKCXkWlkqpA
kYN4NQ77K0OIoyKebvYvxbm7d4wNOonyQ6US6xWKe/sBnJKZtP/7K8+fNPUU945znt+XVMpUzDcZ
hFCN7DejneXpNOEv7lbmYHs77tGvNsjMDcxGa3+X3DcH6XnsDHpI+nE8rhC1pjNQ4miF/qv3nvmE
g6In6zVJIL1HJfYU5payaQacgC7iN0OzPFifx0IZHgVncXqTfjwhVLsD55rlgO4VRT+zyKv4IkAy
2ctBaSB0crpWrKqvyns5VW5sWFqyyztJONRuJvMriorX/Qk6wU4ykJI3mZUmrdsz8oPexULKalkl
wLxle8UEGxrfCdkudZvwU1ts80LVXotsisbblb4M3yCpIr5y02ItmsUrgVvPDoyNNYsbTbLisR2G
6q1jL+gfuTpnKPC2HtSN67lf9q02+zIe3UUyqil/ITdLiAsO7eaeqxXFzH2W7nmmLbyIj4NGPOCe
m7f+H6H1WsixIvfomP2qcnak/VY+hZYYBqmY1sClwi7Myq9WV6M78ywPUDIGoRZvpNEJou9NeRlx
KK0+CoJE99TEgE5aC7X1iPigjL6BwdxIDFGEJNsDmWE0PXP7OydFt2rmr2OS3QfDAra/ADoXKcwm
FqmBgAJ/Hw3Gii9G8t1U9OTJmBsRPTgoar12CiIRLVW10/J6JbS6hTFXKUM9ElL2dPGUfa40h7XE
flp39B1zbXaeYs/brE1uB9/5xXGdSgYeJudvALCZvEdG1dUnR8kQImjPJRsz4VGXFKatZT9tEk9H
4wlgabyPA3745MJSXRXBTR2efsiBLK2zvUf71NKecgwkdI0CcdIv+LPY3utvZVVf2hCAOhlsyhqf
8cP5DX2jWscXKkGl7qvfoeK6QlZfUbiiyGLvN/pypkyhAWK5x8rPbbWzlWdv3qM5Uo+T9zViU2xX
Dq1PoUGV0BOdvzZ6rtjnLzW6FLaBgfcrwdP0N/vspRfFVdM+Dp5ze/zajngXQ4LwXgYnbjH/42Bh
udWx4TQ0t+Q1KIZ3MO5ean8XweSIlefN8inYQAJ6UD8v3IcWgUdUl5x/qvxTHYLslG7CyXwkbRBK
zDvNdey5x9KH3Tq6OILnWd1NDp4GDcBXlF5XNKxB3nlKk3rnLLDVfuD5CetwWo7xQQLgNc6irwcK
+KkWRgNudH1FFE0P7CSs0p4qpZ9ZIixdwME6TEPfugVqtckLpFNQy2BCWAVayKkNtv2WFA1n//cu
gniz4XeLdIEhlZD086EciAjhI3elwGKtTGPnHTVW3yMiXEer1aDMQLP0IQ7JW2Fq870a8zmKgpro
kfJz45MHZ2MMMTQLo31iMIPvKScvpENIV9Kb/ToKuQRZAbUXB0/qljsJRDO6EBBXQ7d7fxEkWRvj
/fuV4KQwk0Ctx/arpoFBPPpe32qSPWx1DVbXEoAx6ejoiiDjyFtEvRvA18BA5IDs1xNayvi6a06u
49Y88KwVL0W765V9f49uC1J0xqmAVuzIKOMH370wlZT5a/cgff609E8dP/bgweGABxxoXD8PrSKv
TfsQSbfuj/ikJHwqwNf9u4uhhfkIeiDCyVm1s7Ne8naHP+zz/9+dKTfXA3RwcvORT3qqzQVXwRsX
FOmBgcjGktIjNybPOF1vmDOzVuFL0i5jANwKvWyHkY5ZVqZib1O1Zmc88MFXw42DzkvnMdND1UQ2
Eo5SPjbsxL/RMfHznL6yFq/gm8x/6YHL6yGSp0OEoWQb7qqEQhKNclJBwt4VsgOCeWu7pCM2X4l6
2Pps+wl2IfTe9D9nsUs7u6aPxUajNv6dTjCHsy15JneLW94Oz73KW4UofbBWTD2ilziOJarqlCQP
muqB0ZuFkp1DlF/ILvzT/9dFnconLAfQZEwIsZq+wdsLgF0Bdy85u058XDbItxJ8a3+BgNlXytF/
nSblCcO2EpRyVRR3iL8+4zo//pwIRPSCgbnrLqSHtHCYjO7SpUkgrbekMH090SJcE8isYBoklkVJ
lZsnt5wuZS22l5KEMqe733ZldRjXxWZEGwmOOsJVdqXEAJZSfZSAMIZjONCWLRp6E6vKWI3UIuhX
3Txs8IEnjSf8s/OdVJ8//3ifGoKoS0AAgZ1j+thuyirL18krbLl+YEUvBVQfo26oM0IqlYRExRQg
mcXZ7V/UPTgkyPyfS7It7HQs24r7ZjVktwIpdgfCl7oEripc603C/6zOsZvMqYDpwxHtDaipfY6Q
1DKa5QexQqn47AOhT2ZxoajyJMuToeQKnR4fyI4pyTzh5jjIGhXdAbDrmFJw5dEuqVS/libycJNd
wPx43bSDIBEUyccyg07KcLqeIZddOLGtLuYR11f22h3QXj69dVGBCxl1obub+SUIdCXf+T55YFY7
YnOYwzmewUcNy9dYorvFfNNv6uT2+Fj8dqPJIvW+PkD1ENjOFcHUvilpsFBTTqBSgd5GDTPcq7Np
Q/Lkpgt82DCdT91liLoSuBZiEfbTxSNkQQS4/esMsuj5McNtCqkCQLOn2K8/9HOMGwjBzCYuhN+w
pkRAD8cwvFzl8yUA9/ij7kHfZDmQSKZIHSe2EO2Fs/rp03DouYz0zQz5F+1MSqhQoGkGKL4PinOA
omzazZo8KnPAN6xPZEmZ+GpHIA948ZW9x2xgztopiH7C37iFYhrQLDSFSEW/SKLqrEX8Intk0HmI
sWPxIY0bnbEFrUUK3brDM1RfnJt4+FZVp66AZzwfdB26Mae8S2OT+UX4bIiyrEP4IWZeq9AkUOCC
xPudTeY3IDWda77zMuMAxv4SEHEGg8wRQC+JLJpLg7b61eOqQqA7+k0kRPL3CRgJ5M/xKOJaALRs
EE6jtk++RGXDOy72sPnpc/84RoxgYQ39dd7qZYNIsvLrxVmHNBxIDc1vXb2B0mRVvR39IFMBNRgT
f3ysFMydKdQOTK+gkcMPtMWrJ60rDPm74/q759w3OqrUzCMFDal22HmXFZ12xvLa6jaMekbiULdT
frUjrGp0wv417zlRjK5xWUrgr2MiIZzXZoL7ON+ATTS0K1yZK9Z0By61WY7rqaD9Ne9doRb4KIKj
1/2kUCzDEDi6y7NWiXG72GODbMUVCCxCu2NJIxuJNv4VEftG5goO6bIdk8nFp8HdI+5O4xtrUgjI
kWEiGAqxgFTuyVpREnqUyvCpR8AxgrYIdc6B5z0IXD5BfJLeHNOCHTrB9OAqneqHNFrHrf41AfYQ
yiBmZhe1M8F12mtjRWGyFDVzWQxVQAc7SZ7bnEw5cct0OCIp7QuEXCIEVE0nCAvye1QYibvByVQ9
G59PxXZ5BbylOW1zbKrjGxn+De7H9JklBhtdaQWJ+fFTkhXaZLm0D6uTmKOkMtSOsoby6cFLUtxl
GHaJc1Xv6rQBBGv9I24qx7u245S5rReVU5gCV/DaMP5erSWMa83CRefdCunXBWZAyjpxP9LeFvZb
X+OWM0WdPRLdYkBFwF7YgelFQxh1FbaYTdRgcjbiAxwCEkijzGNQ+cYDGwFl8byvZ66P9+JJrddl
U18GGrnoJC2Nsh7C+ceFWZAYXYbv3atca3wLH2uRc9CTUwf6za+IhF/JPA9RSkRXPax7gFkqHheb
K9Wee9kxGpZ9AXa0Re3UdMKwqlPbVNNJhwyHlT+3YEisL5z3eeiwApApIUlklDZXsYQWNICSJahI
vZ22YMMOnYLSko6mnTuoksvD1YIr2eB0A15fjepHolnbgnsDknVBSSwQhI/oG007QpX3FgyG9dEb
0PnkfzTOnzkjZ4hIcw/Ti1GOYCwzWnaWSWNZnHLw2gpE8i8NajUp5FdNQe1B2l/IUXK9FyZShKLU
ubqpSizcR26tci9dy6M2JUy/t1l0yMkwhmQ9ZVXNILiSOiNqGNJu0hh5XuXCEWuxhj25+RQPSYRG
Dui/1+fm+B3DZTaqkEyruT5Cj/1guzHkk9nZ0tHD/+U+Zn3X4IDh7o/wm2IwsRpxZCLMNX4QTlYm
f25H8upcT2CEjQ6RMicTpM2dGBElYXYz5yGsOHwUJoiXvDt4NdZweU1AbOLid1IFjsrKZp0RsmA+
+AMkQTgTo0OYHUP9IYbEZMnVufLXNvrdCqsMPnGExZA9+U8rgMFMSYfMrx0UZz6jEHevwuYUV6sV
d2Z0joCPcELbzevM2/+l+rrv/CjaA0KumhwATYnI8s5ClcUKAAHTMi3rFHTq5oaLpS5ePe2DDQXH
LjHspw6u0kl+x+UWqkwIBfrwj0EiMZQzVB3DCAFhnesYBRJ44+Fe7PzVRaGRDsUdG0odk6ymu1un
QW9zXxZFTgIBbmmJvtmCn7ZMeZWSWSQom9b7XPLC575qw7p8wEOWpgUk0ok2hU6m4HCyu4sOv1zS
CW9dENqyLWvjQa8MHmmJCKkT898+qDWn6VFu2VO+y7JT50yBduHMPjht1K6tkk+tJANpVTWNXMmn
hAkgO7zvUllWwUGlpmNEghOH+usfeFhWf16ZICZ5do24kESAYWW4zXSrrQE/m5tsvLVuLKy/p+Go
rxo9sRI9ATATt47t9vmyCH8J9ZVmccGo5KHqaMzMumzuILr/0pbnjdm7pLwqAEiUxKG8moEoe9aH
rFeN5X0RdrOYTegu/ZxQSsgMJP+w/zf53bhjKyUcPU4SVOuNGsOKDD4nAKBxqy7y/T2q3yvF7xAr
tu12ZqtRur5dPKOtPt3j1u1PYI1fgUcH6imgPb501DwnZCCNkEGrhs5nESTV6g2WmgsqD29splZi
8oAG5OVsoXqi99d8aR9WGvRp12Gm96zpSaK+rey6/lU5r4OcJj4+68DpdsAhb+7PSNwz11ESZ4R1
fr2nBx+5na1pX0DlxHEHdqCCFNnuREJ7xpDo38Hgwya7+b6kOWNryQO5ePgt9HMNZHP9HF5s09X3
gOruHAQuULQmzc2vUMzHK9kHO1QmdhH0yGCe5heOyKqZ+Zy0AiRWA7xQ+LaykCzE31OdiXvdMO5H
vl9pZPrNGNas9TOPJhZNvRjSwyryTKsSVu1TT76vrme4ag9d/esFS1Q9hYKh2aoUH2QgNuS2SeFk
a9GwQm0WrPvpF2KF3VQvgO1k3WXPckdDwhxtXHpvavHwHBCV1f3cWBP778+olZz5QVSIO65FlX8x
aRF2Rv5LsMyGCCXPTD2GYntKLEpaEQdavpv/MbVsgseKW7reTYGJv3CJS39tug5krnc8fC7zLcX0
4WDii7zGbK2Yasl3xszpSO67wqhYvd9JokEwm76rIGZpN5PN7B56hY3q/KqZUZgYjqreN2eQbJgc
+IGcyHzTEXr698Bjs9oXhzQqKmhxhBZ3iyJoE9WmzRROFeXQViAHDCy0AvS8v28/mee/6EdOGaCS
zhcPO0Kxc6UdFvyDcq6GTMUKWshf5dVh0mrCDFgAX4lInrshnW17aTFvRqIteM+JDnTA7EUcy/FG
yyQJHhRPY96dEOVBCePaJ+RgXnLdLCsdLkIo83uxMT2BWqwN8tbG5+5cDv3uQmQExnzYfzlN7imB
Sd7lULQwn2vMcY38gWA7HGI4/9IDkMlr/1MUREbZ4UyGpna+M13kUx3s53zU/Ti18fg+7zUi5/H1
OoZnRYIF17MjC7rh0hazwwe40Ajys9vwVvSazhTiJHX9EhWWb1D8QyfnSH6CwBwxVK6hPCJsQFv+
vZApsc+riTA2gYhBwg5vxvFt/5PIU9IfbutTcGbNIukFcbuNwtYYHlaIyoC8hYdLXKB6DsbTJpK2
PZP+6oXP2mDCIVr930fJrQ2xbiLZXuDfv5GucS12Rm4nOVZbm5+g+vRUOwhNXpfiWO89BdD1xFDC
6FnSbokQLAA+pT2y9iLRFOf6BtxWvU0F66HgAgYO2h+Ly8vgd3YJErQDLC/GRfuk67i6Ef1/+ukk
XT6Dn8JuEYLucWYplQIMfARCztrI9YYXM4MiZJSyQ8uKktUXOJxCVSA9UsfGcdBb67NivJpoTn5g
FAI0UCDHKcSYwk19rIKP163Vue4xjLBYd2XAfEeR9pf+LbAQDYzJX0NO18agAZVb3EkhkLGgLJ1l
33tcVLwJ5EijzBHPMZW4Wh8h+cSIe0ujc5Q3UJRBlgdZx4ko0Hg8ewHvZM1VGA4Of9nOnYYj7tL5
4c64c8ydTDwXEWo5JM31/iwdP2bfu5inj+JOPtoBpLkCQIZYGuuYp7AcpREpPkshmbS45FkVo7d2
0wDSPIw2axnoVtl0Osghe7V/V8mSEIktr9kCXHkP1rvLpSuS+EpBA6iozH4vodOxpsDvcMW5ScGB
s2z5qWYLn0JKDMe8GSD2WlyKXc01uZPEvRa/TqS5ipZ9Ukc+lAJY236WMspV1BY6JS8WvTal07lg
FJ4BK1sHYB7A4oa3QYGXGjungR7BA6UKWNGldbSlr5i3SXR45XNe8pnVVkd5UPa5JUfHBpw3f8aS
NhjUw2FaNpYZppKh6ikZnX0ndNpnjFdUAlXQ4f0xfOlrfLnetL8GZCm5uZRBaLWscZqFCfJN0qhS
7YwmfHohPP3bYRK42izcBawPTFe/XBIUtMkJvclAtp7xqEAfW24hvDwc6KOTvPRn8QUhicZjo6Cf
Jt04xS35ZkGMy3E+Ij/2CyXLm+5jUpj+GJDJfmMLc/kzaBxRdc/QUtncU9LY0B0P3Suy95Yx2qs5
43c4TalKbDDs4cC0CPAYEW/5suc2THChhVIbp9Aw0NEp8Navi/b64ZuTQhrnPEBozWCR5NcC+LHY
A9jkTW7+gYlInDkZQW6BhcNllN7zRuKRRf8H3Hoy+I1txWmwyCUbLRnMY4N5bZSpY7NCy9WGxC5h
aXtsraP2HqRHas0SIi37eBu1x1zthF6miIYzWv6If/EYYs9cYxp7Uwg8qkcs5y12oxLgp1XNPoIe
kZz0NmTs5TL6/F84e1+ibr0e9Nn3kHsjv5ssvts3S0zgDcKxSGbTyALsGGoHsRXif3RnuSRrYtMI
mO6N9sscHCDuJSXyH1KYaGdTDh3t0PT6C3jnmA1/TNiz3uYbvWQV4vbAUy6YYdSSRrxhN7kqQoCO
u7CM+TtvRr0E7lsxRG+cYaxetV3zSTl1HuATMynJtnFznGJEMEKYRUus5ltArMBe6bMeHZeXHLo6
uo4IpR16ODjvCbHiP0+xHXMoMOObVJy8H8uW7e6obPUxcJ0L8zFfegxv9Q9vI5CPyVXuU798Uni2
6zgTApL0icczqsd8d6t0FRucpx3d+5DIrMQUlOfbFDfOJc7xFqJRsza6Euw9qeq7n3amuxXQ120u
gy96VLICeXj5NBUBEJfI/Xc+rHvPoVsgHm7f1QtB8L3vfKQV7hx9bjt4eevNyyaGjWVGXBtyNtHv
O6EWOXZJozm2AQMMnTexYs5CspuB3mNEroMTe5YI5SuJee2EH/i9nN63tU4Go+Yr22VuHUeaARTH
EgpuzevHDn5DhD2+rLBNg3I7wZ8n1VrNAl0LMvYQsmfPv2xTYtpSCH05huL+djcE1qoBFC445IOg
J/XzsLW6dtbVxmIuTY+fIvUh+z6DDpW0dXDT83yWCAfezeJYgrQ45jIKwvLdm/ePArKp/6cMORUg
UB4MpwbGYtwuyebJ2qDu5CGKDUag8Ejy5G1ss/iL9bd+xQ+F02wkgytSWU73AxWDY2H4xWbFXXeZ
GZiSy52WtFc8Pu4rRIcIy1dNdo+uOl2GGhYQniiwaB7OEmWid6YOWxP3LcaHYvkj6twhEFDpYYU0
FqNVmiY7Xnt8htnWC9GWLt29Sa+WVW/2pkO/eATjBkz/d3qkP4r5WorQ63Qlv0yzMD81TVSE0tgt
GQ++OTXeyUJyfxovq9Rx0BFIcZ8X8B9PYFP2vund43bU2mqNqWCxuccjucCKSAQfQxa5uIskdCwA
SFHzrgE191Tnh+hRulkrKes2eaTLNA7FeTEZM8KWXBImPpnb54KxGQJpetNosrEzuWUa+SPd0KG/
lh2d/FDq7hKPu0Q4ktOJz0TGd6P9AkW1UBMkcjboLd/qihv580GE0Dz73clWPoWnZkjRoxRaGo2T
NE9cSNdWVD0YRsKL4t79uvRvzLh6rB8wrG6pHDandQ9ZbsfpfpqsiQzdRXn6/a/QkFmDje/j+Sr5
V9sdHyNAa32Zw2POHYEnNeVZTtId+wTESOF8e9NNatqQL7+kiFmz0R0zqxBbIacZGSqrM9+Cq9fU
V1xHhGbbdO0/uTiITJKyUspOUgfo+xX+N3xAtCQ+n5kYRCv4LVdrHOM95sYSAVywuu1cxoDjxJ1M
XPg8p4QVkfLOjpqDSxrUCQS2nDMDR/Kwpfi6e79hwmitcTnbt7vQsYaufSsU5CiiycXSrFHVv3lL
uMQmGndb2cmM8TBMuM/u2G47dvO+XXgGw2xdtsvFdNLnxmVtDNBAz1QPBdhPmbYxNb6hJq6uxu4+
2Za33fnmQHLUNpZImySj5zYAkqcBDWrU1UpIH/5Ilx2dz+rRB2i+UAyfs/LxrN0yunStmnZNNrUj
yXPnQeoTtEtmn2YkuX5VShADHIuZAKb4YdzV9hE/9XjeVs4xEo8Ix9XVoIAWvqJUnCjRP/2hQ9Do
aS8YyBFNdz/ueIqKonF2/m6Wr9vLIiaz+VgjFm/QFmILLnHB7wNt0aJ02G/yBujmfmIrcGWvloOR
Qq8NbRJd43p3wtjp+wznLCel+MKDf1avTRyyZzw2YgR7YcJtt4XvvVAiBd1+Abcl1ROsI/R/dMLh
Sd5Tckh42p7OmIpZrtzq/vfDiLEfbfgK3wqP9pJpoy6HbHdO5kjhR8lTqYpwSZ2xfLFHc9HjxaXd
dU+Q/PopXxgJAU7icWLz5j5QPQZfPAgkDu8yGKoT2JhmJbiKLEbW8VkJpHx8iChY3x5F4d64y6Ao
K1XnQpWr29TD8I6vd1j0Ir/ICl4TW/46CpNr0kuTsLbp5V5q4XxlgrfuHUVjg5bYU1TUD+DLIcHM
jv7ctOUXZDqFc2wbOkdUcxgFi6Jnfcr4sUST5u6cKeXlNpD5asV/jB709ia0/6NPXGq2j+ff5NGI
/NEU8I4iMKi8FfnX8wUkMVZapbpgZk+NGU2JQTkxmodrr3hlXYWEbuyWfxI8Iu6TyL/+3sj3yCp1
8ZbpMgTyL75KI3fIrKUzFTyG52LqrKPn+N8tCZlEmtoAxifEq4SvJvDaJI5FxXRLqyyn9Wb142IR
QvVr2jm9gKRPBD4dV8pzBNhINiI+sh/9ryN1ybnbf3kcbWv8J+Q3+5CZHIcYFOq/c6i22KsH37Ro
83qzVIeagsfYWVEwOirCqaOP0vNkAC0xpq1Eta8/Nax96ZuVdVGVCuLk3v3G6Fwf8zfjmh5jNovq
bZbY1bD7d2wA05mlXTEdbBAy9E5dZAIHYoWNRcUlijx7pgfoRjE3NKAy+l0e06JI/4oJKTqo5pRm
mIFSATWz6pafCBdkyTrN6wuSH7uv5MdaeFA3+UpZ1HbfyUAdM6w/TVM48XPfqAag/JnfOeug23yk
4RWwE31Op5Vsay9VLbUgp1XHhfUu2nSeQWng/IX9jpz5zpRtUeGLdpn3QZmX5xM5nQfV+abwScuX
qGNEQusM6zXvGzYoY5qiAMKoJTCQB7LR6q1IiZ9B8CdBtNA1WcFOhq/8L9ZeBeL9oCKTjWsq5QmB
nQyDOHEdvyyyZGVob/zFPNKGY4mIZddqTqjDpbYJv4/eZDs2cV7SCoGrzrV4FaO2cRgEMP2ELdTK
vTcg5afhS3JMaVmDs6QfPnwOaFaBCqGllpwZi/jbQcUdB3QQkBU2okBaApGJ9XAtq3b/LogjjP0t
nz6I8JnlDWc9THAHciEatLtVy+VlMigmJnKsyqH3wM2wzp0r83Dc9vxh0LoaxxeBSocAPLTKS0TP
kTHkSul+Ca8ijD9uGkzLO8Gpw1fbCvfQ3RRUwS2cFNzGtPLqEIdHnltmWsudONLipxpKj44fSTlc
LpJOc9abRgr1OCX6++ueGeWLEzF0KcdXl9hkCjZaLnApK0VKa8RlT2jJm3SPTmnAUBPTaaII1IQ+
wB4K8+eG5Q0Kol9iGWBaSzWKUX/UYcRMkr1q5RzYgA7pJcGHOIwaNQsxfQP5EDAHinyZD189VjS2
UIGiOnmNzUHydCp2ukoBTpHyfze/IgLUXXwYzH1Y4grM+ntcwlA5AWMs9MRsfS8BEbmWZ2OEYcgC
rZfHGkhpvJWqm6V0ScFP6aQcm+GSu4txX92DIFVUhLudCZhQYwXX4HvrMHhwC6TT8QTkR7+5NyO2
b+OHQ2VrCtFqN4RWXcy5U/mxueavQS0NVjjOUkbkaMetX3Dl96At1G87wB4h7aWvYCSKSY5q40mX
lcJ/c+QF8YiZeXRkeLkfLtzYTms9NRBM026iobnXa75ltr9FrHlAAB4eugnVQ92ox1HEDoFzXTxO
eki+re8dyNynH2G5PJp662UhlWjNnRYBRZyJHAeVutd8gT6kIZMPDKoKfY2Kj0nbnWTvdIk+YRqq
SEZqrAdisw67SuqZQ1KqetdaGVTRomx2mUQVLfWI2ybGT4x0zniA2HS7NBQA+y3Le5pW+EnN3eFk
WJVB3EbSCvY4pOUZ8N+zJce08Bppi7Zk7WKMfsPnN37n6uMq1IaYaRnmtiSgzU5hzR1MQWb/VK3+
keNXDOrVPoAjvwSzOQPBmtyxMiEXfdEOgOT1doXpwzakuGCkoD18NzuKb/7Mi7arJXOF37gYDXNO
9y+gZjlAZugS15oHhEKAqoCNHNhs9JvP8ylCGjTnYqbGOc8B+/u1ClZUXjVR6t3rplqOc65Z8VxQ
tWKgeNfIR+sgQ5UOolBS/OjcWIufS1od4JeivzfSuVkSWI6znV2lHggaWe7BldeLKlcIuWKbOEoQ
dwTrMkG1yX9Py/kzCOrsHH2gG1tIUkl/aHh5qPPZFwgTn6+sIKWsHksKtY+u9QeCggY4iWDx9azN
O92IkqM9wC5VdcQyYF/62rEQVtCT7n+zq9K4VyER1PWR2QH7Xitk9D3H51OLm4VPMDum080sDVDR
QuaS4rfOIVayM9iN5BlrXbtHTTKsGuOVYDYJQfreoajwySzqWMcijRzI8AWvnTQJ/N/77XiLSL14
snmCPcngIb1Wd4hWPtb1czTDx4L6/RS7JPnASnUDDhLn2JCMnbY5HA8vbca4sebnkmZu5ohf9Asi
FiisRn/UoZswfqF86rohHSxQVVUIwzzDJYd+0RWYyhBkhcWze4ZM8DScmCJg5BSAxPq5vpOoQFd+
jWhaeF9jCoiOcMNJCHlEJDwE4IZnbw5mzZKutlPFWdbAOgUtZ2RoApOfP8714T56S086rbJYoZDi
4kK204ssuSm7xk7XxWgRiidDILd7rG65vT0nQMfEwnAcMs0NBSQdKH8Mb1tHTnmuB66D+U95ztGC
v5nmwMSIvAAnAs8/HUIFzV1f5MYBAqMijy99PhLK/ADxzS58SEyHuPZJK60kq8qjfC+I5TUjDmla
gBHGz2wUnYPO+elJ5n6Ux6RV4VxPw/T4PllsoRw8urriJ2ebwdiFTJNKz+BayQ3lHhZdAsWfaKST
ir/uT9ONoGqXmCfI4brajYPcxhzPq5baNYAp68hUeeDv4LZhL1SHDWLUafsAXeUy1LeuhbRP3DlE
ejJOA/wRn5rcIhQQi6Ca+PCPtJtt+2t3tbJ6dDCz+1h0lKSJrHW5nT4M6gwCWjCgSx3czvhdELio
TJLyGphnbxQI9iCPv8ymEXDRXwe8GStghdBTTHpX17nSI5H3wiizGvSgf5nYoiEuBLsVl2g8nIHN
6Ap3NpewG2Zz9tAEcm2xGCWYkz7bUw3t98Ce0FIOvVCOiKIEOZZ9KDEELWZUcmTE6I+mPUvy0FBM
rMInMeTYA6TrzcQfiBIIShguf/JgooBzcJ82lK+/Qkzp0TvOytkn7aj3MAT4cU4DedyTLX86wNYu
FFrq1E+ea5fR3X0EfS76cGGIPkza+YNFKyspaJrCTwGIy0oPOY6C5IX1xXyPmhdkeNLhHPqfEoOn
l0AetlGurrt29MBF78gGvcLpik3XbaF+3x1cPhsadfZgRXDL/k07ksyEAtdz+TjUIRHryBUUNdPh
zsEHe2ufshCi87UCRa13pZvGS6pS9tYylRUQ1qdkJEpWcvliO2M9RXJyJrd0m0tUAAnWBMimEwGr
NsrZcmP0+dzVvNOk7wNCMreHarb5Q3jeiozORjGvDsVHwIE/ZbrQo3DYkFgcAIy0+rsDk5UpALQt
SyTz0d38QAKiC/hu4p85/OutkHYwhXoerj7x0s8BCzYLLyP+LIy/0FSLTHRrnBHtDgu7evrw/7/E
YygR6Pie3gLl3Zfzuw0VRfGZO/Bywq71baCA0F043Ed7Mivr9/370FZlEjU2xDoxKVrc9SRp3aUJ
fTyCmItcdPrXVifYClT6ni2LaPhS0x9zBPwxQxgWuBLYMu2lPf96JjeqE4gglANRpsye+/ierNvY
UOU4zuXRmec/89nWE6nq3WxfeJetylubCvNQwfDhYqSg0A3obB5rPZce22ISDtlFcGZEV6qa96IG
aLRY8G3zw8Qriknnt4FZLEbmHBQ5tYvhBTLNpkf1w947MdSCaSs+sHDTHtQNhpi4kB6BFGg4nrWS
vPKe2U3Ffraxpclb+VWuLUo5X/Gs8SRc8/eZtwhqOupPHGVcGoGcaLjgevWvv5LzRooW+pXMpOpO
GqLjkDfu9FWn0698IV3KzdrYkiNxHsYy0x0G3GJ9r1DakEIscOeq+1uuxGknJ2ObuQT5x1KEtkkV
JBgIlbd6mM5k8IZ+PfkRnKsGCMhAMFZ0OaQEwUoNV9qVK6i72yGR5hH/Mwrdo155kkSqJlCrbCEd
5bpEA9wGNoN7Jjd39sa3e4vl5rmeQP82ym6gJ3NbCbZqA2FVySltwQfZjs1GbRsZwep8uriIHhse
OpclfX2uF6UCG4prVJeNAU4hUdVWwqvrOwHJmjMqpuI+1t5G2ZnujD/ig4EQrcFo4szjzYVLHaQu
iDDJMf0dg9DUpDt9duVSZ2iW1dkUASKoWNIrrQQU0e9PYmH1tqwWUd2RScy4J/Myzru2tF+93k96
38NZu4CbA62ItpAdDl4QkBrvGkdF9Y3QK7/fNxdWEfujHxb1fdylOnt1AXn1PpuaaNRgJj/hRU4U
q7d4WSFms8n8oFys4BCW3AGPM3CQZ+jMvdOmJuPaZjy5hvIvyZxRVHwDura1Jp4amOM+QCzwstNu
/BAN4R2bmeR/lq7rfuAhoYdGtXydTwL2EH+jvJoF5q/0tgVkTE1yxA7X1KBGsGNpnz5fwKY0F4jp
4tml3Zhwb/pbIs9TXxPxtPsLj3BvhQzlBgTsrNu8FhBcctKxffaPejP57pw1Zf6nTl1JgWXMHakN
WqCl8VYs/iwmygfoLZebZCvkwaiJunvBvu2gTJGsbqieRTI/T6VoccyiK624ORaT9HHiHjsIYWDj
Bp+XNwy6UIWWxjEx1/OMo9L+eyx+NpY6ddsRL+d9bhLVOpGH0HpaR1BUD1+iXgVDDNK5szFkkBVK
SBRW2+4wzk+Wm2V9BvLYaNVHWxAJyTqW1RtoeBHaqpqqWCTb+rB37jp7U8rDaAZgEzt+Jd5QMeUy
XJh8vmToBe4jVJclPMjpKBZHNnhav+RyBL1Sy82xCmElvLjjwcfkAScu3KHOrSk5GTb7ShNcRIi8
BJSWOtDgMgv7ehweB2rAUzryE3PON+BHS3y+/r+49QH/IxdwvV1kaZSwvA5//yjGXuAKvpOzEb8H
dghyVJZy8TzWRLyINfn++1A8+k2EtS1PnWOct9GUZEfi168Ah/1phSo8cIsZ/48RC6lgItbBKSak
PjEJ7iIgBCsRDc4g+R5Arz/0rgtPg02/ZTdmct6aGM+1TiFfpMh441CpyNqzlC9mb6oN6/knhjPp
aarhbrJKm9fff/dEm4DtPCyBu/ZOFsyem/Q6UnmRkGjqfr6g70goqpxcgWwx+LB+Kyt5dloKG69w
629YqmOddplLC0w+GkrGoDef4unjssG+13rwio9i5moAt/okDiAxutW7/q50ZeMg/B0O8H96H3h+
JmGM521dSp0Owng/PL0LDSh3k/UfFOVkvv/21bhK5rtGYn2xMYs2a7GACfzMHRI72+B9amccGFu1
X25lHm+REQwLjexVpVH6dk5/fVj0LYoeFbF3/HB8+zKfbAyKGVsUuq9LVDi3WinruUdZmgmdd/3a
OfympJmVp+vS4HiCQjR6+PLc/8+s4q6BTRODgs/MZF2oKw2TqHiIw5N9h0mUtl1HaRy24DEr3BP0
JfNTfAEdexwjyB+FVLOV+0kRSE++78tdMWsh8bMAml2z6+L+SRn61gw04aJSZi9yEGmHwv44jPq+
TGHYVX/l2cihfimugc7SSlgwyr4V+l6vN42JChCaiLRdDP9fizAlPLc4ERrrZkI0aoSpkb+T5bJB
OWMrtNeRJ9nBbE8kEdY5uxc2+o+9NfAGYbbp985oD6WutO81DeRI7H9WnsZlHXQSaadXyVClpULI
mNp3DBv5EJlbk+SKC2vF1PbatzMohdSi+s3wpgWzLirkE/+adv8RcMjlQKTimNJFLrlMKgslAly3
uTiDJpTAlOkINIw7TbL3xIF6g0+fPlnMd3PUQKKYg7Qj3bl8FUkn366t4z3QFtupIUoOXzJxziTK
2m8deOu6QPCkV53rXoCI9EyavVLtBYlH9x7cnmJLhSdvEpPSKmoJOC8KYfnXYB9QGkerV+zXMGIl
O/Hg47rgaOJqDuB0FnSiJCkiSXui9YLXNDxRTUg7b52JvBYr0FOfj/JVqzkZmFn10yFZD1WIAzEz
S3Ch5wDt+JLz+oDUWLxodA0Zka8mwipo0wyUpwGrSNgmpjq0lCsxGw8Ef1YHcVC1Z/IFMRRIxNpU
b9hUpY7R2YUqVPC9jtUV2R/tjmdTGGdCU31XpEyj+ZHyGqUJouObs2Um3UdbPFvqmcYytksqr1f3
AM6ByHBpO2j0FC/+ZMQmoS+T9f1A10GTsLJ6sfl/uJLhIrEanRQFhaGxNf/iJYs9pziyYa26StIG
UfTub1g8Q9Xm159GqKqYRmLVXdc6AsreJt2RdWdK92YZxnUeJ1+L9cD/0BK6a1bhDEDK3Z/r9d+b
r1m6zspu37+nTabYq3Y6pgrMgDMnt5bue0qqdNviS7vHtou9T+5sP3y7kvAmYf2je+p2L/Vy/gEH
W4nXorn3AiUGv4R+E3qsUzFDVJ4ID8q14nyjv4KMT5UYfWVo8lT+J7kekHv4E0VKzh913yNqULlI
DngsXqaJ9SCeRCYmkcKT2MIQhkVTIv6YUTCjtVkxL2RpX1fTtm/+xShmxDWVTZMi/HPjs9e6l2SD
kJj5zIJlNzw3Cddlp4ctKvyZKzyweQf+c4gbOwDNtYHGIGavGWDeBbghXelxnqsKP/N9+vqgY34i
ra3A99RFf4A6zLqSgMdNAn8Uhy2ewRY/d7hIE0JuxeeKPHWS2Lh6mV3spKA375JwXOJpGjIuIv/P
Or9SFKq1uLXNS/UARybEfMkeo+GM3cywE7LdPVVjUjK+Wv15hLr1BvCFjfH0GWbny/VRwVZzKKwV
Pvmvcj3/BpQzb0OippO7Axge/AdCrg//FS24Tnanvx6muoQ9Ly19UlTZ3kt8ubeQ+kDZbpGfljve
k3G4/ad3sYZ2hwsQ7orboaM/Bmv82HEA5wLAyKZ4ayk9KZudy2rG1GvOJlAKHGZgMwLsLYqEW9n6
ZXvUx7MfJu1dnHP8EJYWkL4WvQ+Wizr6K+UFXYkiIFwXQcyL5gUqQop1WSR1p5yFoCjeTXZfdC64
R/NmBqbsg9xV1tEhnHkj4mlQe7kxvSzO/jUaYu9CYcxZgwRI8ERZdO/fisZ6DRJ7xuhHdVWf43cp
HsAFDU9xSFYK6LHW+Gm/je2w23SJxPSZnKnc0nHrYejxHzNxjk90dAuHBnmNICkYzv6pvdImG9+I
BHgWivroRtCeefNCyvE9XJjmYSzKiNoFa4Xlg/nBGXG4nrCBxegzWSBpjXfKOxd7tjY2JBiYwKgc
3Clz0uWsdt74/ZtmVdT0hShQBDjZeOzVz52/33cm0dOhsO14eBoGaT9zEWjtuiMaSoslYJKKJwPg
dtlUUZYAoDqOscXssaR0ced2ENPS7zs4LxCiBvYVsUApoC9sp3n1k9B3CX5IMr8Bq6GJGHvweM/l
anqtFvttKuGIhzV25DHKRdvccPjrmwOp/Nk0vhvOhq80AoH4L7d3jgoFJePLrfxcpb94NLIW7Ow3
ECWMXKLfa0QhfqYh3NykU1KHBGvm5awNBYHDBTK+MbpiMAoXlBPzeold5Xpi8SOKPsj37sejzD8Y
gSoVrkRoCLdIJamKyE62u+7sULy0pwGp3Zm2+4zKn4D2aTtIepzavIqnpXLpmRCTY6IWnM+cUE0n
CQR56p7vagv8vsR1zePr0k3liUQhllja5+VmGwNCo6rYnKUMg/VFZQnmGa5+sSUx2DQ7BusMjASQ
fw7vd/KxJLCtN0PF0yf7kZ56uDekThzDywvhWgOh8YczkHmAUrrKBf9of7p4XxIO+gmA/hfLiyxr
YjyuPJsI04keZ27elmUSNqrwG41sqpGW7U8jtZkrCrLDbUeVB2n+oQWrEXcuQk6jhpsXbghO7wZ7
iyDY5eCJn9mXEf7TpAjg+crvyUrH7izd+C7lqT2sF3D64PT023CmZy6C5r+ip1uDHKCybba5FOCh
CWqy+lgUmySRGAzVfdT2SMiYA/M7iGRPhkXV1I3U4e9e05R3ULagPl3yIG9yylsWuXe1KLPuXFBl
7eOiPGLzGK+o4CDftp4lZqeFuV5r6ZkLSjVyAvgRca2psIqkTrA4Qjmvju3OOuZv/fL8DCdt9oFm
YaUFDtRrzz2SNQHmsAoEJCaPbE8Ae7dY2I8ZiNg0eJW9fQIxA/g33TP78p71GJOTh1JAqhwnScU3
YIjo+2ntvZMIB+F4P5N8P7wWTBtNUCWBZDuKDoKr/2lUdZGhbuls7+to4XYQZIJ1CV+ueC1vIpOx
R6aP6egr+tN9JBmNxadKoMsPwN1+P534k+ECDcQsvyyzTmWto8braROh7QNZaj5uEoZ7iJnK3W6u
/foZy99kf8qeNl41nexWco5W33rqiTvOrTpUrSFGBjt7K60QgEsnr6j8AxFwLJHwo6FjlUWsT+2k
95j8H3rAyBkD1N33fsgr6TNtYfgfWF8Ng0JX9HcRNMGZLaDkEP0lx8t3bZcQwsQx7OIapwk7fn/y
H7OgCjXIE8CenZPPjr8ZqOiQTqdhAFxsTIPzeDkWeXujxesKd/WEI7Rb40OohvbuTg2vlbhm3K4M
NdVdbqTS3Rf5uBMeKBQ6/uAIrDyoAJWuLh2z1k45ycxxCDoyRpZ/xP/ZMmWhip5+jQiAJ6MU1tPy
JyOHlH2BqxmtXcv7U3UfIEyyfwZ8+nFRu91HS3YAK00g3O9mvSROHfmeSV6nfXCxWF31H3h4FmWG
H2jNFdpP6QEehXDS581QgtxtFaKejtTSoDHugPVjY5Xekn5tdKXHdHTEDzHJgrmEwZLCd3b+pEPO
oja600OpMkXtCs7rIe7GJ896KAhFqpdzpo3fVDMc/rseKuMXaAsbCaoSWooLn4izQpG6/y1HV8lN
YItPBQe3e/uvu7EBQQeKHqFupnmznScTKQaXgKQ6g7LlAh/9opruQ2fAAlK5KC5A2dOyKcoaQGJE
R5MjfCTJZJ1DQo5hQh1sblM+7PHv86V0FFzZ3s/r+wvaSWOGdfEUAbIKoFcU0oyljyffHEVZBA1I
KaZXlxloDJ79OuwZjQV0QpPtEWYgoU36M2km8mI83rl/fs8yalaaZYCZtrdQe/Ey/egEohv2VVtd
zFgim8y8+7wzpp1ly78L3pbiJsiIVWUFIoA2Dy5Go2eQoOReTVNGLQo/TO4Yi2bi6uBTsdACS07p
pPZcB8nGszldebr4xaIKfffHJhmWJAa4yIFXaTzkwY8a50wtCeLi1ZXGQb72ZM/QRuGP0ru/AuFF
W04swuG8n2TsgJADRIvOmmGzsfilbK9fQq5dkDhdwCHpoKf6vKIbQ/3JXhSme37oeyZ9ijgh8M0v
nK83VxaxEyF/h133oqpmJZdac9jhrmz1Y+kdWfi5ksftwglPh2U5MLvA4d/i0ngTMXq/o/KPlfFj
10vTw3jSEXziC1TKv1id41I0FUXJszR691W1Ga68uXT0kwIE0JkzziKh7PLW2IXAVWNO0MexN95p
kGvoUL9RtLur2vZgUIziAhYOPlw+wrDaLOjyOB4I5bCXCXcVh61yCUgH79tMfPHvWhxauNzT8Exp
JqW77yTTlCcxmeHmz8AbyQVZPbPVWKNsmz5FAVCaKL6vrbeYW2DplC8j+mZ7fUStFK4sRpmbG1c+
0xj2meSmtqa8UpsyMlJt0AK5NHAAoV5V8KRB043HQqhJJqFgEBOuXLwVZvNhT0NMt5CBzJ7ONIDD
QbbYSAXTGvWg1vopkcPlkhRPzybUYzPyOy3dZo0Hgdl3i90ZMmZOmaLAWJjMOtht9vIRqLlukYPe
7HMmCpgI0/IxCtVNenH7FSHgI1jchPI5Sti201n3A7GpSp5XD6aANjSfJtNtUktKO7d9d27n8D0R
El72nYHSOq05nJT5cttwodUzBoo+IBR4dbIW9HIVYjGB+CRTNp9na6v3kHYDIdNjfZ6ZugS5zvr9
BYQu9iOPKr9gYL13/7ItFTYqLJ2affZLU6aRPJGApb/Y0XaLKhbpLeCOKb684rfh/YXjnGI9cUWH
12Fzc2innq3kNfUrYnPLcFQAriq1KrZYL99QWApXAaPQlj3Gls1ATyj9vn4faXYUhrqaJ2K6YjPG
8jqwjHLup/nG5Y1CoZAlSn1LgHcFagnKakMHT+i5swW+or2be0zcFKb3dQ+aP5ksnV4aIHDhaqcT
Qf8vK/4jMuPBn/gHTLxbbyo91RQtnWFD1MYbKQd+JscFjkZudE1NIefOytw9s6w6BpOcfRlhxTQF
B/GUZ/2EzEVOAXfABtPv2sNVRl+/D/SpITOFVrpfv5KNJRHEn9xgCRHxdQv39BaLxcrkbzM+RdFp
m3YERawlHbSgT0UjV6mM6S/TWp0QH2lrBmjGzSv4me89pfzVDkqiugcUKjGVO3WiAmjW0YIEq353
lhqpLn9Ii6yKoYdZ5DV8lE8YiHwbBjx2FevLD0t6v/Mtma9oUA66PZwOTrGTzREHkGRi2fxL/j0S
gR7qfiLUYZ4CQkH/X2nRR9x2aP9AkGOqEePnnAd5kam6eVmIx4TemrbY02Pmcnw4Uxz4k4twhTlE
8GwFPO95UMm0/YtKI3FNv4x19hFzuZOeEz5cy3J3axnjo1KZSxPdudlU9CHTdW57ZmQ7CiwMrtDZ
F4SJLv5HWt+7lG7JmVhUQSeqgjSKQmFdLbKyoj3iSWLJIyRvrSMqaGMgTeHjNitW+z1yg0KAsyjr
2RPIYUlEzNldAD7pXVztCyzZZBmDBQdlLMcrhglIF96/3QnBP+LC0oUyF+h4ZkjnEO1fvVpOScUI
fYiX3JcFgYq4KVjcWZ5WgaZuQp7x7dHR0v1NlKbBE7URaYWWIGzAFpX+FrUjFnLDXl9KRPhAINdj
1fXuiF7RLjY8/L/pH/uj6en54IoqadBH5Ez4EbfB3gNZn8JWayHXrqYsWBwmfZZg7iW4JTD31NTm
LEHbEXbglhcnY5eO6YcQGioudutJxo/Z/cHqJzrRh+LFO6JQRiwkOHZaOyYmpgNkB5jCrb2uyrQ/
dxS2IO8yyalpR+Psud1l/E2B4uYp+JE7+huJchAury8KCtyOYcnthUqBcOKaMg8WA3mFmUgUQpWB
PCgQTYthU1fP8trQiPdOcYhA7v6ZtT0G4nJQCoSD9apyJJI7as3WRbB1Kt9NQWwgySd3CsbdX+J6
gkzSQ2/Z9vRZon+nVS7wtiGZn3Z4f28quj9YyhHiT6gMdvXU4/7JMc+blaD9ugCwdODGB9/elOdX
WIt9DmUvGDbjyxDX7tASP+0cWyN0NIpWeNmM+S42Uhg/5HsO2Hbv5p+0oO9oR0UuRk5+G/aL4Shq
r5idSvl1R4lGZLZvLjNSO+GH4RjPUl2+bbA8qti+Wywlhg3k1UcqQ/V7bLjxrVKzkP616LpNaYp3
K1OmKWROLiaqGDRtUQ6LfZMDU0lvBLgneObWwVfTRY+ZjbSydD/Lb7tfvCnUEV/sNsV5JOvcMZff
DJ9zo1fKM6Mxf+HsYgld7ARe/OZhJvKTUT+uaQWrCQAjyi+kdW/+TWR8ioHcEqLJ+paaIXgz4/xb
lUCaqdSOcAhfDYv5ASPaLqxb0hZDFZcK3MkvpnuRf61oEdouqOi1XOHVZJCc+czpi5x+N4lh9Q2a
bye+KPnS7PshGqqfWhvOFpzfCjKVm665LrDBH7lIV7n5kak+AD9JejritSuQXr6Ei0zvEf5L3+L6
Ym2qSD+QEfTONSc7J1uMZk+5ZZxRqL+RyedNOlVrq9u0yhkga/w1L/QOXXfTHSycrAJqsjpA8Lk1
Wd99frDOG0Xpui3D6WM/jetAgQtJdorj61Sg0qxjQwEY7MbxGAQEL+NMPoYgjhRYOEKLAx5f8lQX
ACZJb+HXYnzFZDoMnT9q4MnChyQnaXmuWmhSovBVYp9pvDcT71HSxWnh++424lgS4mdAlvCJtdkV
JA4fpq6isDcqI0TbLZWKFwdnYtfUfkz+UbzJ+ho4rb3LHz42wYtR6kC7Mnf1tYuGrATRI/ydzmc8
k6SaANAZPGkVGkDPd26fyYRfU/gyjKD18qfCG0ENb+uBapgBtZCHzBqRHADg7d1SM8rEthUbycXq
n2Gnwy9aQon4tZJOFdpSdIovf4P0NitQ3OMFBvYXkULwpCDwMkZEGP7jVb74azUBEuWSiVG71UZb
U7xmwLvvwE+6KykuCkUIAai/rh/4r/wUEJZOyYVPOAZOgiY2a+aLc3qhfPLxRVAlsxTeIxEBm9pb
/xbwCCHCNSlI503mkRhPmfYWJDQ6mptyLu+cC0zZhM803dcGlRcmFVvy9wcxRoVyvlKULAl3HNJR
KVTAFeDtZI2R51X2/yYhcjAwJTa8ZBQz0s2X8nfWsHd4WJ2JCYh3qUBZfGUiphrTw+AGc3T1JMfP
jBsZccSC7WWfFAyGTf4t++P0kjTi7h/lETXpg9r2W5UvrzInbmXRjZ+R4Zs89BiwAm6yE/rJDOYk
/+rQG9AjFCxYaiUBEbXzwYd1+aF84LbGk89m/EEW77DFLgTIusM0XgefJcowGeUAwkYM5yjB88Yu
d9hNlEM5nllgZ/K4ixEagfc3ne7i1Ii1mVtupUGhtYEthOopAg0pSnToA+ONqHDgVd/YnNVaVBs6
KJiy68yQshQUNkEQ1RuDWBjr+HLYqkoO1UZgMlk+7p3Yrq3gyIFIzCMZ2i2JUmeulfMHwG6Zeos5
cfqHQbJOwrBb6LZBFglYjCdxZWZA3MoOCF5gU2N5lR7n6+3LxZEeVdoHwkxzyv7NvZtLk4hobRf6
TJpvSmB2IK216EJztH7DJ2rJjenpb0AAyn1EMUrpucly3roipREFtYwnSjm1e6sqpXG3axyivW+p
He9oPUFJe9y18vMtwxct5D9iyTctEB5HqRkKP/IOeEvUbsfe7/pVWlSLFkUz7UjfWpL0qqKM0dpo
GRQoAJwQfaMnKO7o6Rp8AL6KJqFUCe8ZypwczjyPwkLZkCpU92elk/wq6j5AMRTQxb6Ew6XdqGgP
d2gbMJeed4yI91kM6hyVeVdh1lqyzcJFo2cs7A6y9bilrktio0kbeor78b8twUqzllJ3OVemaUX6
vTht7kqLfR4P4LSiXAs0ClGdQ9mFe7EqS5mLn7USB/ohYWMPBp6x5FaJ4jkIf+2tzpqWPRsLIOAZ
8mIxNAW+HlSIDkLfjUXXZyvayxODVuhkn2z8h2QLV70QRNNLKnXSxJI4E+02vR3yaZ1QqLwQAGEh
L+R2vsbNupBed2mddxXLChHp1w8CCygkk6866S197LXJXPknigbL2a5mDAE/uOy0qHjRR8od4YE7
PQXTRNr8FqhkPje57oofZ5XgojlaHBkkUjPIxupO1ClIh8swrxXqEqMdi2ky53L4ywITKw5T32JE
jAME94VYKU+A0OJegVFyEVn//jkR+NKOpelYh6jLUPmfsA35EU8JOOW+jjEuyjdwrsC5MVlGBomE
OIMy03RnlfeaQK7jeGZ3/AAZUFmYunJPOROtotyWSaehLGx8XpJUeEOteS8YBrampJa1PkXDFy6i
bHUbFx6Dc/PG/6MebFYK1dfzZMsjUPrjec67a0+wpkrLE/pLwwjb4JT58QMLBd0ZaN07XIOTqabJ
oLYnt7J3SEwWoK8CzU45L/OkR4hrZexhUEI66f9cdpng2pNUpoJXRwpVwDXo5PlTuT5se6DkM+j3
mBp3410U/mLNhFt6+YZ2m6En0bgEFKbe5A/kn/El+j1RBb7hoFqf7VTuwxBnL96wkDQHhZhw/MKA
er+UOIAMDIj60wZK4OsD60EApYP/3OnpVV57f5KUryshvvy24PLbow6jNoyTm/TqUfMcXD5JTFBr
bhLpaT8Qan7URl4W3lkusUo6FcXn+vAJacUgPPQk1/dVn5GETsmDPc7bKVj1kADXgCSw92mzrdM7
dONgL5XK1asMetGvXjlv4rag0lB8DBzFoxAJh4hCdbA07jGzo6Aq8n731HtiNt447NgQzgZI6nGZ
kTpqslyJ3Is/y6hTRBrEY/P0OHS4885fn9hBAv/+5/h3xWLAObsisoiVvY1+vJd7bGSY+2Fa0fre
ho39OgkArPh8zPvRN+98foChlOZN9rWIiQJUGTRShgV3EhW44R8qhXyQwIYKiHm0gYF5DWM+/adf
KXw3E14OyiB3XLMMfqKtg5B+Z81vfQjwyxBUxotfrcNJYnMsh9vqWaMOx0BPp56G8dw0COUUMArZ
klRHYl6hOhyqx37pZb0sXVvNzyt1/mjEC7B/CL+fvdZp6KrYQPYpwRjOoB5s6gJZvdgzKO/GGKPl
5KkOnInre6BiJQVCh4PvgiNks2I6SLjIJtdLm+X+hFW7MI32SK7SKSNIdamHcWmN1Xc74SmXH7zu
aHsmZW4Foj6op1j00rdcshxijGK9Ueiw02DoYFsFCMa0Nuz9MPgJ2cPDWsaoV2VcyxS0gqqmGJHy
Xe+GYyXRrDEomSnmzVfVNqpi3QqsOjMiz9Pg30K5mFJt26TODgRrAHrWrXTQ35k0Ug/7kuQY1s2W
wR1e6JX0f0k6MU9OdsU34cwKiqEFQzWx6sVG8XmLYrSpjeJscGZ4nmSMKnCRs1Mfvwd5iCazBldY
XDCX62chixXs2a9gDouaBo57BZxtM37jOUWZDD6yLk4Rts+bgcBI8ye8YB6ft3g8+WUgiqOK1Y2x
kY4yTj5NI/udus5dPWqb3cusxOyPasvK8/EFlsE2A+sIWZRXPoFdYRMpZ+8ifwoW2bcklSiomdBQ
c9SiAtX2N7/sMoczR9I4LEtUCLd5HiXJALi8qZWui195mCirCtXQwDkzQVMif48clKH6JbGVgPs8
HSDB9tNUmAyhIKlYYM4qXnuOOIuXRtFRnYAo0HkPMMmBXzJ3teIX/DvexWJESrzkRqIeo3hnwDDN
OvpsUO/4ZyxmMUy0sfD3Yd7CcfO5FCQb9xr7ryxqScnAZQfGG7YG7VKeK0OBbEwcs/40INnqciTX
FKWKXiDWZpkB8VX38Mtt2w0U60uX4j7AZhwiyFJsMOHBSchvrLay51Waw3U4X2yjREF16Ap8awGG
ROMGsnYPkUXwocmbvd7WCwrhUQVQaxD56X8KT0UQpwEYjhctQiBbZUanUD7DtqniDw2EcZJvYmAJ
LE01a5hIQLauL6eZGyojrYfZbgyOMZevC62xkldu99NpT0B31D5wQaAkJCTMbZKYUgxI2lHpM/s3
mQtGnSRyBrxY8Nk14SYRcXHt7BKUdvkqrD9zVE6K9gX/B0GYCoh/bjDblZqnPGq7nnmiuTqIwmkr
dGvX2p6Llln2MkOxFRdBlfOlCZmUYBOZeg+y5qZw87RD65NE3exXmFveNRxzI1KD8gKMPtxkA/Eq
USsaGQaZcepPvXfpur+hHqLNd66gmAtrsV+xqOv/8XJ1LYDE8ePxiHQTnbA+0qROevg9t8cCihi8
D2N9AFYiY1lxREUWzod1wwrJG2ZwuYu0PZynNkhZkeRh8EG84CBPs6+8csc/OBm0ZklSmIKmyEdu
bqK7ntoqeUXWl8A5lN6kxeMQa5ySAdxHouHCFhlGK0sbVLqwPppM9c1AwXAFx3hGJFmmYy8e+CL2
vtPEFFvbwUaWgCwy30cD2z+1YFLr33bQP0PHg4c2oSfC9fZOVickQYRYlRDgct5nnUMu1HybGU5u
Zvz2WIKCAkXJAMbwLOYH6WlGJg6KyLBI7UyTgkMF3GmG8jy/nKZkLf4S4W8gcvstN6HTf4z7Gi2J
IOeAL0rLR4DOvH5mLYaeQuGP6u4FYFddVJ/25btJ03SZAa1tMsbNKV8reN0DQJTV8YggmXeYQllo
OW2AsaL2Q18nXcXvu2ZifCSZxnj7WC05QAAgA91nPXWY6WxL8gXzEDWGSv8JA2GOrGC3/TcoVUCR
/ozwfx6FCsDFA7G+kjNgS/rs/y3G7VO8yNDePFlpiLweh9A5EO5Zc97T8+TDIsjzXCfoVZkZHxGl
VQvpRaLOcCilVwg/ljpGwZ5XqRm5VKIk2GCA7teQ3X9Uh+S840w83LY9blXZ9mUmavMrgwXpPzM6
laezzhDD8rj83Wxmi6HR3x/Uv500go5t7EJc+TeZ1ttW066+WyZ8gKrO01GH0SRNLPEsmO7j7Gbx
jTKOlmtVk7U7ucAzzaZj0QFX92WurULn+KNIRBP73OEyBMJbWuiU7GT//u6+RTeZtT57gqxEgR0D
hUHA37yzvD+bSbuwTEUYNa0wYjuIWr1U01CuaSUeNH9PoPRJVZhBQnzZ4U5TlVp/co+hczh16cPi
vqa5jsrp4oZjusYcTREwWhScih8azC4LqouF08QAV/MZNCdTh9n0fyo1OoTppWZ0+KQvd7ZIN+3n
eSdzjJ3CLXCpOQIv2z+gbPY3T5CsNPRtaA7WRBFSmiZMF5/38GvU/dM+XHtCGJ7XawLABp3f9+8A
vt4y/saaYjkbsBCaSnLhkrhJ0elKEHR3wi9X3lvUksvb1lYC/fupu0uEwtVVGf/Az218RyJQeIJP
98Z/Zj0S52rlQ61YiofJ7QgWIH6HXlxTmr9SYLK+AUuT9529wSbq/exqsMZac2wc5qbpbb2z/+5D
1gancUKohjzmYTHZ743hHVjB7lSBW3bAYJWEQNUN/tH2z9r2BnutZh6U80jFxSntEkNlEiSFA6VR
bPogJpU4LAXwJfeqJT9WY/o6QmsChLnn8arZ6HPzhJFSKBHd2OKO7s7zZyOWmQDEa9JbjLIOtJgw
Ietc7t1s6K2lP3wSqLAys/xytTfSsubB1a8IobfcLBMKGa4i+18aIeFivShsY+PNxibN0Dv8RaC1
fqoHbGpGcv2jFgKbMlf85iwjTbcpyJOgF08RvkC7tMnwPKMBiKzrWCxSXnQHdcNRcUWr0g3aGdOg
9UYQ6nX76eIfJWxO22D0oTGOoGjClyWLM19hN/8U3XtLRs2uVHHUtgRTrnKdLpB9jx8iKc18jT+5
K8bsgq00cuHKSA33rRpI/XMS6XF131/d9T8HZIRMZJdC/93Gb2lqmVCqUGrOLT8lh5iSj5rwO8M7
NVvS6TSlYACNZ7x+WbJgII++6vWNpprvAoyULp8PnnI5oIvwCsbOSXDL9x9zw1MTAAPheYKLzuVt
w5Gq5tDJB/rILF+4kVDdWy3njlsjTdLDIwCgDDK0XeHZ/DCnFW2fIYb3z/+5VbxsFo+mH36PbUUQ
HuINBK26lMoplkbe1h+W0X6AEblXaXdXc45j0CWuI3g+w2+hY9WOEPcnNkssxKgeTavmxRxx8jmu
fAkGJ8oc8PW/KBCN1ExbwHaXuLmVCk0MwMfMgLLW39l9HXw2w+IQM/JjfUM67hWLqHmissVCKB2a
t5azJXrjZ49cVctoBSmVfYkLTIcn8y2bAq5Wd5HPxa5OuFzohOYcQ80hH1au6YZC8unvqibKl+NN
XqNU/Hu5oE1K+rp+wnafDoa+u5sEsPlOmnnDyc7GZHdNiJDd4Wk80sjpWRmlTWHfgP3mhxvqRcRP
AzXLG48wwHTKtz1uVykklRuZXH1bGhJFA+j0HGQw3q4P3S62xXoyPHn2Enhx4/cddHk2ERgg/52z
KlymxQCBtiqrkM9wHtu4HljvuiczHZPWh25eUEJYvt5LANg3YEAXZq5a3rldXVG2Zsqnyrcd6W4G
D+3hDzL9NxyhlrNtVINQ5D7OXxa2ohTmD0gCiPNgIrjYc4F9Ky3lRNiXsJAuWJZSPkSlkpndLLIF
q6rgj8fE8tkfn6qqTYduElgDtwKnx0fsEqBwYEn5zhSby9N88YG2QT7ilVvlXCJxwUhGab/EwH+N
9LgKnRQIu1TTpQg9eQZpR0jt/ohg7DJtYEkTpPKOih3BGuXZ3wTUIPGWFwpmdGE6KkNvwEe3Jh9F
tR7Oq916xEJAxRwTHA0iaPJtxcyewIhcPPnslbG8ovZ4PxS1V024ttN8ATB7npXK+pP5vMG7szuU
7dvriQWKalx/IssBPAX3NJZCSp5fAU8qMkPCovoa9k6OPHl02i1u/gBYGbNucAxjqrSFcaXvjgLi
i2ymfqC2Srx/IIVQGG/4EHMm9V8OkZlqzScjzUIHquBAY1yznRuJwj1Vm/y3Ijoie0hgZnSCiAiz
Ku2TaQxmuad0l0yBE42sjOrZvmVBq3VCCxKRK5wZZ3qJf8Li9xv09+XZ+tkwQbODcN4g2s8As+Wf
iO+wx/DdakQHvBQB2SZm7bg2WzGdOzN8boiXFaTORELayGy/BgvboyTyeVJcx80bEtip+Sftbdn9
gflQha7+UxZPAeFmEqCNQNmfMeVvdiunPw/RZY8TiCVIWj2zApu5LJzOyVxOmoVJnyzCbJXZCy9C
mSGyiOBYSr/cykunjd/GJ4C25GDFFY3XYva3vyUwFOrLLP4hkp2XwCIq3Q4Sj0awNEcg+JNNgrhi
5vGd8ws8mMpiI8c9xUljDzp7AOJk0aCGcSwtPmu4HIl+EF2easMzseGYFy6CUSWl4mXmNvE1gk0J
p+bHvc/Vzw8+yabbn+7gW0Ke9xRT6VanxCnTzvbdR+N8QPWtYSP442dAGYo2IuKlfkVMD41Xd4AU
HQ5JvmX8LKWWFI81x7UNn1BsS/r0o96Ain5tssSNGOGFXh/NLKBfbFIPP/bQbVw+RA1V/VqrqIeL
skC+I5TrsyKedVhMxHCVT8lutZ/LqmnLsWoSqhalDYYZmXCqmYBj4v3dDxryqocFYsAEMv9QSSMs
lH2OP3quZd1vuIlk06HKMvN8+BWoMgmFh6qsH/7h7wXYcP7MRKsRwFyeC5FxN0k8cACA1S0iL1oN
c7ww+gyAcCh6pM1VpGrt305wBmSK2Wk8OYFwa37qGqXu92IACYV8UiZwgPOpmO5VbSnWjJd9mR4j
nyMYfaWMhrJGrY81ppqBSlHnnEML1Um+5JqlhLv2lS0YxilPTW5cJNaHdSlczW4cX+mTLhMLCxNX
+wZUUI8ko2GA5iWXs8whsgS8/Wwb448/AAfkgxJz4aVWT5G0Yebh7oAuK5eyoVI6Lyj4mfcSSJ4x
700rUOmfXHJp53wM7LYTVslXK+zSNEjhebKEeuxcfXyTGTGcIpmjmGufpbi5cd3t6IGetWk4uQ4U
VBd/0ATjCZWnancA7q5xbITkeLb4XqxJnug4SbNuW5CpW8Mxz2jw/1c1WmxDTj3EGrxV64VKC+gs
ZRAw52U8PyVtQiB1xIGpEImIBdie0JVXzNG8lJY2G09xBL7EvGrVR+h8OIJzktKSKWa7tfLKarqz
aI+hsUv4qBxk0yh5Hp0lPObzMRJ0h02YUDUURwK5j536vzEr+6mlALVKKBbL73SdWjzf8bOZcCKL
yFTnMdCUS3Fz8rL6LGiW3j+A3bx2ZhnIKFMcDU8tYKEsJ3/sYRwN6iWNP7EIayvb6yKTy6q7r4/4
aF9gKP7HmnTxepzJXOXeqdVnLqA6cgnIeqdyDrFRJqEo6W7L4s+zBZXGm/oGJU7WNQu9qZOuRlNb
AsUURNYsYN/O5rhJC1hyewc/avO3VeVcP9Cy0YGiQa+X9xL0pcIs22JieQXMFEwDaKi0kPwsPmX1
LrkPfF06nPA3RmlDWAt8zjaFg9Wb83LS/oYf1eSlKrdpwSnAvQVdRcrdKgHl4WUptm3wcD6YD/9y
go6LzBErehTP2kKlGEWED6KhHCUwNXUpXG4iPR3VUlumJV9yntk636xWOxW54atpRZ5oEpgF3r72
KlyQcaic3ryiLIhWtReK/w59PhxAYQjr8TcgZgnnMWcg1yfPrydEwt56T/jvN+P5+iOYv0+mFQ1N
bqH78zYdiue2WqoUV/vdn3gqVMSlg8guHPaUbdLJFW51SigfDwIhK2cuRRHZgAMw23G0AF86lR+k
Dp+HhMctvik4pBGMaSfqNd8qB86qCnvJVaN80U2mekRjhKj7LR5jHtyQ0vtePLmugczn7hc/77o8
i4EZ2Z+ViVxZnRDciBRSC9nrQ7rISSHvlYeLBMfmb6cRWw6ZT06Ej3sciyBlRz1IFdnh5YgwIAYS
oAY3ekpfbRSaLxcq2kyptmyny4abirYDlRnCFBu6Gd3NqUUVS1SMKR0SqIlQ4izWIBQ1e7W731Mv
URWDtiKAt5bTciZZS6vqaFWDLNXodwNIfMB5dsyBxp86/Fd41a18TAEyirJXegbklTQ0qxN5X4ZF
ySdRbQ1SKXYjTjGdqa7H/jaxv3wY0MAosTKjqcKQCldean0IwG73dWMP9BvCHwRMtyXBSYvufm+4
Dx0meXqkDW+oZjuIqLJoW4kB+aJK7iFFS7qY57oYQB0AY8N/IkuVkS1ZlzgRBB9xtDbPHkL4SSVS
NrmlAP/1sTVaheFgG6BxrfcJpCZ3EzPETLxnjg4zPNYfDOqGFXIMaK/Y44qQ/nLNT0HngyIIA4ja
vURkizBB+3LzmP3D1AXync7/1GBXYb65ORwhWHl0GDXM888JJtUAiBXkQL4K/olvckIk6Zx0l4Bn
39Gw4zkbzBIR9Tur7tB3K/pAfnLNWykkZVXX8aM9qj2m6GBCddhLGRhPfQEqxkBLnLb37LGUy5C6
nWdUaW4lfPIvWUa+ffMDmzziuxVnc6zIpSqNparGywBBgoxnUK+rVT4YI4nIC27J80JtbolID6s7
9vkAt5T3Ra4uGY3ztzRraUM/Ej6NcC3ijoewKST9RUMY/f+hVftlecUKYAcVypiUyURw+Ek+OU2h
9GPXIxfi0HCwA78w0mZxMhHbWqeiekFxjc3IQdg0i4d+FVOkS3TEnEusvOtNlafpk81Zh1ux3J8+
pA7TDTG08zauBo1oNd1BjePgVZCkAyfh4X3GYTVsq9iykQgOqY2Ff40RFqxqyxr4+dMWsW5bneN8
Na5ZVHv10Z8KaL1LnrQbFdQqy33vOyJbMUk64j31x8OUHqY6T0nZyMpk9aHRekHYJ3uFchFkwNkR
hGGJwijKb2HEVFyzdGTgkhfCbEEI/IJfjMBwCB4X1TOBvfPhHn7vxdwI7oPYuVK1uTFllGqi5DDV
2O/x162byHKW8be/qrsHw9QrQVGjznNz7AMFOXa/eHFWbEmS+7GzjoH7BhfLis6ru8f39qZ/tgFF
+5pBcNflN0GvtE+JEBK61offAsUqSSSFE/Ye/+HwsAKJbni5IGyPVk/Llru7qfihgKj6f+oSOx3V
WgvSyPrheW7gb83rZPtQBmkotmZOiWwiG1zbWoDGcJfFguVM1TE60NyNUU5qWEtbe57aL9Y72HVe
Ub+JDvEfgTFYWccYd+9PPEReGIdc1K/3Ph8ezxI03sFH8NWE/eePeC862iNcEAGdTrthnz+sRByF
YDHBs18/VJXJOuEi1Q+Tb1Qqlt5VgiCh50caRQ0ru55gWsSYlpDhEPzaWMa7Y4PZmfER0dQcWiTx
2Lwjn0eHhwUUBcnTru/UEOPtfqDIqq2PyRqhUmSBktmSAGYqqeh8mG/c7Uza9YzCA1KqBiAoRgqB
2fIOcNNo9nCpqMwjwqh/f/vAIiP/i+sTwZXZFvwaC+mGPF/gQ/+sDILGueHESQpJ/Gd6uhB6uIQt
UuLjAo8jO2T9rBeA2kBS1JoRy0Xa6UXqyGWH8X3BtX+ySweaio1r4of3ikNRtDpU7rlLW+q8GKac
2mD9FC8GrTPUyuJAgUIUk6QBxViRE2XlPT64szrsP6Vx1mfnQJOZ30nc548px8Z04jjD1BcxOaCJ
BuI6C9OQFkzEUGE7M2tI7BizJJNgaONFWe+Dyh4+FzkJnPXl4mUfPT08qEnvtBA+AyO4MVky6YM5
8weYnnm/ZHzjZk/LpfHHlkSc/7hTygxgH3hoEfs/XcS6dveI2davVbGXQUWCPksyc0g40H1jGnhH
9+Cr3CoAk6xFwJY/NxK1d9FY+h1z+LxUb5AS31qDWCxE0IGyYJjoKFYRl60S+GuR4AuSYdTDuBXf
zeGxzP26Cv1OU9t404hjtFGJ+FGDwkhSd6Lea1dE8fnbIDZ1BLcdaZOdanWdzCRMbD/giIvpJRFE
r8UQSDgS+Xv6ZCOl6zEnYuzPMXUbjIiG70uAEI2Uyexidb8UIwvIHRzFlG6yrHiqYNwGk/cXibXx
VkdoRZQlOhy75uvhNusVh89exRtUQGAD9S/lU/d8hHgMHuNs4ndVVC0JRROYXx/hV0kUCUcm/vF/
qOd3aZVbuMB718/v/t6LAtC19Z70wV+LIQz2+crGaIpGj5MExlAapBcKKQxNVBKvbOc+2jFbcQWY
yvsUD+VIfAx5LqVABafrmOyPYwEL7cfQGcfBCsJaU1T7wCFER+YxwPXRr4sjWaFNSr3AHPuElgxf
ctenD68Q86r0XqtxJsklXM3foq4sK4y7VmHxgToukb6NymINKr8V8lazEmL1TjBGRYLm6IWjKm4l
8M2ziWaKIVwJe4Icjn4NqKDmSBXj4dpNbO6g0yvdHg+XtEnqBz/YobLB3fYwaSRYNDxORDH8Z6vP
WOXv6fvA3slJ3TM1Um8OVlonG61uxrWUMzxyMdmpk0VYRQ+kchtuc1n8d9iSv2133c32cDEB5uea
/rDkDDouu0Mq4triI/NIOfGupKZaUirhLYTPpXksOmMT/R91nvLMOpFXGqG9upcRYATn4geFsd1f
2b5FR+VWJoHqZH2JHGFOu5B25s9WYAAYyVPQN+Y++3TuS7WJUNB1NsUCbSVC8kBSrwcCeOwck+qa
pNlNPiKfj7x6m7Rvl7FSoOMFOrwkpUm9QGrwKEJPbjuwCAwQXp8sCxKG1iEtIltvlgbQ4eJcSpwX
bQpnoC/1ES7LYGpeuWcAPrUwSSYAactDmhQ6iGt4m0rV8dGVnSO7PtII4iFXKVOyps1boamIMgXH
vDKeOefd9Utog3mWA+nmGXrPnL8pCnlFpHu1JajOIR098buoBjLYIRIerQGY/pdKMTbeMm2VKlIr
WFKjarNyiTAZCwD4BPvGicqTASDl/vAG3ATHHMiUR7wHq4ZGlkFABRGeHVGC0xpgy3h24OqESmHs
ZS6j+fkhNCyMIp0R1Fmyv4DLktnRdoPd7gjZvWsDFxJpEMenZDYXk/Y2aIPDGy/mhWSPOPezc+gR
7XiP3GyXXN47jc9OncKvCBa37IyS5g20T7LWA+8yaJyWRIJCkzquDxSJ1gyYawNfRukCkBpebEzj
IS4vgOCIP+U9ekd15EDWosvtbbjkNEeQbKOtngbHvwB2N6XevLkS1kxx76nleLI8yjjn+MEMvo5J
R7Yk8ra5/DWcL2mReQs0A04azRFFSShK4NQkMRreqVZ1LqfxB8MP/Xm3E2PIPlAeITjGyaehiaGy
1z0nDeebQg3M2OrWj63HMUjY+rxnKPKmohHQWeTZoGiUtR7mZ3u+oFgeh5B2UPu8D7PNfBTDJfko
o5RVbYQzomAgZ8BHsFCV1M1WBHrFIPe1TcOSeaWgslw9eQKwkpuEfOzU9lprYfQ+gQ46uNSoiv9N
Wj2nIS/9J+s4iyz81MAv+F/tRyvBktN6z8xj0bWHxXdRTO7B6lqMa1saVS42UY1o0uO3j08XvVpn
wMJEBIr0OzOQKsDpW76EVmOEeN0qtqqQSRIK4X7dfK8Gwu6XYa9AK8rIztbAryAJb7sR8KfTVkMz
M/Gb/7MjxCjqEtq5KkbGVY9mHRDx2wV56xZrmbyQ69iu8vKNHxzcGv8e+gdprRrCUMqVwuSF2MLJ
X8CdMQjSO2qS0wQp2mlbFxTlTlXBPXijifmNlcIFNYnYNn121JXM1d/KIoucCOHq+jwvzv7Q4oOt
ZMfNA770s2XTe9/x+AiX8v9R6cfb0h4BLuZnMnZMDM20E9t7tTseU/dye8CxcGRHvT2/8NshmQNy
Ez9wUhbqq9/2cQFHVVDYHK6WecgahMEza8wgUZUYn4EPbZgo4XRrPGbWfhrnhc1M6NrlIpJ/8fI6
Rpxw/TTBROKHCqzed2Qbs3r+x+LnTHaBH4bBW3uNoH/0Yz6V63VzYuiL+87g8d/pV7yBakSrLA7S
hyhHmVE747FSCnDcPS8NfWFAIz4srv+SEUkErh65f4lns0wUn3gZJNiAK6kTEgzjWCsWwA98odmd
MQkasaraaS2OEvXqemJ2mJR8zl6Aw+jTM5+BUOG7UEgGAECzbiwBwyg5qf+rXidkAZzgShx0Q6EP
vbuDlcyyn5ppqDy2kAWPasBRthvYbILu+LV14X7moTBrKXuiufKGoNQuJ4+8lT1l+SLMU2Ay7Bi1
iv89Lmv9nHk/b3kq00v3IoJMm+UBFiCVJBtEf3an4xAsz9XV216whmbCYYMwE4W344+SSuqKXNy/
O0cAKvCQ4mygbZ6tNZmIJedXGHYvKKIwyeuC3RdUyNN/ZFHR+Hy6DmbqtlcGuANUp0HaBdNXEyl2
XdwPrLD0Vu3HBExRYVl2yxAIyOFrqRtdF/oVoFeHLHMziuw5Rs3RJZk8hCKYsevIoxtG4sCJ3Frs
5cc5IFb0cdA8fUQahkajfo0EA+x/pG1SlBkpSAu4qX/UfppQIR/2fNEIL7rVDItHvdGbdBvlq3AT
t9+rdefKoUhpoyzDwK2tsWaGSzr4fkXxFilFHHJjBIuBpZzISDfGnQvOQe3fMjihnn3JBcqLRrDE
U9ntUHWulePe9r6P+UJ2z48JEP2DOz9+QJF7ghWCGcjII51CN5or4souJVhvUkGv62h9BlUMIsdr
o0fDPyBXKHcNMVxrz0ROs4d6d5I+h449ezfyVeHWtAHg29m/eZoi0+A6U0AhLGupxF5Gs3/zXBEi
H7GVvERmjfQ3Eg6XMhln8U/r5a+vtTiFY9bDsJRX+ihDlx9/g2Ftpb8VkpyFA/as1D+x8sJFnWpp
JDCHMSUacWxYpvmIbiFUkNhgMmkxqfLFTkRkDEFUNc4pT2VlUCUcoZIXYyR0mN24v2wkKDU2+Nur
rAnsyY/cPb3hmYmPOHqS+T8KWLXvkFzONtzTmAfZPqBT0FfJExcEvVS5BJyu44U1xdat1HHaje/k
QG3QJk/7/9UhoI+WKEsd/tn5cAgEyOy09LACW+8UgwZzKm5VaXCxJGMm9FiXkX9OV5C6Qqyda7mN
+ceHNkUn0897BYTHLxk92oC16jHzckzGn82I0wTK8JTdk7qRMY6R7nJOu1A+KLRGDE42dIPLd0Jm
Ltp4TnERp1TWYXWne3lNMi0uB0fkHJSf6py7J2Cvf0x7jEmhTTF9vH+/9ey7E6xhEx1DNEpsFeVz
V7uDHjkiGKnwcEan5gQ1wUFGjtbyB+pRGoguhwh86hC6hj2+oDyKmZS8WIVmT9UYiH75bc9svxzR
2bLIK5V0mSfBjsWuRr4qZAYfWdVP7GQ+Wc3HD7m/K2KRUQg3YzypDQPHcYB/mY76nRvHJcCIVCkm
F84fWV3kI5h3ktsJqxdfVM6EJokq6/dLvhPN+SokH2lRJoPodfw0IxE0YLicjBY8ERkthrB9PIze
9TgBr7mPGQd2mTHEIg8iq0P4Y+WYxj7rQ+8VnYpyHi6WLN0OpuwGan6ieM7GhRR9x3PjqD3nv7xn
rm3VE+GyVfwJSvQBCiK4putTxLKMO13eVCf4FexVRMJmLwKPE10a74+GB2NO7ltaE95LrGr5NfVd
kXgucSF1v1ysaXNY2MpA5hiS45OGbgdKUht5AjjkpJfPvf/zrPAX5Yufq4neJ23Q02FInu1rF5lK
YXHw2Jva5fgtXGW7PpFFGa/jo4t6vQS81qOhmJm7tVwOMrF7Kjv3cQp2U7UqOUgekETrrPj3U1X5
HR7zJ1HjeB50G6sEiEFaf1k5GBOM8phPRhYmX6e9bqddqXX8GtmU4+XoybuUbVdlh8cDa8L/7ijq
uwTM0+fFvLiput5A9fdWa8B2mbJy6sQfQXPQJFZLS4K6DvuzkVFbiX1zEgLHV+mptQkhIhj0NvmF
q+erPWsGJGWXzDQp+I/eMp6slI1GBAkXMJOe7iqEFEQEJlrclj1CRzsDrxtoeum0vwbbBuKN7hQc
416Nt2mCPUHY14vMOdMohFLqNADql4G6WX+zo2Qvgz1agvpDGjsi4+jMmwhyrSdUiYYfvXu4PvlX
rWbteLHyZLEQusapavAvKKQOSird6unSVBovOCleo/LTTVrjreB8mXDAefRVdw6QzkmHJ0778Uvq
GoHYyHRgfrxSAml5xkJdYUuHEjzRJvMY7agiwgFI3hiGvpx07IQRE9S4HjorOCILmdOLrz6QFtPC
qpupXoOesqGwI3Sca4ce5hmcV0YbPLBYxt8lKQcOl9GR/FQZJuFIEiNwYSqJEgTBQYjiVfw4Dhg+
7PqQgsiYOZ90TfyH3ZonID4CzDYSDsPww5g6QuuNikZNhrpDRcxwXXKdqCRRHOYrvv3JBjNIqp9t
/gJWZU+QyJV2eF7czub5dvPqS3xdmJYxx8FMssrKa3Hp6lU6j49u5WO7GADJQspJEN8E1OXkAi9f
d3R/dkG9liGbTmP+fOwS8VDJfIk4ZA42jmz26vjZPZBTfOZIiWNKBFCmCNGTsF2aXx6HpJm86lz0
H5/NCBbZ5c0u1zvdodHdG/otAvdUj6A3riJ2p2nQfKXbbVDvFm2Mz0A+ANw696Z+Xkmw4hBInTlp
li87qXVStz1NGn60VAn1QlUaMMdcZUTyLpcZ5fQNdVvD8mdnoyKSkBdnijhmO8d8Hp896BKAvQdI
9tiiiYySavEEHOO+eWbm1OyZVjFHgmS4bOrmzdq4xAxB6hCITO9V0DM6a3JUyNL2yhdio0csQ18I
IYxOl+lnK6OSnxGwZkgPsy0i/0R/9antPmu4FwSnJnihNJ622aDN6DPXQmkZLjVhQ6gqqh7V4W7u
zK1wBMou1hLoK1DImqhOknFMQIxi62D93VLw05GSStSH1XxEHoqirvPjNqsTuitnbuItpGUi71b7
USSxJdasIaFj7d5TSEPE3ReACL4leENkzfwjSD7M/BXekJ5ZNzDNsmb47E/3foMqZrWj8Kzl7074
ck25Y5sVqmN/U+AHiltoSwCu7EPxVIayxSkfnJKU+TLdfjEZktEoPSCJQ7zUMPprVGZYKGN62Ilm
hczxcZbyvdvyt0nLFM78BA5IzwIwbuJcW2JIShPYh559/bZ4vn6Nvo7+BJhHSbbG88al4DAv6o+F
j7kIAoGWgS+MdC40w+2tsST0qZQkxBzqZBnaWLhErcWkdxm5HhxIzGLfMzcUk7GKGFVHHVBbPNck
TowLpZFPcGy2dbbns+azN8joju145EDeqVa2T3WntklW90L3R2B25tbY7siwUoMJIpWOdnTC0Tzf
PBxADI7pDodCcVlO5mGGg++RF7yd8vvEQMsDSmS8aYoL3/7E5y1q1VdhQ30nSavT9R724gSou1/S
iG4Q7A35xxmfxUipcQujxvhqrn2JMQVyGBHvcO1ynNDyL3OunBjlGU4wYK82x/MrrFAWVu7Ie4hh
d9hY0cODh4FTk5oPee2iyyIN6XBMkwI/o8+ljiXmOvwOIYjMdJa4OtZx9lH/3nTSFBcaisS6Ou2n
XcIFV2Svo1hOIgAGjrl5iZEjJk8E3G86XbTBSSWNNaAFwUNhFiMXH1i63Car/0PHXbU7JC+BLRNe
+ptlrBoL3TqlScC9ceZ+F0DPBBSRAWeSv2S20Nfo3MfiE9sw47btu3+zAUaCEN4Fh5ixaqVIdihQ
heeeniYW9ZxvehB0ijzWrkk3rZTQoGJHyVNdCPrh8Fafbw0RnB6R1PZJV8Vz+fFfHcZ+QP9dD4HK
4FUWv6ucyJEFNommYz9BMQsegKGYh6w5m5nxbXTSYlv1Vd09dPQVtrhsk/I/cBNJbEoWVSTsX/zX
5wccvu+uZyGomTe1ZIY2JAh7C4lMqqF1z8S1ZwSQeALMc48D82fdu393ajaj75rhO0/V3bVBJhVe
hxF0WC2tDIj+elIdOCEUxGUI2S+qTN9z+9CovFJC1eqHPICu4s2t8fow6NR7w/VRpPGtbWvQp0KX
7AG/FdczFGKo2SMgLwMr7bJKa4SfPd26MPvmL7bPph1KNZoCwfKGX1FFQhbGmak9VUtr2Vs2juvv
MJxMNbXRV6lRUOW4WeySyF4KslKaKKON2Zfv8b8es7IP1leNjJGUUVq5dtov6zZP1V/+mvocMRe6
Uw/XvVHh1XRGbSby7V8YYeaIUw7c7G7+EL9nGn3JtTLn491UCpv3gG4Zho2BpAyzN6J/5VCcXN07
fyw2QC29bt7tkqnZivRtMdqbkYzyiP+aEAQt2jStHh5UvqprytKz9obqDYSlfH7X7X+d276gcxoe
1CYi+qK8UDS68g4Ntfe5UzEHwvF6SGUEcExv+erx5Auwowe+izAnoyCMzpF7BtYbsxfeJIEdPOIH
Ls+F+h0bqdqKhhIthr74l7/F6Z0N294RTEN9AhCzLuyf1jnhQNZdFMoyVXm9kojw6qSh/3W8qzpx
0yA88sXjj7ucszWMeIhNEQHTGYAojZ+ojEWZ8QcblFUcOBtLzOT30og2iIj47RuYfBZYe+YrH6X9
cWzzO/tBf+2y4oiKT8/tu2FhjKoA2OcsOormmoe1ors7Mefof3GmPSBMyX91VX9vk5kt0MhXxm4P
L8s5oLRUUluN3phxRuDND1LTk3cfz6OIkxlXMF0B2rXqZmPWxWx+e6rChTVW85ANWGKD3asooZFH
nneOAGkzqSzCjyNts3f7aJ1jjCNWt2XOR43EgAaWHf+ZuB+1otrYqO+kBeDROsjXzbozgDMYlB+d
c5+9ocXZLoANJkqhfcVrIXT0fIsYeblLwe1Fjr5ef24GSKIISm7XoQ5iO47a34LR67mwbL/Choqo
CBL8ZuHpNUHpkfRca8U4nqJ8KcddeXDK6bVXQyQGrgRTRbFChAXiyHdUqFWHMFF9TLjkRHNXez+r
S2nnlZyGl3mChkYbbd2K6IT5rEvcwXwUDud0tKPl0xoc5VJE7PwqEoVWKpnfzE0dsNaz0xnqiqtJ
33LhyZyu1A/EQTDw0pLM8R1iHJmN7Ec1FWEXx+p/V24boyX1JQD+dm000HT0lg3ngA/wJFJD4KlV
IKYKJmKGpEIf5haepVOXshPOzBG3jgorX4x1ZtD57fjfQPFKJFMYKbvfPy9Bo99c7GQbZONi+Jlu
vE5KBDVeX6SDt4AgcDoe1g7qZS2m4AP48xZwIukdm7blbjem3fOgrVax8JcPxFW3sSml9s6UjPZt
pSiL1gwQUG53q0zKGRGZ7zgdPLYD99MkXHId61VAYbnkwX68PwMTw2hq1de2qqhAXKoaGh4L7JFN
E9wHLsiMP0vZtu0FlCbk305HZHS6sSh0jqv5434M0H2GMi+MVde6iRsUAn7as9gEpR5deqRzCQe6
xc/ccdTiok0M2qTcVFutwnjtHhf7DHr7VJOURVLHb1ZRJ+jvb+SBeKUJFGIPTM64MsYmYxRLewSA
rukI7ml/sJbMTVvdZ+BKGNoWgoRLtgUgqIjvSQAysXKJEgTKODf2anZXg04OMECMpmLqZCF6KgCK
WMRPVWgDiMu1CGtNUPPcbQNSWf34/yZsk86EygKbdjkGiyszOY9CSBzV3xM367QD8b6+RasEtfPQ
ghZ+qYCAhl1SxmVb+hzCH1P1QY4YZGUKswXxgvQWRJ1K6tUCxbqovJJst3KFQhY/GsOlXD1xJeRu
pTbUt4ZScQ2+nZuwZUZLKAstCToPFS+ueI4q3NnWE00pd1ATEG/dTLIg3xzOR0r7uJpJPy/B/nid
tXYRwa2w3Jk59zrzd3JNjySuuVgrFY6tyMhbZt6Zv9cBn/1FmYFalzYQ141WyeXrFmWeUSjKbP+W
DYoafWS1V8NLuy+pRQCkVur6nMQGM6Dstijc/WRlyrN+MQP9xJ26vKcw1oOwrwdEA0LvMc9itHyI
gLnSqbOeDjbKOL+az2M8Br5CXJcttTTF/DT8RA7+t1MGfpj4VTyjv3io7ttv6IZgEcmeRaG1ULfi
clmHgRgc6uWsTgLSl7YVNtyT52jstL4POPyNE1O2KIPbWQ+9+laT5f7cBfbRt9s1ZI4vmPZvaZov
5738igIeqxVDZM38ZW73A9FZH/UaLiRXnp1diiyJzwHIJZJWv3MHcYJyCwpg4FeiavOszCI8GDfU
9gD8a7qRpUrEzK1YqPko6Uk/C4kMDQ3c2sDeOwK8v3mGkJSjwGlGr3jnda6HX5tpmx5hd2sgovEk
LfUEId6SSmBJ6l1ebxXaohUYsD0OmM/U/MbXUnFjim0/LnRlKLcg34TmKZVstJusnePfQ35Aa8nE
QV2qfoYYgxjRbB12c+BmjjNpOy1efqeI99JdfWBcd2QXeU8jUrVfbKquuUOCQbYOobd0nEx3VAX/
JmJWRXu3Cvy/LJkp6R72uLdXPBLedsSvtBzQqSak9J3F0mN6G0zUQJR65BiqK5/A7GruiIxOeso2
xXzw58HROSlDxuNLo2j0PUoUZstjqJ2tAZw5cCVC/saxK/rY/duzCfCPszlB/nRYXfYObsBlaEnm
3EyRi4Bnx3jHNvA9vmfbYGBAyltXCTgCkNyvbic+0/thzy10HqgXVB3U2M1NBb6cbNpDanMtfHFo
2DRRm53VDwoEh1po9KYUGlnu8R4FwL9amsSbHfoKRRSM6R8oybcdV4J8KSXHKGOohS2gON/JGDVU
zWCjhTycZkx15/Wb1lHtqHa85CIatuBGvRcqjK/o/CvD6a0yNhsDgLE5q1JGzjvmhAyCBPvcWJVx
O04+wdP4KEAPVRZcXFtrQ3PNa79nicYA2uVg25rR8xNB3m30xpBoJgI880ruD9VWW04a7qD6zJug
jSMyIDK36s8jsM7C5XzVqHzoEMFTb4190TaA52WC+Xh4+syMLV9wuDhvVkxFXBRc1cfp+uC8rBx2
qWsrJGoUPhyZ/58R5z7eq9zZctyPBjrkjbAc1d+DsmQPaoiMRAMHCmxlG2tLuEUjAQnbdK0skAbA
k4rOzS9bM3Oba2DoexjQoxaXa3F+mbvXKkDnrCj1MqoQrI48kA1k9J04rNtf/2DeNsVZr5guXUL6
sSPEYC8THRo40b9sxeueCdKfFjthm08wAN5N1TGMzsrQr/+MjpAmq6q6IphIhRc+lWBjFkrDmk7z
h2jZ5uD8RAH/o20A+Z9o5Qe4V9cmtE1dy/G+8soreNz3ThkhGtJWwFSF+nHbilQUm0xIQ12V7deE
TEXk/LnQZjt8k5IEArE1Ondk4hDECC9u1eJJe90vdYO99cGpIb28iNWagu3TOfDLfI5etSArSybp
oC2vcfcWqumV5atvynS76oguo1EnV9Dliy+9g3C9TcJau2cOMh5W5tZX5dG5q3ePLKGxKOH3wXFk
amtCXCpYjfK0XFCbW9GhDhpTRxaIYY3oeajZBp8Er+r1Y55c3duGFOJ3IcdxWttzlTlcZXgpQEC3
XO8BZz+zKVTNdeoTIhLLE4uAoX3NxERV31orhotu+yAZ6MPjc0d2iY2Z/9ijXw3BGeitvfucSkCR
OoD2Gyy+cFvZlUgAnUHAGGqv5Ms32YjsFZDxEbKnAchPSteXZI6C1hJpr8IWk+wMe9sp8+NTvS9m
ItDo9rD4I/tkdJWT+pLF04adL4Iz5T400Dy81oWrffOJswXUHNlUHEQMtQtPh3dc4AuG7YeJlPKg
X4RBH3gM/gwjs174+V2Qp1spnl7TF/hXB9R3tEV2/J71o94Huj3nPoxm3vMQBlQf2hIUh6xqLpig
A9OTHrqa44i3ZQvM1knSChSIDvGyoOJZ/rpXpawhLJCSeM4WspLJ9IzAOV3SYn5fXOujwl0FWhkX
T5ED1UBa4ITkE066ExkyjZkISbZOeYDrYbJbmq4RbbN5O2n9hvxzfhxdLbAfkhvSx3ln75XC5CY3
K6pU2EbzIwaMm56lJZRaOfuCFmUXZUJTNPFq0Js0iB9TZpTr8ldWZx8wQw05tPFk5ysnm7lkr/1p
+CQV5i6a1hr0sl4PB8Ao8GiL4jG+E6EdpoC23sUGuDL9QX3b47zGu1vtAIedxifJwsX3fnCb1Bop
RIiw+oCMoUopLdzu05m/0AwzXuJQvHG65D9TQX/a/GtJIkjLgn9mLp19DAiJqfQ7kdJzJ8+hVeHh
uewzTWrhPLfL50l8PTevjK7SVJw2e+8N+r5EzFBetVTG74pwWo6Leu1/xyoY/CCr192aQfSfYote
5VOQmAUGddQlAmRKUb3Kc9fgVUaLgje5OrhHHbnxfiJkeUwnqIJ9nUqa8sf4WaoqUz4yv3rAQp11
3TuUZNdL+G3XRAPXsovzfVkUhSHy8Tjiq5VgWBNiVUMGGFKvYaTnypf2pDxrV6OZhP8A15m8Jw7+
GUM26jl4LAx5czuth1E4FjYwRP5xeNHWXQ0ISTLnpevZDf7RITiMtb871i4egUY37cx9wNsoA1fj
rFQFdznbdHgRxzf/jxP58nB3C+K6P3EqOvj9y4yFcvEps46Iax1dTv7KCLM40MMkSFHG+9j19XJ7
GLe2EdTReZzZZWxTG4QXP0F3vv2hPmtnnZN9ufq4hRfhsqXcsZK52E4rnCu3DXbpBqr/FQ1S+Rl/
wPpamnGLX3nnU9i3PfZNmsvHRYtSxwYaN4YFc5Kb5eRhrkI/KWGd04cu4Ten0fja+tmHdLQ/0wAT
NPjmdbWbH98g0j5YoKVgcSBe+yEh+4R242Dn6RPKzUPsK5ujOBmZrE18jsavMIBUVA3czpjz/ll9
q88HuA67yggkQiQQLs7DMUTTba8zMWIIbPK980VLQm/YuPov+TKpbnA5DNIaoOZXQc+QWXW9ORcL
VdjCLWza4YVI4ALOcHojltdn9o6pAbGJud0egr5TdL8R68648ysuNmWTpXLR7Si9rMK10dqZB/wC
4C86HuGrYl3HdJGXXsH8xtX6Z/3FbLKno/Yba9g/o6P0NIQvYSEWTKmuK13s3r4ssPQEQErfkmSo
SM5L/Ahh90BSuSWlhr28Zc8L99ataea4rjDnIJalJiSku8st182jsPrpoMW1WakGa2SmClUwVqmd
cHbeyVW0Pleter+2gCJOuwEKkV4P8ZS2FSleIPuqQvXmA03u0hm7E9T/vhyeChQ8oEuXF+1f6quH
wtXGmopxEhFC9VqsehPTloP/Xf5QKlMVwhlkvq7hJ64xl1nWP4wc6+hD8sZpWxm3ue8hHXmxpS0k
UToyHve+UTRUJKbbp6sqK7I7wcOoJUWJQk6HtHih39fJqfCgQqFenlyqgFTEhPaUqiFr/bs2gOF9
lP4kdKqkYU6slF328y8l+5NrY05LOPXYwARj1686PJRy6I22ASn4E9ye7q5EeE7HlGwpuZc8/6H4
QjZYWqDXAan6n/Ou1sBnWjXjVhMyjJBDpyJ2Ffpv7uV3eDXiIOag0rsxvCtbu2ahVmxrNdW4vje1
RLnw2T/f7BIPk5yWy8UTZE1xeQRUK32NA2yCSMVDN7dEr3ENuOeoJOmbE5lTYfFVfHfYWRHjgMjY
yKz9YePF2s1++orbdr6D7joWm6DfXo9RQAtRzJrbOkSNEwkM4IaWYi+XgTooL3u8lA9A3chm45or
0c4p13QI3SZ/NmabmtpLOLRXrj1Szw3zp/RwjK+SmElC5eyseX7+myR22AZzjnHfK/25mtTvvIeD
/R8Jb8EhD+PvzQcPeexwUMjmCfwd1HXaIosqyOVjXpakThwYBrIdnMlAnJOhKTTpQiA0TMJCkDia
ZRqQXvllx36OTKEFlG2/uHmA3L3FwgNESlffIHWeAw7uGB4Yiy+mUnIvecvmdEY0Y1Y3RAJ0ztxs
nFIQUAOvfLqJfG6a4HLpceRMXbBU0llMZrJxDYr0Xsc4p5LI4kZ25okJ2QjC8ku5+/wo8+P5mczA
rpTw6q6EBDdZHaLzmJtwvOI0h6hg3uka2qmUJhcyZRTUtRzeOZAlOH/vXANP8RpLWvpoVZ8rDIND
L+1IIIYCJuY1PM0r5plM0icx15ZR1XODWWTg2SCjHcBKMgItPgncxIuEMYmVYGxTde+6slgZmrnO
wPCo/gkwD6m8OA30UD2dCyLfbA0++qraPiPn67ZDkyCXQHhvw/JznLCxMXve9DweccS6dcN6o+Tf
wEbK2h25giRfzqB4twZTQ6ZVzlXkLprcPB7D5irSNG9pPRP6Ek2P65/x1SsFsRYh9gFq8mh0irVe
5RANQuaj4WtxfwlJOzBhh5a6BvyHGXlxjsY0lTI2NIqeKCy+WsuSSUj1xwKpyfqjwlF0ZtepqWzV
/mMLXWRv6EgLUSqNjL7dV20TF8GU944cwM7u7Bj5wynTu6zRLabv2o55S7TpSXhdEx636sDyvOTN
e7jRhRGdtu7DthpS/Yt6JxTA3qYUY1PJ/abQfxuP30edy6Huo13DTR9GxxYNMtB4lF4HSgj+vrAz
4fJ9CZqKhpFzux79X+NDtIOPfdbcsMQEvG/ZsaGDaovsc2EavpaP8IXnC7yiPJGMsoVjqG3AViKY
F1eqz3N8aLkHTcbR/nkvXavKEVeezaWDsc+YqN6OvnMBM555Drpo9YrhfIic/4/CXS+TayMmUnFM
mf1gIDtHtsiobpf5Z414R6qrJc+WW9AYkjAI8n9okqxnRkPyhBFxIOyfOaAyxUOKsgvZGG7OzCFr
jH2f6CdasHpvpVsZp2RMxsTKUpQgtEsBoctPtTPVpeWqO/5faZEhuIk1MK/BcFbrVJV8y0/eKUPl
Ge6G1tc1uZX07St1jcxvWZpWdG6lvSSgRKUDIIXPocXUUSozfI0KZG63fyDl0+DadlyCx4e5/nRi
DgZMM8gxF1JnS3JWfE02iC/oWCcvDAr8KpXh6xOfo/coHOL/2SDt4B8jtpd3uAksAeVNr7jvi6d9
vyfwTKoN5fWtH1FBDSf67xsebzguc8JY+/A5zx+6iM3HEjgWp0OZdGte+7YPuE9996KQjjte+MTe
ZbiDXflkxZInx6/V/64xsv4xlNPod2BMaSNh9a1RCG7xswD3gDNN9gFDdAKPuARnffUJeTi1ZVOC
u44cZoDG2PBKfAM1H6SOMIY0YFysSuxNq3kPJVmgP9SeCGp8k/Zygz7KxE+lyjrBuZzVqgQoWHh4
AUwiL/0sGuLhq0J099ZvUXdfzo5rtchhSq/6DCeZQoYkjevEnUATo8QvzgrvZutlCGh58jxI77c1
lIHB3n9y6rFCt5YoH2XdGFw2PanEyQKV0+8t8ADqVCZRWZmo5mppznXN1WsHXKTSt1tPESp+l9rW
ztOXTqOblRTOLdhR+NNEqG3FOg1vC9j+F75iaSmX29+wwmhFJiabQvI7gBtgHJcN+/yt3IPUU8WR
lB9uDAzGEruC9NhuDarOAvQdBV55teXYw4p1NpCDV3SgCAf0mfjEoiUINE9QPhnYsZA1H5tezqUu
S4iKkn4N+0JeL1w0khPUfIx9usYISqRyk8Zb0KT6UAjAMVULUZWupyPodvtp5G47JAhJzx28263F
QHgV6dDdc+irR7OhfvrhM2yqMMNfFi17sL9ejsDQPI+CqGerTJPjUXigpfnpdDrhQbk7MAtkzOR8
F6vl7NtkXiesLOSy7Ok2vISF9B6gMO/klxnbt5nknhq7X9dOS0BKCb5BvuchHICUsYjM06quQMsB
mQo/x+8QNmF7Oa9F7s5nnhjf8pFhLy9VwTVucE2YAFSLMPg7+PicympKtbZYESjkAG6ixtDtNt44
UP5hJxFBXDW7zXG9Uj2GgzR5R5lvZuY4xUz2yxsjgZTHKYoC15jKYTLGrD8nrmklyH4PWpFYOHPG
vPVRdePJ4rH6VrA0/TX4cZ6aPXOwIz03/X4KXgY7l9Uks5TGKqN+7ik2mFxS+Yt45VUKtaXwQJ3C
RErQZRSlZA0cekqRUnRKJ155MMuqTZYhCA4zmVdjWEKaAD+trc1DdSAhxZOdq2PJfJPQgS+DR4TT
JZ1FKswXlvGavhCMFZBtklKKoOga1ZzYkgUBPsbZCGcDCu+y0rfBFrViCtVnWnPYzidK3hz4fNlR
OL+DCzPoxyJH236VsmrC8sF69cb7SwvUX8QmrYTfBwf6eexjb/VZW0nIIJz/a9K4vNwiO13DwDAr
GidvgeAZ6/lkDddTe1TlMxmFISqr8954QTUzXRokdYCuW8TXdIEzcbAsRTHq+vazIBTzui8MmqGK
Fj6WVrUOZG90uKWQno4J47zZF8VgI9q0itNSVA0TwnhEO6z+ZqbTvX8qn3M0S18YSB3KQNuYfxX5
np481ikSWilLMY+2cf5Af8Odjfdmddin8Xl8sWarg55E7Ej0SeXKFv5SJ7Y4WQqe4d7PpV2khG9S
wJy/r3datAQn1FZ2s9es12g53SSkbHwg7akDtsOBai1nGBDcSiWg5DEPFuSK7QjKOqM6tXexco66
+AevNBLQLffw6QOc+R3xhO8Keg0zE2SIesRWkjo84+wP58Wt5GNsVcnLX62GtaQlz7HvtxT8fV3U
B3faGo1qDrsEKhSOJP0n2lrzm27xRTqY9X8sPLr192ylAvAazlAyr75y7uTVu0Qjo0ZhZ8IR4DNE
5NAQ2MLtLi1FGO8X4gDHjk4ZDHyeSAkvNc05rxpOWbjzsTihHwNRObhQ/J0EJmWxAaJMZq5yTVTs
/8DtkSajPYZhrJ0/iiSMNOXe6t0PzGEZI/o/oRbYOqUwHQiy7XX3LL4BB7UHUK8bJ9dXXtDTY9no
GnN1ES5G2LWfUe1hMmxbZ3HuV3y6fWj2z9sTt+xeYm/Ob20SOnw0g7ORCO8wsFI8e0TRalm5imsY
Z9VShOMXRfQ/nnhlBRDiJ2qq6Nnh+k0ffpPOfjlzFD3DaK3ZU/MuYwjRdMEEf7zqcTYO27mt0gYe
BkjlzE+iXK0egOB9aoWeud20jankvQWVq35zBkVo7QsVaFzBpmHYPxgNf/QfEYXzr699Oiei1txc
Ec2OIcS/hP6GfzjCoZZNubBBi9P0cMqmtVpXXp8BzBLGbjSYjHUUi77AMJsR8GLq4yJGpsAopjoD
POM2gTNgXDxVflyLkO7kS5hn9bvx0HyW+/Ba1FeiWYFt/T2fiThQj+BQgibvexUzS6rhaeQ+3LFo
zkQjYknLnkSB+r67Ha+iE3NiuxFC+tW1fw19e5zfv+LhjglIrEqLZnd6TkxrG3Sm2KXtIgDlfctG
hH1PtoJjOQu/5cQ4MJMR5jahocCIMJ/9XEB25zfACLD4lgPaajViR/wruIYBKOJJKgQr5+Eta5xF
JcCKE16ZqZyvHFN6VW1y4J2QmtvLYcYUDR4lnbLjMivu44tVFgEIt76rX8R80VNBLShz2VMcPj0x
b1an2/nmLxBOOPxIcna8/C/xXaJRCoO8/nGNNDwhZbIAMJceon/qOby7Hb/cymRtt2prVfjLBFlm
N1Lrws01NgMtOklWEUSz36RZusSftxv9DVYmdrLjPYXLJ7wz300EVuazi88EhuAs5/33IfkokyZu
oc1/6kCtVlIK88gJ0jX/8VC+L8yD1Mp/guL7DBOnPpsFgKVXO6spPIutoN3vUHpnTy0i1caw/66N
iKeazM/dK6xzKFYTG3kQrtN4lggz8x8PjRLpz4OxomyaoiwhrkNXPRx8sJ4aNs7Yg+ba3mC3Num6
VVpRAOuN0Cli02K8I7LQopttHVv2EKg4wJshieWnTMeqf3807ifggntF7YFFKBnxJMBAEjlJGRVj
QECyad7UyCn6Dv+cRgAUag8swpClYX5mUYrpqr0U3IfjYIwl/9Zk8+E9MaHc9Fp7qJ3UtVyPF4Tr
ik4iv/097lrRH6Lnwa+fgcU8+9omSLgNjBripPV8ZI6nWy8he9sbmQ76cEwBfpTLJc8PKYULWtNd
mpCMrkQu08+2lx3efsX4zCBQ41720HMyd7/4kKW/KV3MJCFxc3vNWlZsLq8U6ubW1mv3Hgk0QnVs
AAKFi3v9b26TMvGjDTv15WBg1PRJPn3qodIfzir2vgAbVQjA6pQeLRu+ouCnvObwccgM297rNJhl
QQjYsfiJxRMZn7EhQdAy7hLF3RNevWELMcI6PUwGhMpkq/Ebo32Bw2hR45VAaQaVqaQvOlsOmsL7
YvMna3rZFQqy+WkrIolmIqC84RtLIoZE0pgdiY5En9tL8YqA+FGX8aGAxY9h2LTQGGQvXkSt3q8F
e8mcUhDZaxZb0ZgnHFMFYzX23zOgFPE81vmtwi4+D9BPi1V6KuMgvvrACLVAqkWS3wkQKcm/DcFO
VicNCfuaPtLcBKwAtvRY3Y3nEZ1IV2JlG1SRaIkRiAkAD04n7osSPZ6yzKc9yGb8elpjK6J9pHn2
PGDPffANShDB6tJD3XUwVQ5fGHfPNlptMktFaISNAgK8PiWEw9XuJtl4539X77MIG9DPZ5FUefjn
aOxzlzUhsCVSPCI0kH9qXDUVx2gOiPcDypSZmZDreAtrXx5iAQ8ZJ7LYyuYgXvNzC0Kjl/rt1ffg
qgmtWWqMl7HvVcjm2Q9n6Pl5eqrhqdMGo4PI91mKUwry8Cp5bbIwnwg7wrtJ/HU2H+7xb5m+bzUV
RMxHQKZXRBEs6vTktmzz9AjMgr2SB5EdgxLjuu2YkdjwPMn6PA7qQJJ8e5L/Rn31hk27Eni4qHlc
2U3EN7Vp5nKJgeLAwsZwt/xYkg5evGPY7NrShwiQZc8dByRBU9TWs7Ps8DsuXZt9lH6D7wa8Cgh8
oHpwHXY4ABSu6i9GJexl1QWJjWfgBw1/eRCU6QvtEX0IvV3F7ysliS2bFgADZmsp+87Gdj4cqIOB
35Ut5zi8GT5zBY6r59qYIB3FZGTncH+rWNoY3ENOAtEP4lzkc1S3BlKJrYx8P1PMA7i8LoduJfRF
dM35GhoyMVkgZoD1zu1tVcYSl3+HEsKf646ImcAO5Hwy2wKm8ClvkYKdBkNRVU+i3sfIpkXhOeiM
xF5zYitbTl4+biideX2Xe2bdtb4dtsa1KSjbg/v326vX/2gTDbHHJtxcpJ69m+ZcHYtTT1uHa8Dx
sBdpb3FEwIM4P5YLToK4U+jFFFvkvVKC0xejfnK6A4AFS8p+rN7dm+uQCtJKFrAkORy0AvW84fae
1f0ReF9oOmh+G4rRGqKKAqX0JpYmv3NsSUBQEUiHUDcCts/BrZ0Bp2mx6XElQ9yOtPx0jbkUA8Ck
yA8BWDUTBDQFbTpxQB25npO2umXjm4QYcw6be7XUPTiP3ML0eYqBteUVHjulvlL+EgIsDHzm6TEv
0W9ZKgB3ED/MtB8aWzQDTVIgn8e39pqWZij8Gn9cizS/LsL/Gb4tL7vmnx10cnKo0f0VhTQu4tKE
+S4rQm20875SWz6BiPeQREI9uR+MuQYxmKaJ6S247V8qqylOQqxr9u51ihdU+Vwflop0BscnKNCQ
I0obD9iHH+MBjXP9uxghR5gFp7Dh5PjX+/EVPZCTgwJrrehhNJp7zcJO3FpTx0jCJTp+YCBuUYGk
9kXIqMU5WVXYSaK+rryJgeTdEBSlQY3WZCIlLkS2lCWpmFGzp0vGz6hmT1kbp/TncrekShchPq+2
wJOdjW29j6caHKdzb39hXEj4lheMxzGszp7CVX1gBRphGWjXfxk1h6IRRR/Yp2BuJ5dEn1rKXkp1
4FHKRkWmCCzYXOoye1hToYepr0IPuvfRm9njldCemN7YKeOL81zS3H5Jz2pQH1bpdQhfXh2Wm8mb
+Z0QV26oVJ+q5SakTBjMZyaopR7ZoN49v5XgORl/jFWOT1cyQji2x0iN+tByJqoZeaj6a2fUjy+A
Htm/JXlSEDUj75e1TYoJazOvpaEVpcHuXZPRx+j+5Qzg/W4+J8n/6DmmUPo8pDc/O+PTlij3iuCS
Nbqf0vRi/PTR7+moLOlVPGH/CsFIMzsWe7i4a6+6kV7iTkIn1B9Fs2r+iCAS1cd7nBrZflgz90ky
w3mYky46lORxZ9i7E7apZxxVn+IlL0Zo7i5QXJrDQScAnEB8D/Dc4QNiDReyN/ymODMHWDMZdrXS
kOdcUiHJHzfWoU1IZv/f8EUM6F5FiZIBE1EupFo6Q4F8Jd/kc7KKGExcjv8Jz7YDqty5V5pgSC4N
pS4bx4zeHMxhpfU78yU1barPyE6otYRDE0VZuHhe+C7rBRz3Fr9nFsKgL4Pdfj/bwgt5+izaRuAm
pkVLtfzrNUgezIIL17G6Qa8tvS/AfTu3YxWojhyA37oHjE7L6rj/YVf6sB/2yViSPypnBxfmlhdL
ENLnM0qS/VaHE75eCB94bLX8PppTxdvgt1XNdEY5LlWx3CddvObvbMHjd7WkwxbSsgXeP+FbLwft
eZ+KvmMUoxFuNJj7dVZ6wfZymTYAyugfzM3C0iYCshfcnwabfe+2P7TyLQgOncuN0LJw80CZ+dPd
287Ak3zfhuOx8x+FsJhNWJiXBijzB9Vdwc9IXfXcTAVQ/PCeBAnd5mO1nobu7BEkJorb2HBc5t0r
dC3j2q5AcILPXi73B7U4Z84jqfSJgpIrXSTaeRJiqiqRwfnFb1J85v2SSrVFWLT7Gof+cyLvQI9k
dtwfWQe64A8V4EzfZGFxC7RRZFOW2wyUe4Fb2YqyhMnzxjuieTevrTaojqCunTsYKaKRcJTZ71/s
jEQvw9PS382/kI3Jy1Guc7bojVdP3P/vErwxr4ERfqnX60ZPI8icMuh39UOVVZadol9Gvxdy615P
BL0LLNSvc60wpEfGUjAz/2lLOF1VvPoniJu9UXwJsnLp6eWOgw30kWawwk4UVXeG+ueXE3JNDtqs
Izh9zPJV+LAYXBSC26xzrQ8cLSUyZB374snXyhydLSwPkt0l877PigIkJQd4tA88J55l2cnzjqlC
kJmnD7p66oLmCWKq7O647NzyuAndWgr5JfG8yhwf+TQVEmWSMne8Md16965h5BpBP52J4wKNmwUf
3IGnjffqzhvpL5k2SuVBoxuxnQUgyn4EENzDJlrKHIGkgbtteN0XkjZmOVb71vMmh+9lrkcl1ppE
A/fqwi+DHDt24AKO5ew4kRWyb3qv0JB2pXGvt9NOgnhLuaF0c9iZOZDCesl5Sys/fpQmYgtOy0+7
yagacEWkHEhV2iG/M9/ymW6JdZy+ZBuVx5vDyRvPK3lG6RV7HYbtNsWVgaK5B8fKHiKDccr66Zyr
yFXXKSIYvBfFNAUrOLBoivj1SB763m0BckB2G/kkftp5lppp3EfVT2yn4o7KR9E/DqietE+TyehR
62kEmm+KlITRtEnNP2PADqPwfTdW4Rjbe16rEakc59eAy9QzzIECFbPKz0vDlqRER19vTWLxDNGV
KA8ogPCBCnyNwqg2Wi/E/EHRvY6aRMNYysven+BwalS1N5j9fr7n95km7EgPtXWpcr5DDFNisLVm
/99i6px1ofHBIsjX5Pw9DmNnPZsWhmXtKZAciFLaH2wkGAtbVDi9ezyXFyWZmlcOOFrkmnq9GBTW
kkqN92es81nO4Ves9EIU1ng/vF8LN451v8IhWtFtgTm33Fvq+OHvb7C9JjaUyC7l3OALLt4uP52Z
c61giAJQLXjVQ+/kHqJq7+AK79DDQBqYpTBrkzV8PTBLU7RyH0ASQiFEwxqbIZX/PI03c5wxdwFK
15INg/DaYw0dz4QnAX1kq7BJDW04Ut0wRljO55J+lBacHvgH7x4BDR7kEKmEl2e7pp6x82V8igHs
e+dUG7fBxFBHb5EYMrgZDPsqH8rwfh1Em3vwIJPPMwJ+i9Lkg+g9JF8qox7EYvr9m2blfhBUAsXh
o/rHRsmSJJkbSQJpfJjP5uiN/e9vxmid8r/xz3bsiY3y0Z/tXjqI8ROL8VdM8cVVkl76M9u/x4kO
3Ggh3I0Rj1S3T8KLAK4NnDlZrTjwCu2mmIaS1j+R+USWYhL0cRdSRZTKRcEonTug6BJsWA+PvTRz
PffDbCovOrXJ/hRWnU/OvGCK3q860EnDyWPom2LjtQDpE+u7lTqcYUDJs740xVbMxy4cReylMJ+d
IPBcXy+b8K+2UqDNkfDzYuVjNik5RAQsa3S9RV0q0cptaFi+KJe25eHhD0UfJ6x79xS8He02zZUK
4UI6BiJk1orD+uZLwKv2wA1gBtyE6rF8twbPNd6mdjzQY7gBMO+P/fJP+8kJfK6z+sBRL6GQALEB
xQStuWjg1C2Yihz+iN78oFTCKxoxFFv+O8MVTwb34e6ivQYG1OkSjcNEzrQI8tSn6t/3MkSofUOx
LzoL0uDGtsTQdYnKq1uRcTfxN6Mkx3Jcnx0YyqHySe4ASzOeo0X4xr7h4LgAqMwxDVCCvXJGh4gy
gr9H6WDiaRH/lgxqHSoh4mUnB12KChYNLzuYsMAF9uQ+8CeoT4k/R2SBDy4eZF/olaNAN0JIgTs5
Bllr83jfmQ5ReXrozUQC9CCvGVJHAQefHwXFhI8J+1f+rRqs9GxWOcmn1ojWmupoF6ROE2yWH6Ae
0jKyKA++PVKZbW93lX+Zm6gmtiQwYgWpnZod8BfmyZ8xjRloRXkUx2CjZgTlR4Bfu4LW8tTvonqs
/x6D3ch0xiVmAD6+cmHgv2uW85D9Rv3GPGwxUk8IZHo0WhbNp/Mjs2c2Wogd5pSu72My8yjGJwP3
3TvRyO9dr5a+Gt1MSep87KLUl6c/nnWFW0sJrdmp4KXLecSEwkwEAXv3EUC3I6mjQaykYlmMY2GY
E/r55PonixVosWiEysHNJmYQn3TjeqOV1NvM28d16nNvvzb0c6LqlPBtKA/qypLpn4TM/+vEhxJr
rKT2h50Telnm1nvHgZwwfJhLCQzut80T/CTFPo33mcN4nHJPvz9WNBZUwshM85wpg/OBUtJ+H70m
c6fMvBOzv61eha3siDWh7iwSYx7GOckK/esJtCUJvSCqm2c0FiRlF77SpD11Tx6kvUqqW766cowC
fHpPDAbecGTu5mhIONBzGtUxoSUYXBXOnzPoe+9oS44YKhXTPbLTwtfp2ASpZsefzUXjm2KaAWzx
WN2bITbBo6k3fehaJUyWv+XkLIxafpREPLtnMphtvRQ605iT+gc0mE5HKMZBlBoFjBu+K6d8ckai
iN7//nuTvMDZKqCuSyfkK4NMLqdTjrqcEVQl3tirsy9SqKxeUaqt1LhVD8NUZzLTOBmIxMWwF9BP
yKkeE7OCgnPV+xSZdYWUh8ZrCzSF3b4QxGS3ogoWttz12ro/BviOE5WgXRvCCDRCIYIxDTuRp5pH
iDd4smFZYg28juZMOO/sCQ9geNNK0mIjN66bEuSa3wtHnwmMb0txh1s+u8WR46H5Pxp530B41pmt
0hbQuIkMewBzeU7wuVi5euHHFzZnN6Ri3ZLYv1SqP1SJm4JAM/5BG3bYUsfhitQYXChAutZ11cgL
pE80U44FgJZ3sKpogse1HkRSei1apt4dnfA/ZFyUBaGwESLgWVd21gl4D3RJEOrCQi0YAUwI/RK+
BV1xg1Gpqyoo2gif2idnLlClt2VZIivCJ0LYcbquogAdQEVSQ0C40NQ5Bm+aGa0dCsW8K2coxgDv
J9/gvFm504fLle4vbFPjAuZiTBBEHwQnbcDTFGr5WIA6IcmiI41UUdzghQPQ0cS9L60Wiu2evs2c
EB7g9ZhvH3Ih8w6ft0G2/R/9364mUAb/rJg9bolDA6PujaSYGat+URlqa7N2daCrMuVIPKHkYera
pL9g31M4liVZtcLe57cbhYxjeQWW8eO43tvNEyJGuMuAIku2bvy6/voDT4sVDOU/odAIlQFMYkYT
S39lRLFL5cZ10Av7m/HI97obxscvbHo3bzTQTUih4f+AOtHFy9gzA/SRVLbz70G9YXVp/kPWPpbN
ljNl1uCaSDa/2xQt7D/JR7laoPM5suSEDJmT5MbKECbMWcFtONY9xmpH7ogM4tTIQn5CzITzN0Hv
fJiH5UjR1Us6PGg6P3kAdwGeY+AZl9fnuvFBb2FrYpgBbK4S8+l4dC/gxlVpAW1X5Qbi1hKPRy7A
jlp6gyEO5pGqXi4DSlP+ixy8Kbrv5P0lZ1TTrSrKfVsRa8SzQaLDW4YoGJxmS6BNQUpopyVvMO1Q
A13DXvupgwbOjTEivt0gpyXKAyTq31SSsFwoOlwHdY+6kRaG57Ke/vb7ZNWt0pVv4tV/LH3CfV1c
2qOVJrejlOuzqMmUK3P5X+lFBECR5c6tsHBokvKOCIqgtC53GVHAjm+fqAlvbx93OH7W+kIltCV1
D0aoJ0r8VyjJ8XimKVuDXh8auvuP43p0/m+UuobhG3MNekUiR0QJDnCXfjKk4u9yQZbCrWNfBdFC
EiqROrF0ju3/HEZcyr0UDecl32cJf1LVZdJP5fsumdnY/HzeZAbNmWUHJfk0tmpXdViwp5uOFV/n
yHn1UFlG7jOMTyWiKdgVpYEZls51Yd1mrLaMuJZvxw2fz2liRxv4zTz/3ULtvlbcr/MqAjQAJQf+
YK29SbNnXOJmlo8D+4CHtgLKs2Ihy6Nm82xsP+69Yy5sB4pn+3r9wKX3R5pXoaFJFQf3d/Fs2iHE
0bM+VVScsOrHjr28TBochgXMnFiG7DddiryY0k3v/sjMj6vUMK5Tb3dFpjPKBFTd83iSfb7ICuWa
Id2NoDjkQRmHFOIFbupM7Y6PGDUdUojxrbqwL29SK0AiOwxYCZewzo12wqG0x4Mp0fgsZRXTx3J3
Bu9HS1MY3jTmj3R3duUQw5WIXkAfzNweGocCQP8luSf0yOZvJcqHAe9hcEiyj/E5hBIPCEWEA3CG
51nd/6Osn/D9E9+AGwg8XS1wtJfplOHkYb7YAyM3C5OncmvvPYz/GLhwZUt2bgnAq86thix8Ee7P
uDth0RpOfgGn1pFy9vdDZBaM33TKdYKIFP2/FnvdFS1dJrrkbgHpGslniZBQIjcXcKM/LzEVMK4r
70MXT6lMyLTYvR0K/8RTdoBLJmhAjYK2DtZbWtqd5qy68q+Vutw9PrTco4XOqpct2S6CbJE+YQ0/
NeAUvHCYCVQdgmgRGqLSEndp3aP5fQkiZd5ISBkPYKZMY3titr7eY9KievqcLqJhLBF3jX+fRJf6
laNndEGRyEz2IrBljLDgob6z6oJZ/47USwgT1uWmZRPFbnEmcJ4Em9zEzlUEUDi5zp0sTV7Y+0mX
HvUwg5vfloVPpEh1VEo8ZEr3CB1K45NUy8G863KnzhGXvCT6h7a+X8RY6bqiIbjpXGzqOAh405md
4I3SW62OcfzYiyQYUrj3MWA9XjD1ABCmI6f7G4eaK9/k6kaTv/1KAC148dPoZpEJxB5Coz3DFhZB
WXYnRZXjiEKMBuNoY2NnWKVcgiKlcs/OPiYCmPyZJT+H6JafBKVq2I4Ik4zy/HGcwIS+H8bYKwX3
lJLMoHP03Dd318jhDSuhv/csZyHwkHzClI2iTby8xXSI7+cu9HCPZOVOwv1hu9quojcmxqIIWlUH
HIvGm9Yt9V0LNqZyHGlKnveIpHfILDYSuk2ivP+PMq/MPMZMm2I7uQbC9AOuf52LRlBwJbPrmFY8
4ZOoAPHnyHWKMSUxJI2ho0ttSMyA1+McYIMk76TCTeG9kVjMwRPzXRzfQyAzl9x9Pi8QrnebYLxu
z9s/PfrQ25dvFt2erE7xYKNEErxqhg+h0j4L5EJepGyyirrGDnhwbiD8bcE/PSXX10xXBHO9IPpn
cm2+j2ZoDZBP+bTluFqyedRcVN1RRK1BlGCLCtjHYR7t4BIJBDl1kNK/JldqcmQ68Ne+GFY8ys61
5i+x2lv55/W5ZcmGYF+/4sUXgNDi16Dv8BbHniqq1hbSD9N0yokp4kzG1x733sslfmsDnsco1Ob4
fXL7I9ToLy63DGEQ8OItoiG3HHJw/7qoaRIuNWFHT3ik6iXeCzUHh/Rb9E6JUK04KIwQXQKwBz8x
MC49rpaYf5BlXRawIFmEELnS8++i1L+qvP5QkyOLOFhKp97RgNErTQj2UGQBQwEpg8KHAvym7g5r
VA2rw36aBLRQPsh60Oqr2Z8JunUbHv1hE4tp7KBnpAyU7hu4i3Sbh7K7rYdv/XImbrPr88jWJzXJ
y3mqF9mMdsXfhp7inUNAB4bHhDqGrtXfP95JRZ74CECimyMxKcoljNjC7ClSEKFCMHWOQg+JQqXH
OlaVfsqC5PyPP7JDNrmq+Idc6VV5H4mjVWxHRzi7NvWcV/I32uurmCDHqH4u92WWBpXL96YRGioI
n2gcwUexotke0W2vQVB3R9UZbxJAWhFkNi0clapcXxWtf7nKb2dK56NVKSyU3N51Momtna/kBkCO
rnu6+kLfYnFdc+3B9iCzfm/DBdrcfE9jfmfWm1CfC3HtV982lboyOS3CULxblHNy6sYlGNS4fGee
RnbgfP7G3ChDr7fXr0xF8Clmhj/Kgg/ssMHediaNkjA3lPjYY3RBvr6TcSyU6dEYF7gl5QWZGuxy
9yTLtU9jmc6AtOrsaA3kIzh8+Ut5mN6URaCcMVrpktzGT/IjGG4rb76UrmovqvVwiMqFFeB5+MJe
Bb+AA8RPWG9PfvSKxW3GZ1OcjJE+OvscnA5RCkOZROcMlsvXvdVq1pOPONz3EqIsWkwjx8SFiG5c
3Gi5h/uoXrA2Vu1HtU6p/uLIDnczU9RYbClfWnZpjy1aJJFAnnQpo7pK9OAODZGuKAtevv2UENs+
etMmoucozr2JB6PVATx2f1j0UoHWIfhxsfbSIJZYqj/6JjCS3ML1k/++i9pd9MUraO7BLFQi56KB
ccHK5XQ+gkpdNOzyhw15lJkfEX3/MS/KWhIn+BOYgLuk3S+jjM00Znxd4NTxNrkhd5psQNuAm2FL
FsAhXduOtwyrEempdvmSh08wVJIZxrGadYkhVI4h+9YDwfXtdHdqM/HzFJgqESWbknHkCUuQ84kR
Y99unrIeQGYVO8Iur8pqYaF++jy+yb/802H5+RFKm5heRvDx6KyV7QDWKAF8gzHanSWy6Ykcqr9f
zCTJ4VN/jjGl/NiFy+5QE4qJEkiVrJaHvpkMjjKjSkyBcd844bpNdGs2GiMqgadC5tMjV0MGg9Wp
h5H/OezR45jclajaJPv01c9TZzSN/RcS0NhdMGdZHv00n+cuOsHRqd4W0O9mZXfQovQeKDvojnLG
losCfdm1Vz5tGH8wv5VDfzlvnS08131bM1pXw6AZfZR08tq7X6wlLKT+NIqB2Di/j+q7hkhGn9iO
RpplBfWp6mrXce46A/k6AosAUoYefEaafn6tNDwr8+vJOT/yIfax+nnSDauqtyTBeQpOiWKA8Ktf
0Of0qXmE+9bN4ZFOGtUxXO/fQM56sfeFmvE5A4pb5W60mpUW/JSlihSTJ0IC838H7sq4V0QSZGOI
BDjgZtyUTdesjKRdoF2WRBy5T5/vGX5Ks668Q3eUC4gbQaRqPr6k09ITzCIBdV9pbbbXrlPkePTK
by/HPIAS9M/Jj0L9p6/r8vz/hRdnTJxVffkMQMuLPA3uYSZ70rYbVLDfn+TFE8awCKTjngHoWYjP
RrwRIsRueesPSNwZMYyACxUFMcmZHMVBET1yzZc1EtVPj0OJoQLhuYEx1m2y/NkA6CIvpCkQkB80
RAAEQZ6D6V9ZIxqCixxH4kUmbTAhG7MLwRjlPbfnwgI+kgaxvZhMd6Bzs8FeXtv7d7E102xkf8Lg
1/TuxOHqrT0TAw5tc/DpmU/sOTtF3YuU6GyiDgKEcGiGAFl9PWaAWQyevXNq8B7TlU5ndcq97/Gs
pwwxb57HngVTQnS2Ydg4buprY/0NIFvA5z9+gPU7ksO5M81cMjkTdzrnky+Oc6JU6C1kVNwahPa9
eEQVW3z81yyJ3yxf4dNXnlaiphPN4DoyzEcqCd5aP1da0cgUmxkjc9s1D5rNTJvEA8GHCOMgadax
4XBWKtyPxwT6I/j1rrh2l2SknE3YrpbPgDCzn1YOX0IFtQpvz3QM5zWCnV+kWnMpKVJf+AOOszY6
FNlRIq0ldvCYZT7+b9hoMcbmVu7GCrqgMWlNUbYfc5D3uMfWpLFDHuQSBUPv73UEhqb7vYH/to49
o6v53Aa58o72HefiXnPHGt96X9kidTE7yBFWcIeLWTP2yKbKS0cG1ID6LFDOWsPPwz8BocmJt9/U
1+7KgQIGNnoAc4WST05SlVx1mvPiZU7VP70QoOBfMLsQQiv5BqFQ/iDg5mS0s9ZZ0uORsU6Lda7Z
r4iYfqu2TvgOKAQLsdv6gIrKE1CAL6SVO7SdW99eLfTzkDppcLnzCHu/VU+PUnBGUm9WZP7zF1kR
t+BsOWLjaDkwznvy3NSbxcIW8yfQjJZxyrVEnv/Lt+MVe2v4wObjviy4oe04Fpt9ODGfQV7oT68Y
nDyAAPmMq1CiXVQ0bTsKRQbQdnb+0OkfPL9BEqXnB88ynkfR/lgofKWJAtErEgkmfjqPQbdW9+O5
H3DSVNoDEgL5tO+jT3157SnAe4z2laxnS507Kgavg9loOWI3PwdIM0IC2iS9XJ1QOSX8nZV6IVt/
ogZzRx/tU4hFedqEhNoglOKOMg+HOY2lXBO0dPzzP7xAkx+H5yr+OYrPxguv/pDMxhBkyE4fNtSw
HJa+AKCWYvupcZGDILZLJntvge3iutLqxR6f5mOcQFjFoxqiR4qT6g7hvy8kJetf/QkEEhbyKc7x
0o+B4Y10aXEdvD+LxjunVkMSsGNnDgvucYTsuuhSnILTFn/mEa3VwcDVMkYCsnIHQGbeQInnIOdM
ZEddhoKV4dnwmBqBtznh4Bgo5qlptnPYdbDHrwsUib9PKMKK6L4gZwPiKrwreViYzzUjB5bz51DD
WWid/1OV7ICiu3UE4kFQ5CeCT/Dlvi+yzaiPvz1jEBYcFqSMJ6XKIMD1/AprbmiOsKA92Y+3v7Ds
zu9AwHCDQUal9YMShDLiymRTRbdD1uBZhawaUfxe4NPU/vDn2j+dqDmq5TQErBfftCBfTfZ9zql/
iuyEyAkzhA1JuEvgh9LNISmj1I4E3ugludqxPkPAMGSVk+o3AobhaLl0o7HY8sTpQLeQzPp0kio6
cLkq4RVNp2s1VVLUJYDIZ9HO9BqVhXfQc6fpp+mVYQNzqZBtF5+o1LSdUc9LtZcP/2vgMVrDlikd
UX7fWWBEjBu3CF5qwBLkzntzyXwTIS90+gHPp13GUChMNHNyXuB0zE+JMGJ2oxf+NoRsR32ps5qj
m/kYEUoPt8x6FqLqbHekySscUEIMePjDwEgbPk6w6/RSUDpVcRJq8Bb2GMs2NCE0aHkksSGZZxtl
XIocUazv6+sk5Nmu29s9GhTrcmKDUB66kt0QqIbBp5J8BDHahXjXeSSOqhzxRbnQBbS9XYRKcNCd
yE1o8sUYQbpZgj7jxmRpegBpUhqKUrh2JhtVN23QgepdoyA3jvOiYkMdon1RW8u96q2CkAUxLEnM
pgNLnC84RQsj4k9s8ac2/WtHo0P2m8BjM/uuc92ZDhxld6Fm2UbFpjqApVfJavOFpONRtqmpXUUm
MdZFQ7jTJp7WNYF18KJBOVN0+rOm7i15q8EnDsdVpCB16YdCW8VEMzHmeLXGUA63TauXS37/kA3h
MG+cZ9mV/AE38e0LlV5mF/JYDYAkZnD0PCL7KE6bGkt3HovH0uSRfKw5420LLmnRNWbbUjLYSjqK
aCW+CdD3teFtvS5k35wW5rqkSRhhbxEGdGSmICYKFbAHFOmP1xg9ghblkdfbatKeHusDZalrTUKO
+OIMABBbBKIj2O6eR7yQ2/wzV1QYGiN6eJbidRgFZCVgqFkoI/YWDT8/jInxsQagEvOEsx00KNzU
4T90t4U04oFip1Ezb8owTX8wewJgErbfESwxFotYLJ3r5O5tw40sZpDYuYZ7dIPs7P0RF90DN+Cj
duLvojogISybGy7KuIFR6RXPpqQUki/u1XGbdwDHjS0TLybEOdLegdoZ/FPYAYdoMZHc7ZaZyhJP
T8We1Y8xpBJDRD1I0aXs2qGRJ5TskslZCbZg0TQ1Azp+toJwHniESIx29bGi54jodf9wrFYPfVll
upWCfPi8CKBK58dS2aDK+nQMOnY/xAUlwbo23+MCfR3edzuHCtfVmsoc8q7SL1tzgpkfGhJGyDgb
Mo89k0aKlsq1JIgL5dyGkcNpDFKA4VUiVXI5KXZFwGrKcTuVB2gnIxWF/8MvpGGLUPa1OLDessTn
+VN6IZ/6Uofg1zRRLZVA4jzBCKcL/0yYvOxeosXR8PgHVSLOE49zmtHszXgx/U6q6sdYnTYcbX0X
Q00xydNYwKfaYmV+XetJRekTrFRpcZvccgQmGnJkbimJ3CTi86Gyt2pqDpJ5R827hl0tNWH+hHgD
lo4hRQVp0YFe4rBP32eautqOvgaZgKDZKubE8JOzm6Q8NJws5TJgTcYmHAbvhz3X8gRoZQgzSSQb
V8ymmW0KUaCeZUMTJ+dwZLxss/TRSF6Lk9JiLayPZpxkFT3Jk41WPwrOEspPNH2bEzagerQQ33f2
5ppwo5tjaLXJFRqoFxokixAnynEmqPManHAcaAMrXVTxutPBDCoRPH9Mc6jKWQu2QVAgPM7Br2Tb
evARjV51RYZkuz1RGzTsfIp0pvG6N0NBxAJrbQZDniU3KxNDkmfQaiPjT5keGnhgM0Qywum0L7MM
yZoULvoMHXFDTFMZbY7aPWF2nYM6Pyg7ycYoOcUITOF7HeCnhTqUhGsyMfLsvQeK58D31qw0mkRD
dAuXP0l4GpLo9W3bqZBUz3Xuoz5X/xd1oInOj2VBIrvvDea49+nutnVrtndQO5m7slRQEAzeJRBw
XT+I1x2f05DxQMsU1g+/GHbPzBJ2LN9EgyWXZqUDUINo/2rQnh1XdV4orn4rEXZ6jkdVfsHesNXZ
6ifNrSeGC6H7O7TMYqZBtr7a8n02aitLG6HLrXA6kpIewiD7Z319UtNN195s5L+CoQlp8lEP5/Kj
5A95TqFkaZK1iq2sqiGytnG07GL6sElKuuG3wnslQpfqmgOrOzxeFTCSJV1BuvNvp9hxCskpauZs
yQkU+7OM5yx3GKIOP0wZNQKuKPtrqIFqUARZYDRuuH46ZGEkHm2rf2rdsM1jaCq7HemNcGdTkMWZ
mBpQChTYLvT0WsuRifxVXgslzbJC1wkNqXrtTxdaZouORy+8WKlIyZXRr1U8XfQcX5Orxk0IVEEd
1BwQPA9IdeEqiPtC58CzaPYjx6xpKVCOQHRMBjrYEpQOI94uQKcak2Bwn0CrRwGYPxiqmhDBfbOw
Rg5YwC7YTyay6KqUABeTDrRuAdf3GCuUVMWn65IQ7IKaH1F6IcInrISZKa+LtRswGOrJYG8cQYh6
oMBhmdBowpks+EWQBEk9WMHZBwvVmgagMtBdEJatspdFvnaEuUeTNJnTaI9aQSxEWV5TSGsU0gKg
N2o2eoF1GuJJfL/U/+fgb9FKRu4cC/3XEXMBlje+/mhnouglYU0qcHSI3aKwuqIQxpaOuYvltCVp
qj7Yujd3iPHzeJa6Y1d4nhhU0wq88AUC8vyrlOXbCdD0iXXQ/uSax3JjY7AKmnl3pj29nz9ykrk9
2bFhrf2Bwzlw+On0THB1hqgMwBv2mtgu2iwUr0z5BkLvtfFiQo8nsc1vQS1LuTl9Dq+/mj1vS0Aw
hS++Rv2r1lPFXagp50FmXFi1hZjyC98a1yg1HJL0xvQJTD+Ap3b6CiC06DwCu4NDcoJEFUHkjWa2
d08awTgx9twagrt5dMZy19wWNTspW60FJoUpJVdBkaGGj9DIwo3dza/S3uQiHveTmYodRvInp/Vd
pl8iW0v6WwDgRoSya8RgilI0JvB3nIOZ6tfGXVO6bGg6TKmU+QPdGXFdHcDybcva+qDmPfAZxby/
F0m+dVFhzGp+iQJMYBePLrAdY+t8NIW/CPXscuEdsv884v+dy4hCuHTWb7EJ9YWk3h2blyVg+a4B
i/dmTSDJ5OPn9JAbulDiAv9x4jHcPZgyTgIMBQpRytdMc1E87ZtverwnhA8Jp/pIefWks8hsiWoY
PaGrR3nJLCR2LtCM24VWnL/sT4+rroz5mi3D7g1JGIhElmIiH+2cnZbELN4RQACzoiyHCjFUR1zC
vBld1q6OplPKlc7Qxgdoa9nCFp+1ns7uKSrKI3/q4YzHYGn4VQ47CpaISommT7RduWsV/2jF/P0d
WoeCuwnHZuWmuYJF6vnRlvocanuhN7hAxOZYUIWSLkt1B8N3Gmnw2Wucj9+n7Ffj1q1rtANwUNT2
0/Zw8HV+6gw+FJ3LfoUMaZPFhO94rkUr4Rgu2KAd9DpYSxVVJQvOcX9KbySlwqWTECIT44Gue8fg
Go7LdfvSY2RUd3m4MZ5Rfd/TJizrKhtB9Kf06YjzhUg+GbgOFe5mK+xENXhWFbFiM4LyQPs04Fml
ujamcwO+MWwTRTwLN/MON5awwU8/txRm+6pmjvO7GIusrowEZk5dudKLpccErIIaQ9Y7ubBP30Qi
Jp3If7AsN7WGpOUds5o+0Q+lcPQKnLNW/NT5kThg+gXp1VGI10FtH+bzpjZoiWj5khXbRmA2pgxX
FG1SBQYI3p0DsMNNF1K04Z8WYBPA0rhSn/JMwOYzrKy1c0cB6iLmf5AZ7hXnGdPJMN2aoq5PEN1y
T97ic0xtDHFhsouJl5GuiLazso3zAHu9p3ynuS3KIz1W3aNPUs7HE9bp699y5VVke2S/XDIpbVcn
G7tquvIBUhGqEhGG1f9P2pPdHZZ8v9A7u9xxZbDhyAsjjCpNx0DGmbSigvSR9aKqf8BhJRRF7mQA
RncX1G8pxMNJSTnAo11j3MEzFQU0v4UQG9/8Q/7HFba5BEpAh1/L3vQPskT44VOYW7N2UF180Q1Y
oD3xXi/NnxLdQqkBVmDiv0+y1Fd7H3FeTc+n9PQGdnWY2dsRmTSuF+2GZY5Xz1bR2ShcXgUrQyI9
nyjYkpweUR88824ywXK062FaZMiDGvr+FuXCSkVKrastd62WHnwtsTRESIf/jL7qtyA4sZU7Y3X5
jMWYNe/OaD47Ouk/p3yf/sMnko0kbmOA2wL+KhePqxk/aQWoJeI0O5KhFODEX0bXFQsn3wScJVBv
iVDsc4jTIvEs3SK+lzpTdkLyvb65OC8HW1wJx4sNuYsScNCoKKweDr229k7pFuDZj2imPoXBnij1
9d67K7JxYa/gY+g/8w2M8m/5E0SkHmW1ttYwGvgBA07wMm9ffqtHeEHyBL+/dpDzwPRjzCuQSqtw
dKmFtW9OBpPrjUNRApSzuukMg9/NZ+zArxL1GAofUgJpDEtiilVoVbDW0/tAAJmqtrQ1qWHgXHNA
IFvRMrrcWqw5VN5mV83jFf1a63eCa2mm9kmJ8tQL+sQaucDtteNT7MkrA7aJXpJ7heItQnp+BxWR
2BOlgfxQdeN8XKaFLhSBiT2K8WxCcD7+o+aLvp1f/ytP/TIns9ZswGoQlPb/uMmyDciD6UqwpRfd
nCREelNTnSZQ2vTZHONez2ssO0/nZOV4VtxSzw+R4e1XOH4Uy4fSXLXQEfUeq7Jmyh1PGKLImb7f
wjH3IfeaVFl1LcgC7NR6PPlRwMrRsy+/UwvyRb8+uMQNYVNlO0GYm/iUnWgRr1LTGXBm1aYas+yj
WqaZYct1iauDOTFnR6Ofep1eGyTc76n5U86WWg+pIRHk2oIzV1TFfgX56+asFXXkbpJTbrzjdrxB
epOTzT848bYMfm5kYCfJvdX/CZwU9pRDwUKDCHCAgqqqN2ML9nX0GuCOaVOC0F54Op4vWbiqhT7O
kkh818dox8n0qDeC9UqgqB5FzAL4E241616uJtdEzhtWey/CnuEnh0dh1C3BZ+sMSKyfgD1kbfr5
Qo+3Dspigm9Vuwy7WgaHF4Iw/6XE/yKXMIUHGuKFQPg/Wp6Mkg6KJUfpetl4rDQrma9CqLPKegfX
0YDG/T8/z3usUlzGF+F03f7Qhf89ry2DpYK2wmUPQKGjiZhne+6jXoqX5XonyKQDimx3Pp3mmIIb
xW6PeZd7cLfTcvGYuSgvxM2MdCfhlBPPaRpVwyQ6kNcb+EnufAXWTu0vHjjzR9ZjqGGhmoBKfuax
bOkhRl3dQ0KY8QUiirrlM3kmi84rCMjTM0dQfqdGlBxOpgfNQh9sHJ5K/nOlTEqLRZPd96Xsai2d
M6POQYymc17LAGoMR7FI4G+f6sXV2mBuKa3LfGRYlR53ql5OBW0sXQq5BMFGhCeTJFC+B7wfMVFj
fvbQKYY+lWjWgp+yEUjpEA/SV4gQy+KzgTE0m+QagZQakyGya3C3hKPrzBkg7yfFemI3ngxgjwgy
YMkb41zoOe/mpXVXwDHOFv4B+7trHuvFBHso37pmaMBUyKFpdrzcqjaM+lOt+VX3+ZtUQuPM0ofv
ILaUSmduFtMwqY36PoEtyrRVtTehf2e1iRGZpBMxiEfnWrCm4avflD7ir0OAN+y2W5y+Azbte8jo
k/YvPamKwEsKehfAMSGLAKdlpOYQGybyPZeqYMH4bDpLEbcsBdKPGvTTZM7EyEROnIcQi/rI9s/s
l77UakUbo2N6aJBnRqum+LHg4Zj08fCNYeMk+yYwo/WAft4edMxOJPSUxTyfdNIP85rTNZHxiGOe
XduQj1Ewd8dCcqtPP//mqOm2Y54eHND99s73I4tYq7qhMP4nYd+0rHi+HtsTGbYQFtQAZV4eI/Fh
ssfbXU5NqVgeeTkaEptiiV202hVDAMDXYcd3v/MWJS0wrFiPzz788mycCd5YXtx/D5htxvp0+pyq
tBQqSBblfB8hYqncxXkVbXhR1e/uis7ZTAhadSkPb6TXAbZPorqYN3Bkawi8UxOXJ2B3jsRKecTM
QeDT1QphZe1HLYGtQDEYzJPzMqA8utAvMCPJz6TC00BrmhJZUNzf0EPkb4Htf14Bubx18DzhUrA0
mCN9/lBMNQ4JmbZkqbNZ0kGqn6V1hNMj3SvfRME0O/YLZcKiyDrjDgfbT2leaxEEvdWz3mc6gG09
bbf0HUbwy5TGujCO9iNRqI9yuUiBmMOO8VdrcBgzYXcY/8K3bHj2AWw/QCSUcIWkqFAsLR8hi6O0
lqFw/vdDqZ57ICvMubT9nwKXHQtNDPBUtHEr5grslcRq5Aywph8c/lOmR5jo1U6YuKdU2mYZx/Ej
CdJ4E1samQprtXfSaFXbTHWqmMPkPRPNes+q2tYmKG5WEszTckb5RsE91lvmw+11SoxQ+Onmclqb
95u4vId/7MG3ktIZJPc0JXWB1VaBTbxcmy48aWVRuFBzTGpYuT/5NDnMd7RQfJvLpm3u6/w44kXU
FV5WUzxYZckxw8xlW4n+NsIF2Jcd4TEgB7uQw89fBLQiE5VH0Okd6q+S//qE89/Y8x3B5HTltHJ5
zZwbW/Vgk/acm9BODfEZkd0i/B9kfdCmnTxfJTauYmNQ7yAd348hWsBu9pwB44wM8Fp810uadIOl
bFSfx+O/stPBfPKSPr8B6TJ3hDGGakaGXdVRurQHAHgtp3j8Ph0Fat0Lqd9wyaWGcbiu+tI2xBwX
Bpb5BK1AHU9N/202wkWYTCNWSe093r/cDRwyy42y1TINEAFilFIowbNl4+1b+YYYF4U+TdUUkNat
kKqeRj/+AyJCb3cCyHo4VvZ5rT+ZUyvOPkF2gRUOQzmFPwohixYzzZkBEYiboddb59PEbGjv8rM5
RAyD5AxLbxYZEsUpHplODoTaIIkR4OLZ3S1xx3eYfq5MYxIJuz5TALcpGq5b10A5YNOj1UqnADTZ
+4ir0o8xu5MnwozjOwRMe/TPtHUEbbDuVQlZQrImVAVDDVDNaBacCXjUaqOduQrSMbAALdqxDZCv
K2UIS1V32P+newHzmhZuYUtAEZvaFmF25SeK1OZJhsqkOaz/xJMrrmG3m1LIHTssp0iwAlOZkljp
0LI9pw6qeIkklHQGrLJzRUNoCLp4sG6k6M5gJrhTGp5juoQ+IRPCvkkldnCZe18upnVxNR5qM6I3
68OGsWXxYBWvhmfxi0U892WEgYu1M8YCoD4yhBp7OqdCLa3+tVjfYBGuCs8DXWq9k47aCMAh3gqb
na9xthJYuHrMHvMTTcbtihflvE6RkJrJwdpAYwjD6D8fW5O3bgVvoOdPgFeVFW7HJvpct6EQBTEn
rv2HY6O/+xzZvr8oGEHAaj82hHlizIMn252OCcVewGX7bvhIoc81bb7BNuJ5DufnfB0tskfo5xkD
0m3rDiQ7XeW5VVEjB3haFuLrzvBzjfYqRsvQrIxJdbrFssUEicqhjwF+RRlu4OXKy63VgjxxBmDV
wi23nxK6LTXEkYqzJ7f2GgYhB4vpbtdLPFm8hfL09prktSyIRkbCAUQlN+sK/eYa6EejQQgcAekD
KO4fF/8YkSO9XGoTatEN03hxHTsgFUO1xuhDl1Ex85a0rXmBwI2VTNUz7ht/IYa9d3fT4BkqHj/W
zJIMTor2O7iTJQmEfTqRNtRvjApVPrZg+pn1q1ZrQpZtuj6RbTfQbVG/63YEe1yOyH+cJWSO5GDl
JUqfehxiHhuVUSXkOC/VfAlVMaX0HJwNlD61PwASx4YaGNFhkmGSKxB/jPsqXJQtQsgQU/qDrlSr
69H1kCLNyE5XmvOHXE+oPlrTaGZTNYpTT6/LcfyQULeZOp29Tt4UuPC/F6/W6i0pLXIOegV3+Q6q
mdvnSPvboUKgXJjiuUgdYUIioFSPMv0m/w1ZtAXnvE/pqKK7qlKYDx+iG6VHG++p+Ej2E4aAmwVd
VoKeG+5cJIj8VyW9vi4zP+r4naB2eV6tVvJ9SkMAqnWUxoFC/jpF0AgFT9Mos0ZG24EgtM+g9Oib
euqvBsEaFwFbD9lajLMwwzvYe2E0XuYn13guSX7erTg6+HCLG7ZRUc2B6WHTDqCN2rsgEvrjmHBd
ZmvJhsHIkbrg6EZACHeRrsolPu1m4LNeHtu5TnPf7mnToxpqWFVJGAb3OAfaII0L38bnIpadNWjE
lNnSSPF4UXOduS27ozMg0Jx510WWIUURpKNkAnzsG8YhpwFlf0G/0pofOGN4f4XCzvptHVuSbfLa
YkklaOaQ2UFbHLPZWW+GzCQxvseDqUNpk15fkuYVWdBhdTkILo3hTShkk/3gZEv/dPJCsv1peb58
7Y/B3yXzhEwsiReQweumZ/10FHF4gIAwu0cdfJeBYczBmfA9e2ACjebkYWg+SOUsVjB5LPnddhjt
jL/N3G28bLqLBmgiDqfwIP5CeO5c8X/wW6Tye7IsC/pZwGuZ2QWU5OCFsYlI0E5zXZ4kl6V6s8Jt
EMziHRfGTPxb/yMTQSDQl7JWTCKAEfh0b85PypXR4/TCDm9zPNls2NIn7WyWhvSrk0XnX2LA5uVp
62yfTmBFc7B5axuCuoOhjE1Gsk0FQQai63jcS67HBl+XgkhfHY18ikUK24xHy6C6hLUmeD9L9MLx
WpgJUEgcWkmeEjrTokeBdbAjHLxgApurrfHFDQE0IbUW6fx4cdZk8bIhy61NQI88X+LfrKHNa9zG
EFVfzo4cURD/eE11Wp4dHUtxEIxMkCOJQ0VOrao8TSyNnE6nNCz666kHAPs+UXWJmBxWH1cUlgH9
Lt2BhOfV04BCJvTIhdU6BhPRVTRYc3yIGza9DBRAXVVLv67m1Qmo9jbZd4+oa/9lpnx3WsNJ1EiR
8iHy5oWf7PJV/PzE6yDGX0hvgOevvXOGdjv4b0fU3NSYUvOG43jIv+6GL72T7lffuMXgmHdcNdRG
aTqFSIWyHRlBCChJ4uWiBx8I0oYwwHxrScdyRTdWeR/vOwNLMwWA9zGYBWTLdB7lFoomB4ljljoQ
z9vHU0fN16wXejhAdlTQ6PKrC613RUW7NGMzYCbCLHq58lBES/1CTCLg73hc4RbsOyX2yX1NCwBt
Rr3VvZFgXO5ldm/N/llRcXoIKfCM67/rFfN+LL/wWxwMa/l0v7DY6kjPg3n9xlTJtCSdeC3sue22
g4hGKFVI01X2OrbGF43TB7irSQomBxjCNV37X+ycNg9c09qhNkWTjhr1mBsN+3gwCRbVYg99hQrC
cAVE7XUzk475iwUccDxNAL3Ynyo6wFQd1D0VeaVhQTtrPgg80EMPcU97APjbGU9zcH3xe43ixT+m
WvL651ZFcKgjtfpMY2cUhICvBqQAI6TAhuzhdWmb49hxjqDV2XAb7l/YYoABgG2R8FlrsRmZSHcj
0yT2b86Us8REF/DflU5aWchOc4S9CEpVzzOis4PVcENlgmq2wApuXrNXgaMApmcpuccekAIpx9D3
9fwqg2BhI2vL+sjgiYFAzcLg5sA3HwxTBWe04DpLyjUIiTsKFwmmZASOlukiT0ftVkhs0oRT+CbD
oj3J7/QCyTcRTgH1UrWSrhO1S8n3MFxSzsX48UbI7WvpYEUfePYDF8pU/UyALaZntTaHx6F4DvLw
lsqidyTE63MCsxFAcuyImqSbsiYEoE0GjcDGEADmmpJhWnRD0n36DSBSLkTLDN0Ku2Q3y/BuplbH
7l+iEXaw3wfmbVOXaxhtOjwlpPNruv85MRg29ShnXYzhJajueIsU0GsA9Asg8TUM5V8W0dto685Q
kqLMtLM32Z6j4fyQkmqkWdic59nsZyEmhzguGTAHjZcVJvljxnraMCNIfPypWKIIg2ACx+uIQ66N
f97FHiiqLcnZqtEW2y+9JS7b9jtIXQAph9Wy/FxEqWWgsEgnOE2Ofvb0WJc0hv/BjcaaBCgplO0M
oRTBMXrWaQ6X1uZ+zu5mDf+FCZSkBQ9PKLeD32W1xvvJNbZ5l1C3Fb69/sPUVdqXzIt98X9/05I/
jdz5MbLRbc3M0UhKpTIIrB5+G1YQuklaB6lWphcV1Mvnsdare1V3SGHmgwlOs4xC8GrzzH7wpsNV
cNi3Elo1GgApeZCFevgboPfWwEAY7oMeXMuepaM4J8tBTWAZEf8b70gW67vu7RKD9i+BgA2bCCQl
lVkDRSvTzT3q2wDNNDOKa9FkHv6wu6yCEG/krT8Xlk92WsWN0z88Stnb7/0C/uf8Jq7I7rJZQlbi
AbzSOJyxljl2tpfbL7d2t2JBZcKfFcjfenh7+K3MAGzxDwEbdfnwBquJifGCptO6QEy+K7ykyIWA
9oR4LDROo37h7WQwiAQj0KhGabFn1jTxs6yO/tgdldtVArE3wPqrfpbgr7z4c8b02eYmVjl/qIZF
4E8UIVzzecHv18jGIoCFYaBpmh/EeUnmZM8FPeKy0tm7QDehpC4uycR5HEzjyo6z0u6sGo6C3ZHV
DzJs+IPUuBSbPzVoWrjbs0mRJH8CMXtzObUw3jqyJZwdSKdI1kLB3xAj6iQx5mgv+7Pr6JbUHFU2
8mIQuJ2caZvRWbRQrutxUr7WqqyPB4KFXPrVXoxR4sdF+4PobHJIbk64cAxdBEiMSn2asF/71MY/
riIhUiVSNpeLNxKA9mvhvI/uMFrag7jYqWfBtEGglvgkiqGCwdAizzR5w0gmJKVZqSfgEcSV+eXU
j5W5ZI1CABokQtozMBE2UiJncdfinsxy4tZ3Ez2mmtSW8IpMFGjWPYRvHn1m0e+gEbAh88Mc8KSH
pGQvNMtwCydJUCrlFU7RRfo7Usvf13IEzljYe+qT+ADXO4QyXjdl7Narn6bQ+VWXQMdlJtakyc0/
0/RMcBZqcgwbD/uAa+W5cLVSaqf8M1If0xysLdwAzlURcOmilQ9NmlyReMWiBRYsCJ7359F7qbTo
lrFpVsaCG5js9iVRIbpYlkV7K/Ok4hKXVDErPKDjWWKlFzvCG3bqgnTIPfuoBxgKlSbna4+Voz6t
u2M1CvfBYGacMGqXcnKKo9tmv3a+yyifHiUge00K0fJQxU34V8Sb6N0we/e6nrBlmj/AWbZ8FPg/
ww6C7RjD5Gd8Zvl1Bz2ykscxozdhZpM6jp7t9ZmGaaXWdK1yrRD8OnEhPwGS4AHKZYf0pI2WgcSF
p/8CwCfQhRLC3QavH1QkKiZv1nCeMzmBafqXZxupDGlE8vBB6g9F3JxTwPtaT2G9dY5tMt4JB6nm
mYLaMcGfVwj8RCNFEx9rCrZlFVhF5onSnqID5NNuSbRPQEhH6dOVd1DYZKlS/RiaGbsw0ip0T6Rd
8ar+tzmhCgE5Asap0Mi7kA1Lt9UYEVQFrXJz6CWGAx8CHP4k+Dw9xnCLoibrzdxj5VFhAHT7IAmf
NcNB2jM9ylY5IeeqOHqDA71EQFAPhm9u8mM+OPmcNJCUJfCTNZZ1hJ43FiI4b5+71cLqCVcW44Vg
7le/BEiHQt3avSG/MoKbqJirG11rrE29cMWcckhNH7HCTjHkUKiPNMbe5Xf26QKGzyDQqxKMm25B
rhzTlyVoOXYtmmcTdL58N85H9CRC5YfbGDYg8c9DmnHchhYFdzVWmFcDKiT4TkaBAe1aCinj8oHl
2bnMbBY+S8wD27iOmv6RUOgOquRidaEpHElH5JF3l9oUm8dXmPiM5Fv/zN43JkJZkZ45JdhOE26K
n8APQPvA7g+qAEkrM3KuSmgT6W78O8/hFXplcFu+T0wk80w+stGSE88zVGx6uUP44tGYmZAh32ZK
w/hTJD8ZKZsAogqJpsoefT6/wsd8MD8b8lljVdKlryVHn1kK/Av5xMHgIO4yF2AmoyucJLE3RCjb
8/0pt3/3QZGFxQ4nyPhWBfd+SJQJd3NQWhKGOrStuOnoaaYlWKdJVYqES6RRAo5HgBWtlaQ6sC7f
00lMnqW25igs46blnbXhazboq6P47naQ1/wmrqwSweoyBN/A9ysaEuNHdwfl8j7Rea4a6HKPOn70
Yn+FHbRLQ33Eyqrt4hgTXGmg7XHTm3dQQc8Eujg4yg83HmANATGI5sDAQ639R0CrkUnuK+isZCnZ
/gnnvcOT28KUrybGLI220dqbtRdMGK4g+4q9K2KS337iXPY8bqsPUtuJ3W5rdOCXEkLfHBCWlaYC
LvFjNB9t1hxJOD9qcfWi7Oqwi43wV+Fk2S3DHXxfntNx8N82GhxSnxn/aROMQsODgO1uhXe3b3q1
PAel7CebevT3ZhknYCvGmjFM5D1AkgQisvPd2NSVO4RnphsmcRL2m+sV64GNjwUme7tKN665bcOe
+sXqNNZIrfOMm/xN9rsXiLDe/2zA5vGe85O/d+le1lMc2bq9y7yvt2jNmid6IX1xqCWOmVDrWTO+
s/WbWozSjqsBhuJ81lWti3YSdsiu5SJn3gCGP6+Fml44xEx4MHsd6ZYPL+YCPlDFMlBeNGV9yYt8
/tdozFrTGy3fyajBnQnUo17wDlIEgIkMeFpKLAZgvRbWgq0FmhgxoGLhPHJTNyEiRXhZHuZ5Pt6r
SCCmGuyXWAx0jjonx5rQvS5AUufWDskQm/cf69B0uBvSxMpxHT/4yZ4iQUM9yFbRA7mYdUP/tTRt
frEUHi9h036nUHWhHahthc+sZ2vZ5pqakR39xv7sk9/6K5Ewvk1Bq/qLJbY4EF7ZW7/p2n/qJOn+
coFAR2UKbBEb4tbJdkzUZiH0+3IkAuAwpTUP8OqI53YM31Zdd7MZ6OKfT2kiMJe2xHFGALbqrWiR
K2x+77jV1kO8WTKwJfKy3dPUMa2QUzJT4zM6y3wNR4sJ1S9qYCahRGZSHp8vNLd/JrSkpJTobqx2
u+lLwMPnAq/8+zJjWPVJx/MKAp3O/RPrK9nAnM1OvOM4lpKSEt59lyZ9m6IhRg8NZvtCRJZqheeM
MmygQNbohRBK/wyq8ikrSI1mQjVv+sfBi9uRl6V4J1ejh7HkKghszLw0+4DJ/PVyTJXEfhnsPwHm
/3Z/4CwWZ53CMPe+XvdENKUoyMdyvL2BiIdH1JxYO4sCOI7qJCu1Ux3UYFig9MZVliVOPI8yJ0FU
XgEuMuS4n/X38T+0CAVWFvQzCl6HM2h0Frot0xl3vK7zTtON3X/Vjxsg2a32TaQ4IbARYXH9mPW5
dxbnwbjn/io+r9WFaZsrigd07BZznvhT2D0w38UWwctykhZ0voMCR0+u0e8rEZXmH+XVC61wFZat
m+lFjAyIHSGDF8ykd2pWw0JHwlNLk+Ry/gAmjNCb3Gos5x2aLWpUeotALnchjGHKWcRs6auC0D1L
izbRanMFFu2a51e1KWXFWMZ8GXRs9/UW+tT66xbBaLLKb1YTOIu9c+W+E5RiAlzv63Fko+rGgpPA
CVj/N9/jsWVp1QjEuh2QcG47TYO0l3vADtuIwAlOf/zuY2tMvJzABsWSFr9+sj5uPnMu0Uu+0a6b
lnX3Kaoj0ZziB3Mwk3z9/EOPS4BnEHC3iW1IKTlxGoqzI+IGL5aqwiW94MZVOWM8H7CbCzGA0DME
wMFjTeCxGrtGXkMOJolSdaXX/OiIUNfzNJJn6egJyyKKn96KUMrTBW4+z/UWvFX6GyQYcrXjriog
WBe3NYSVbhZFqk7XVPYmW9YbUi2fbpnJ1vjEtoEFL7Zbxo64kL7W21Pi3MqvuproMPzPP6JKLjSt
8aBDjFJcjuZ2EfxgqgoeBRXgYXRLZLPbmrxGhWOnVBGtjk8i0S1jvWg51vJYE6YGleRBIX1VXdES
VwBS5Y5nWOLCTB4B0CKTE3Ach4teqoXiu32TnVG/Y5k9+EADNcSTIYSWfDr5cOJlXEcX5hKc+KS9
UEAVfYwrgGCWzGzFTcQzwwYsoMjd0HwP2h2HxYw1g4cd33dQWCa4ecDqDeN/rwUyjqAxcHiw4q6i
IX0r2+H7Xy8Qw7THeLIj2yqdu4Ial13jl5K6S7YZSqd3jb2p3Ez79syvKHtZiWvLC5u2FpKhD1Ig
78ehux50nYb7GZQP3frxM3E2kxptsBhFMwCx8+YoPHzHqxuhRN7JvOghPoOFxApDrUyVgj7BqugW
mK3Cx/al/FdJuxT09qGT+QNWX+VZ3iaJyLkrPUP2lGRRikzXkJ5MoTGRAOWyBCqlQG3gDd4=

`pragma protect end_protected

 endmodule